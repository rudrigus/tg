 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 03 03 03 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 04 04 04 08 08 08 08 08 08 06 06 06 07 07 07 05 05 05 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 08 08 08 0d 0d 0d 16 16 16 23 23 23 2d 2d 2d 4c 4c 4c 31 31 31 28 28 28 13 13 13 1e 1e 1e 3a 3a 3a 4d 4d 4d 45 45 45 34 34 34 34 34 34 35 35 35 2d 2d 2d 2a 2a 2a 2b 2b 2b 1e 1e 1e 19 19 19 13 13 13 0c 0c 0c 07 07 07 05 05 05 04 04 04 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 08 08 08 18 18 18 32 32 32 57 57 57 6d 6d 6d 7e 7e 7e 95 95 95 98 98 98 99 99 99 84 84 84 5a 5a 5a 52 52 52 50 50 50 56 56 56 5b 5b 5b 54 54 54 4d 4d 4d 45 45 45 42 42 42 44 44 44 46 46 46 48 48 48 66 66 66 93 93 93 92 92 92 7f 7f 7f 55 55 55 44 44 44 3a 3a 3a 1b 1b 1b 0c 0c 0c 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 12 12 12 2c 2c 2c 4e 4e 4e 67 67 67 81 81 81 9a 9a 9a ad ad ad a0 a0 a0 8d 8d 8d 78 78 78 6d 6d 6d 68 68 68 6c 6c 6c 6d 6d 6d 6e 6e 6e 6e 6e 6e 66 66 66 63 63 63 5d 5d 5d 59 59 59 51 51 51 52 52 52 4e 4e 4e 4f 4f 4f 5d 5d 5d 6c 6c 6c 71 71 71 69 69 69 64 64 64 66 66 66 78 78 78 64 64 64 55 55 55 2c 2c 2c 0e 0e 0e 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 0c 0c 0c 1c 1c 1c 42 42 42 5e 5e 5e 63 63 63 6c 6c 6c 72 72 72 7e 7e 7e 90 90 90 99 99 99 97 97 97 8e 8e 8e 78 78 78 70 70 70 6f 6f 6f 80 80 80 85 85 85 87 87 87 82 82 82 7a 7a 7a 72 72 72 6c 6c 6c 6b 6b 6b 65 65 65 5f 5f 5f 5a 5a 5a 54 54 54 5f 5f 5f 6a 6a 6a 6a 6a 6a 6f 6f 6f 71 71 71 69 69 69 67 67 67 67 67 67 8b 8b 8b 94 94 94 54 54 54 1f 1f 1f 0a 0a 0a 04 04 04 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 1b 1b 1b 4a 4a 4a 91 91 91 90 90 90 6a 6a 6a 6e 6e 6e 74 74 74 76 76 76 80 80 80 8f 8f 8f a9 a9 a9 ac ac ac 99 99 99 80 80 80 76 76 76 77 77 77 88 88 88 92 92 92 95 95 95 90 90 90 88 88 88 7d 7d 7d 79 79 79 77 77 77 73 73 73 6d 6d 6d 64 64 64 5b 5b 5b 61 61 61 6f 6f 6f 7a 7a 7a 85 85 85 80 80 80 72 72 72 78 78 78 73 73 73 73 73 73 7b 7b 7b 75 75 75 50 50 50 28 28 28 06 06 06 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0d 0d 0d 2d 2d 2d 6d 6d 6d 97 97 97 97 97 97 75 75 75 75 75 75 7d 7d 7d 87 87 87 82 82 82 92 92 92 98 98 98 b4 b4 b4 b9 b9 b9 a5 a5 a5 8f 8f 8f 7e 7e 7e 78 78 78 85 85 85 8d 8d 8d 8f 8f 8f 90 90 90 8b 8b 8b 88 88 88 82 82 82 80 80 80 7c 7c 7c 79 79 79 73 73 73 68 68 68 6c 6c 6c 80 80 80 94 94 94 99 99 99 8e 8e 8e 88 88 88 8b 8b 8b 87 87 87 7c 7c 7c 7c 7c 7c 7b 7b 7b 62 62 62 6a 6a 6a 27 27 27 05 05 05 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 15 15 15 3f 3f 3f 7a 7a 7a 70 70 70 6d 6d 6d 75 75 75 76 76 76 7e 7e 7e 8c 8c 8c 98 98 98 95 95 95 a1 a1 a1 ab ab ab b8 b8 b8 b7 b7 b7 a6 a6 a6 9c 9c 9c 8d 8d 8d 7f 7f 7f 84 84 84 88 88 88 8c 8c 8c 91 91 91 96 96 96 90 90 90 87 87 87 85 85 85 87 87 87 89 89 89 83 83 83 78 78 78 81 81 81 97 97 97 a8 a8 a8 a6 a6 a6 a0 a0 a0 9d 9d 9d 9f 9f 9f 90 90 90 84 84 84 7d 7d 7d 7a 7a 7a 6c 6c 6c 84 84 84 5c 5c 5c 18 18 18 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 25 25 25 51 51 51 59 59 59 5e 5e 5e 65 65 65 6d 6d 6d 77 77 77 79 79 79 7f 7f 7f 8b 8b 8b 9a 9a 9a a1 a1 a1 a5 a5 a5 ae ae ae b4 b4 b4 b0 b0 b0 a3 a3 a3 a4 a4 a4 9d 9d 9d 8f 8f 8f 8c 8c 8c 93 93 93 96 96 96 99 99 99 9f 9f 9f 98 98 98 8b 8b 8b 92 92 92 96 96 96 9b 9b 9b 9c 9c 9c 97 97 97 9b 9b 9b ac ac ac b2 b2 b2 ac ac ac b1 b1 b1 b1 b1 b1 aa aa aa 98 98 98 87 87 87 7c 7c 7c 76 76 76 77 77 77 80 80 80 9d 9d 9d 46 46 46 10 10 10 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1c 1c 1c 6a 6a 6a 67 67 67 5f 5f 5f 66 66 66 75 75 75 78 78 78 7f 7f 7f 84 84 84 86 86 86 8e 8e 8e 97 97 97 9d 9d 9d a1 a1 a1 a7 a7 a7 a7 a7 a7 a2 a2 a2 98 98 98 9d 9d 9d a3 a3 a3 9d 9d 9d 97 97 97 92 92 92 8d 8d 8d 90 90 90 90 90 90 94 94 94 97 97 97 9e 9e 9e a8 a8 a8 b0 b0 b0 b7 b7 b7 b4 b4 b4 b0 b0 b0 b3 b3 b3 b5 b5 b5 b5 b5 b5 bf bf bf bc bc bc af af af 97 97 97 87 87 87 7a 7a 7a 76 76 76 76 76 76 72 72 72 ad ad ad 83 83 83 31 31 31 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 3b 3b 3b 81 81 81 68 68 68 66 66 66 6e 6e 6e 77 77 77 7f 7f 7f 84 84 84 8b 8b 8b 8f 8f 8f 92 92 92 9c 9c 9c 9c 9c 9c 9c 9c 9c 9c 9c 9c 9d 9d 9d 91 91 91 8b 8b 8b 90 90 90 9b 9b 9b a2 a2 a2 a6 a6 a6 a1 a1 a1 9d 9d 9d 9b 9b 9b 9a 9a 9a 9f 9f 9f a7 a7 a7 ad ad ad bb bb bb c5 c5 c5 c1 c1 c1 b5 b5 b5 b0 b0 b0 b1 b1 b1 b8 b8 b8 bc bc bc c0 c0 c0 b7 b7 b7 a6 a6 a6 8f 8f 8f 82 82 82 7f 7f 7f 79 79 79 71 71 71 70 70 70 83 83 83 97 97 97 49 49 49 0b 0b 0b 03 03 03 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0b 0b 0b 2c 2c 2c 4e 4e 4e 70 70 70 73 73 73 69 69 69 6e 6e 6e 79 79 79 7d 7d 7d 84 84 84 8c 8c 8c 94 94 94 97 97 97 9b 9b 9b 9d 9d 9d a2 a2 a2 a3 a3 a3 9a 9a 9a 8b 8b 8b 7f 7f 7f 85 85 85 91 91 91 9f 9f 9f ab ab ab ae ae ae af af af ab ab ab aa aa aa ad ad ad b3 b3 b3 c0 c0 c0 d1 d1 d1 cb cb cb bc bc bc b3 b3 b3 b4 b4 b4 b8 b8 b8 c0 c0 c0 c1 c1 c1 b9 b9 b9 a7 a7 a7 97 97 97 8c 8c 8c 83 83 83 7f 7f 7f 77 77 77 74 74 74 6e 6e 6e 68 68 68 65 65 65 66 66 66 28 28 28 06 06 06 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 06 06 06 27 27 27 49 49 49 5b 5b 5b 68 68 68 75 75 75 6e 6e 6e 6f 6f 6f 75 75 75 7a 7a 7a 81 81 81 89 89 89 94 94 94 9d 9d 9d a1 a1 a1 a1 a1 a1 a4 a4 a4 a7 a7 a7 a2 a2 a2 8e 8e 8e 82 82 82 82 82 82 8d 8d 8d 9a 9a 9a ab ab ab b8 b8 b8 bb bb bb b8 b8 b8 b9 b9 b9 bc bc bc c5 c5 c5 de de de e7 e7 e7 cf cf cf be be be ba ba ba b9 b9 b9 ba ba ba ba ba ba b8 b8 b8 ab ab ab 9a 9a 9a 91 91 91 87 87 87 82 82 82 7d 7d 7d 79 79 79 73 73 73 6b 6b 6b 68 68 68 5d 5d 5d 67 67 67 43 43 43 06 06 06 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0b 0b 0b 3f 3f 3f 62 62 62 59 59 59 61 61 61 67 67 67 6c 6c 6c 6e 6e 6e 73 73 73 7c 7c 7c 7f 7f 7f 88 88 88 94 94 94 9e 9e 9e a4 a4 a4 a9 a9 a9 ad ad ad af af af a9 a9 a9 9b 9b 9b 8e 8e 8e 8b 8b 8b 93 93 93 9e 9e 9e b9 b9 b9 d8 d8 d8 df df df de de de cb cb cb cf cf cf e2 e2 e2 f7 f7 f7 e9 e9 e9 c8 c8 c8 bc bc bc b8 b8 b8 b6 b6 b6 b6 b6 b6 b6 b6 b6 b0 b0 b0 a5 a5 a5 96 96 96 8d 8d 8d 84 84 84 80 80 80 7b 7b 7b 76 76 76 6f 6f 6f 66 66 66 69 69 69 69 69 69 67 67 67 50 50 50 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 09 09 09 46 46 46 5f 5f 5f 57 57 57 5b 5b 5b 60 60 60 6a 6a 6a 6e 6e 6e 73 73 73 7b 7b 7b 80 80 80 89 89 89 90 90 90 9b 9b 9b a1 a1 a1 a7 a7 a7 af af af b1 b1 b1 ac ac ac a0 a0 a0 9d 9d 9d aa aa aa a4 a4 a4 a9 a9 a9 d9 d9 d9 fe fe fe fe fe fe f6 f6 f6 f6 f6 f6 fb fb fb fe fe fe fe fe fe de de de c5 c5 c5 c0 c0 c0 ba ba ba ba ba ba b8 b8 b8 b5 b5 b5 ad ad ad a0 a0 a0 9a 9a 9a 8c 8c 8c 84 84 84 7f 7f 7f 7a 7a 7a 73 73 73 6a 6a 6a 60 60 60 5f 5f 5f 64 64 64 68 68 68 5a 5a 5a 0a 0a 0a 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0b 0b 0b 43 43 43 6f 6f 6f 57 57 57 5d 5d 5d 61 61 61 68 68 68 70 70 70 75 75 75 7b 7b 7b 84 84 84 8a 8a 8a 8f 8f 8f 94 94 94 9a 9a 9a 9f 9f 9f a7 a7 a7 aa aa aa a6 a6 a6 a3 a3 a3 a2 a2 a2 be be be d9 d9 d9 e4 e4 e4 fd fd fd fe fe fe f3 f3 f3 e9 e9 e9 fd fd fd ff ff ff fe fe fe f1 f1 f1 cd cd cd bc bc bc b5 b5 b5 b1 b1 b1 b0 b0 b0 af af af a9 a9 a9 a3 a3 a3 99 99 99 93 93 93 8b 8b 8b 80 80 80 7d 7d 7d 78 78 78 6c 6c 6c 64 64 64 5a 5a 5a 55 55 55 4f 4f 4f 5b 5b 5b 5b 5b 5b 0a 0a 0a 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 12 12 12 4d 4d 4d 80 80 80 5a 5a 5a 56 56 56 63 63 63 6f 6f 6f 71 71 71 73 73 73 79 79 79 7d 7d 7d 81 81 81 87 87 87 89 89 89 91 91 91 96 96 96 9e 9e 9e a3 a3 a3 a5 a5 a5 a5 a5 a5 9d 9d 9d a7 a7 a7 ca ca ca fd fd fd fb fb fb ef ef ef b2 b2 b2 c9 c9 c9 f4 f4 f4 ff ff ff ed ed ed c4 c4 c4 b3 b3 b3 a8 a8 a8 a3 a3 a3 9d 9d 9d 99 99 99 98 98 98 95 95 95 92 92 92 8d 8d 8d 86 86 86 80 80 80 77 77 77 76 76 76 70 70 70 68 68 68 60 60 60 5d 5d 5d 53 53 53 4b 4b 4b 52 52 52 59 59 59 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 11 11 11 57 57 57 88 88 88 5b 5b 5b 56 56 56 5a 5a 5a 6d 6d 6d 76 76 76 77 77 77 74 74 74 77 77 77 79 79 79 7a 7a 7a 81 81 81 89 89 89 8e 8e 8e 97 97 97 99 99 99 9c 9c 9c 93 93 93 83 83 83 83 83 83 91 91 91 ef ef ef e3 e3 e3 b0 b0 b0 9f 9f 9f a3 a3 a3 cc cc cc ec ec ec ce ce ce b3 b3 b3 a8 a8 a8 9f 9f 9f 9a 9a 9a 93 93 93 8b 8b 8b 86 86 86 82 82 82 7f 7f 7f 7b 7b 7b 77 77 77 72 72 72 6d 6d 6d 6f 6f 6f 6e 6e 6e 64 64 64 62 62 62 5c 5c 5c 52 52 52 4d 4d 4d 51 51 51 56 56 56 12 12 12 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0a 0a 0a 51 51 51 8a 8a 8a 5d 5d 5d 57 57 57 58 58 58 5f 5f 5f 6b 6b 6b 75 75 75 72 72 72 72 72 72 75 75 75 78 78 78 7d 7d 7d 84 84 84 85 85 85 8a 8a 8a 88 88 88 88 88 88 82 82 82 76 76 76 75 75 75 7d 7d 7d cc cc cc bd bd bd 6a 6a 6a 5f 5f 5f 6f 6f 6f 8c 8c 8c b7 b7 b7 d8 d8 d8 d6 d6 d6 c6 c6 c6 a9 a9 a9 90 90 90 83 83 83 7c 7c 7c 74 74 74 71 71 71 6e 6e 6e 68 68 68 67 67 67 67 67 67 65 65 65 69 69 69 6a 6a 6a 64 64 64 62 62 62 5a 5a 5a 52 52 52 4f 4f 4f 52 52 52 59 59 59 23 23 23 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0e 0e 0e 3c 3c 3c 7d 7d 7d 5d 5d 5d 5a 5a 5a 5b 5b 5b 5a 5a 5a 67 67 67 73 73 73 6d 6d 6d 6e 6e 6e 6f 6f 6f 70 70 70 72 72 72 7d 7d 7d 7f 7f 7f 82 82 82 81 81 81 86 86 86 83 83 83 72 72 72 75 75 75 7c 7c 7c a4 a4 a4 79 79 79 48 48 48 63 63 63 86 86 86 b9 b9 b9 da da da fb fb fb fe fe fe f5 f5 f5 c5 c5 c5 91 91 91 7d 7d 7d 72 72 72 66 66 66 66 66 66 66 66 66 62 62 62 61 61 61 65 65 65 64 64 64 67 67 67 6b 6b 6b 67 67 67 60 60 60 56 56 56 52 52 52 53 53 53 54 54 54 65 65 65 28 28 28 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 19 19 19 2e 2e 2e 4f 4f 4f 56 56 56 56 56 56 59 59 59 5a 5a 5a 64 64 64 63 63 63 61 61 61 67 67 67 6a 6a 6a 64 64 64 64 64 64 6e 6e 6e 80 80 80 7a 7a 7a 75 75 75 79 79 79 7a 7a 7a 76 76 76 72 72 72 70 70 70 7d 7d 7d 4a 4a 4a 4b 4b 4b 83 83 83 d4 d4 d4 fa fa fa fe fe fe ff ff ff ff ff ff fe fe fe de de de 94 94 94 7b 7b 7b 6e 6e 6e 63 63 63 61 61 61 62 62 62 5e 5e 5e 5f 5f 5f 5f 5f 5f 60 60 60 69 69 69 6d 6d 6d 6a 6a 6a 62 62 62 58 58 58 55 55 55 54 54 54 5a 5a 5a 6d 6d 6d 28 28 28 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 1f 1f 1f 36 36 36 45 45 45 4d 4d 4d 51 51 51 54 54 54 54 54 54 58 58 58 5e 5e 5e 5d 5d 5d 5e 5e 5e 61 61 61 66 66 66 5d 5d 5d 61 61 61 67 67 67 6a 6a 6a 6d 6d 6d 6f 6f 6f 72 72 72 6e 6e 6e 6a 6a 6a 66 66 66 6e 6e 6e 3c 3c 3c 59 59 59 af af af fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e5 e5 e5 95 95 95 78 78 78 68 68 68 5d 5d 5d 5a 5a 5a 5d 5d 5d 5c 5c 5c 5c 5c 5c 5b 5b 5b 59 59 59 60 60 60 6e 6e 6e 6f 6f 6f 64 64 64 5a 5a 5a 53 53 53 51 51 51 60 60 60 6b 6b 6b 1a 1a 1a 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 1c 1c 1c 5e 5e 5e 5f 5f 5f 52 52 52 52 52 52 57 57 57 55 55 55 57 57 57 5c 5c 5c 5a 5a 5a 59 59 59 5e 5e 5e 5e 5e 5e 54 54 54 54 54 54 58 58 58 64 64 64 6b 6b 6b 6c 6c 6c 68 68 68 65 65 65 63 63 63 62 62 62 65 65 65 3d 3d 3d 5e 5e 5e c3 c3 c3 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d9 d9 d9 96 96 96 7b 7b 7b 66 66 66 56 56 56 55 55 55 5b 5b 5b 5a 5a 5a 58 58 58 58 58 58 58 58 58 5d 5d 5d 6f 6f 6f 68 68 68 5f 5f 5f 58 58 58 4f 4f 4f 50 50 50 68 68 68 59 59 59 0a 0a 0a 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0f 0f 0f 59 59 59 79 79 79 5e 5e 5e 53 53 53 5b 5b 5b 58 58 58 60 60 60 55 55 55 59 59 59 55 55 55 59 59 59 58 58 58 50 50 50 51 51 51 55 55 55 62 62 62 6a 6a 6a 6c 6c 6c 65 65 65 62 62 62 5a 5a 5a 56 56 56 57 57 57 3c 3c 3c 56 56 56 ac ac ac fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe c2 c2 c2 8c 8c 8c 79 79 79 64 64 64 55 55 55 4f 4f 4f 54 54 54 55 55 55 54 54 54 55 55 55 57 57 57 5f 5f 5f 63 63 63 5a 5a 5a 58 58 58 53 53 53 50 50 50 50 50 50 69 69 69 2d 2d 2d 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 08 08 08 36 36 36 70 70 70 5c 5c 5c 4d 4d 4d 4c 4c 4c 4e 4e 4e 54 54 54 5c 5c 5c 54 54 54 54 54 54 59 59 59 5c 5c 5c 58 58 58 52 52 52 54 54 54 5d 5d 5d 62 62 62 66 66 66 66 66 66 5f 5f 5f 53 53 53 46 46 46 41 41 41 34 34 34 46 46 46 7b 7b 7b d6 d6 d6 fe fe fe ff ff ff ff ff ff ff ff ff f9 f9 f9 a5 a5 a5 82 82 82 71 71 71 5c 5c 5c 4c 4c 4c 4f 4f 4f 53 53 53 53 53 53 54 54 54 55 55 55 57 57 57 5c 5c 5c 57 57 57 53 53 53 53 53 53 54 54 54 53 53 53 4b 4b 4b 50 50 50 13 13 13 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 08 08 08 1b 1b 1b 4f 4f 4f 61 61 61 4a 4a 4a 4a 4a 4a 4c 4c 4c 4f 4f 4f 5c 5c 5c 59 59 59 5c 5c 5c 5a 5a 5a 59 59 59 5c 5c 5c 5a 5a 5a 5a 5a 5a 5a 5a 5a 5f 5f 5f 63 63 63 63 63 63 5f 5f 5f 50 50 50 41 41 41 36 36 36 27 27 27 38 38 38 5f 5f 5f 93 93 93 df df df fe fe fe ff ff ff fe fe fe df df df 89 89 89 76 76 76 65 65 65 55 55 55 49 49 49 4c 4c 4c 51 51 51 54 54 54 52 52 52 53 53 53 58 58 58 5a 5a 5a 54 54 54 52 52 52 51 51 51 52 52 52 4c 4c 4c 4c 4c 4c 39 39 39 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 06 06 06 15 15 15 38 38 38 69 69 69 45 45 45 47 47 47 4c 4c 4c 4e 4e 4e 55 55 55 4f 4f 4f 50 50 50 50 50 50 52 52 52 56 56 56 58 58 58 5e 5e 5e 5d 5d 5d 5d 5d 5d 60 60 60 5f 5f 5f 5d 5d 5d 4c 4c 4c 3d 3d 3d 30 30 30 1c 1c 1c 22 22 22 48 48 48 68 68 68 8e 8e 8e d1 d1 d1 ea ea ea e1 e1 e1 a4 a4 a4 73 73 73 67 67 67 5a 5a 5a 4d 4d 4d 49 49 49 4d 4d 4d 53 53 53 54 54 54 55 55 55 58 58 58 5a 5a 5a 57 57 57 5c 5c 5c 54 54 54 4f 4f 4f 4c 4c 4c 47 47 47 4a 4a 4a 17 17 17 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 18 18 18 31 31 31 6b 6b 6b 49 49 49 43 43 43 48 48 48 48 48 48 4c 4c 4c 4a 4a 4a 4a 4a 4a 4c 4c 4c 51 51 51 51 51 51 52 52 52 51 51 51 56 56 56 57 57 57 59 59 59 5c 5c 5c 5a 5a 5a 4f 4f 4f 41 41 41 2e 2e 2e 18 18 18 0d 0d 0d 2a 2a 2a 4b 4b 4b 5f 5f 5f 79 79 79 97 97 97 9a 9a 9a 78 78 78 67 67 67 61 61 61 5b 5b 5b 51 51 51 4d 4d 4d 55 55 55 5e 5e 5e 5d 5d 5d 5c 5c 5c 59 59 59 56 56 56 53 53 53 53 53 53 55 55 55 4c 4c 4c 46 46 46 45 45 45 39 39 39 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 14 14 14 2b 2b 2b 4e 4e 4e 45 45 45 3f 3f 3f 40 40 40 46 46 46 46 46 46 46 46 46 45 45 45 48 48 48 4e 4e 4e 4f 4f 4f 4c 4c 4c 49 49 49 4e 4e 4e 50 50 50 56 56 56 5a 5a 5a 5a 5a 5a 54 54 54 49 49 49 31 31 31 19 19 19 04 04 04 0c 0c 0c 28 28 28 3a 3a 3a 46 46 46 55 55 55 6a 6a 6a 60 60 60 5c 5c 5c 5a 5a 5a 55 55 55 4e 4e 4e 4b 4b 4b 51 51 51 58 58 58 4e 4e 4e 50 50 50 54 54 54 4b 4b 4b 49 49 49 4e 4e 4e 52 52 52 4a 4a 4a 45 45 45 46 46 46 21 21 21 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0a 0a 0a 24 24 24 3a 3a 3a 3f 3f 3f 3b 3b 3b 3d 3d 3d 42 42 42 41 41 41 40 40 40 3f 3f 3f 42 42 42 47 47 47 4b 4b 4b 49 49 49 46 46 46 49 49 49 4d 4d 4d 53 53 53 57 57 57 58 58 58 55 55 55 4d 4d 4d 33 33 33 1a 1a 1a 03 03 03 03 03 03 0b 0b 0b 1c 1c 1c 2b 2b 2b 33 33 33 53 53 53 54 54 54 56 56 56 56 56 56 4c 4c 4c 45 45 45 46 46 46 4b 4b 4b 48 48 48 49 49 49 48 48 48 4b 4b 4b 49 49 49 48 48 48 49 49 49 4b 4b 4b 45 45 45 44 44 44 3e 3e 3e 0b 0b 0b 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 19 19 19 35 35 35 3b 3b 3b 3c 3c 3c 3d 3d 3d 3c 3c 3c 3b 3b 3b 3b 3b 3b 3c 3c 3c 3e 3e 3e 44 44 44 47 47 47 48 48 48 47 47 47 48 48 48 4a 4a 4a 4d 4d 4d 52 52 52 54 54 54 54 54 54 55 55 55 3c 3c 3c 20 20 20 03 03 03 03 03 03 03 03 03 05 05 05 0e 0e 0e 1a 1a 1a 43 43 43 4a 4a 4a 4f 4f 4f 4c 4c 4c 47 47 47 46 46 46 46 46 46 48 48 48 47 47 47 45 45 45 42 42 42 48 48 48 47 47 47 44 44 44 44 44 44 44 44 44 43 43 43 45 45 45 28 28 28 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 2a 2a 2a 39 39 39 39 39 39 37 37 37 36 36 36 3b 3b 3b 39 39 39 38 38 38 3a 3a 3a 3d 3d 3d 42 42 42 4e 4e 4e 48 48 48 46 46 46 47 47 47 49 49 49 4c 4c 4c 52 52 52 55 55 55 5a 5a 5a 47 47 47 24 24 24 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 08 08 08 38 38 38 42 42 42 48 48 48 45 45 45 47 47 47 49 49 49 46 46 46 46 46 46 44 44 44 43 43 43 42 42 42 45 45 45 43 43 43 42 42 42 43 43 43 44 44 44 41 41 41 40 40 40 0f 0f 0f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 37 37 37 37 37 37 34 34 34 34 34 34 37 37 37 38 38 38 37 37 37 38 38 38 3a 3a 3a 3e 3e 3e 42 42 42 47 47 47 4c 4c 4c 48 48 48 47 47 47 48 48 48 4e 4e 4e 55 55 55 58 58 58 4e 4e 4e 2f 2f 2f 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 34 34 34 3f 3f 3f 45 45 45 47 47 47 48 48 48 48 48 48 47 47 47 43 43 43 43 43 43 43 43 43 44 44 44 43 43 43 41 41 41 45 45 45 46 46 46 45 45 45 46 46 46 2b 2b 2b 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 22 22 22 37 37 37 36 36 36 35 35 35 3a 3a 3a 39 39 39 39 39 39 39 39 39 3c 3c 3c 3d 3d 3d 42 42 42 44 44 44 4b 4b 4b 51 51 51 4c 4c 4c 48 48 48 4f 4f 4f 54 54 54 56 56 56 51 51 51 33 33 33 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 37 37 37 44 44 44 4a 4a 4a 46 46 46 46 46 46 47 47 47 49 49 49 45 45 45 44 44 44 44 44 44 42 42 42 44 44 44 43 43 43 45 45 45 47 47 47 49 49 49 40 40 40 11 11 11 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 2f 2f 2f 37 37 37 35 35 35 3a 3a 3a 39 39 39 39 39 39 3b 3b 3b 3d 3d 3d 3f 3f 3f 3f 3f 3f 42 42 42 47 47 47 4a 4a 4a 4c 4c 4c 49 49 49 4c 4c 4c 50 50 50 51 51 51 4f 4f 4f 37 37 37 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 3e 3e 3e 45 45 45 42 42 42 46 46 46 46 46 46 46 46 46 44 44 44 42 42 42 44 44 44 42 42 42 41 41 41 42 42 42 43 43 43 44 44 44 48 48 48 49 49 49 29 29 29 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1a 1a 1a 37 37 37 36 36 36 38 38 38 39 39 39 39 39 39 3a 3a 3a 3e 3e 3e 3f 3f 3f 41 41 41 41 41 41 43 43 43 47 47 47 48 48 48 49 49 49 49 49 49 4d 4d 4d 4d 4d 4d 4b 4b 4b 39 39 39 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 34 34 34 40 40 40 43 43 43 45 45 45 47 47 47 47 47 47 42 42 42 42 42 42 41 41 41 41 41 41 40 40 40 42 42 42 43 43 43 46 46 46 4a 4a 4a 3d 3d 3d 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 2b 2b 2b 39 39 39 3b 3b 3b 3a 3a 3a 3b 3b 3b 3c 3c 3c 40 40 40 41 41 41 3f 3f 3f 3d 3d 3d 40 40 40 40 40 40 42 42 42 44 44 44 45 45 45 49 49 49 49 49 49 48 48 48 3a 3a 3a 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2b 2b 2b 40 40 40 44 44 44 49 49 49 48 48 48 46 46 46 3f 3f 3f 40 40 40 41 41 41 41 41 41 3f 3f 3f 41 41 41 43 43 43 45 45 45 42 42 42 1a 1a 1a 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 10 10 10 34 34 34 3b 3b 3b 3b 3b 3b 3b 3b 3b 3c 3c 3c 3e 3e 3e 40 40 40 3d 3d 3d 3c 3c 3c 3e 3e 3e 3e 3e 3e 40 40 40 41 41 41 43 43 43 44 44 44 45 45 45 43 43 43 38 38 38 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2b 2b 2b 44 44 44 4b 4b 4b 4b 4b 4b 45 45 45 40 40 40 41 41 41 3f 3f 3f 3f 3f 3f 3e 3e 3e 3d 3d 3d 41 41 41 43 43 43 49 49 49 27 27 27 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1b 1b 1b 3c 3c 3c 3b 3b 3b 3c 3c 3c 3c 3c 3c 3c 3c 3c 3e 3e 3e 3c 3c 3c 3c 3c 3c 3f 3f 3f 3b 3b 3b 3e 3e 3e 40 40 40 43 43 43 45 45 45 47 47 47 42 42 42 3b 3b 3b 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 29 29 29 45 45 45 49 49 49 44 44 44 41 41 41 3e 3e 3e 41 41 41 3f 3f 3f 3d 3d 3d 3e 3e 3e 3d 3d 3d 3e 3e 3e 40 40 40 26 26 26 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 26 26 26 3a 3a 3a 3c 3c 3c 39 39 39 3b 3b 3b 3d 3d 3d 3b 3b 3b 3c 3c 3c 3d 3d 3d 3d 3d 3d 3e 3e 3e 3f 3f 3f 43 43 43 43 43 43 46 46 46 42 42 42 3c 3c 3c 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 26 26 26 43 43 43 41 41 41 42 42 42 42 42 42 3e 3e 3e 41 41 41 40 40 40 3e 3e 3e 3d 3d 3d 3e 3e 3e 3e 3e 3e 20 20 20 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 23 23 23 39 39 39 3a 3a 3a 3d 3d 3d 3c 3c 3c 3b 3b 3b 3a 3a 3a 3d 3d 3d 3b 3b 3b 3e 3e 3e 40 40 40 42 42 42 44 44 44 44 44 44 41 41 41 3d 3d 3d 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 23 23 23 48 48 48 4b 4b 4b 4f 4f 4f 51 51 51 4d 4d 4d 4a 4a 4a 45 45 45 41 41 41 3b 3b 3b 2d 2d 2d 14 14 14 04 04 04 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1b 1b 1b 35 35 35 3d 3d 3d 3c 3c 3c 3c 3c 3c 3c 3c 3c 3f 3f 3f 40 40 40 40 40 40 42 42 42 42 42 42 44 44 44 46 46 46 42 42 42 3d 3d 3d 06 06 06 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 33 33 33 74 74 74 77 77 77 7c 7c 7c 7c 7c 7c 7b 7b 7b 77 77 77 69 69 69 50 50 50 1f 1f 1f 06 06 06 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 14 14 14 37 37 37 42 42 42 48 48 48 47 47 47 4b 4b 4b 4d 4d 4d 51 51 51 55 55 55 55 55 55 57 57 57 5a 5a 5a 59 59 59 56 56 56 09 09 09 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2c 2c 2c 6a 6a 6a 6c 6c 6c 6e 6e 6e 6a 6a 6a 63 63 63 54 54 54 33 33 33 10 10 10 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 10 10 10 3d 3d 3d 60 60 60 6c 6c 6c 72 72 72 74 74 74 76 76 76 74 74 74 74 74 74 72 72 72 6d 6d 6d 68 68 68 5f 5f 5f 0b 0b 0b 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 1f 1f 1f 4f 4f 4f 4b 4b 4b 41 41 41 30 30 30 1e 1e 1e 0c 0c 0c 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 0a 0a 0a 29 29 29 4a 4a 4a 5e 5e 5e 60 60 60 5c 5c 5c 54 54 54 58 58 58 59 59 59 58 58 58 52 52 52 4a 4a 4a 0b 0b 0b 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 08 08 08 13 13 13 0b 0b 0b 06 06 06 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 16 16 16 1f 1f 1f 1e 1e 1e 10 10 10 21 21 21 22 22 22 1d 1d 1d 16 16 16 10 10 10 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
