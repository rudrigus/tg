  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 04 04 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 06 13 20 22 1a 13 0b 0f 10 13 06 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 06 1b 30 41 3a 38 34 31 3b 3d 3b 24 1b 19 15 0f 04 03 03 02 03 03 05 09 0b 0a 0b 0c 0e 1a 22 25 21 22 22 16 04 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 04 17 2e 4b 4d 3e 3b 38 3b 4f 56 55 4f 30 2d 29 24 05 03 03 02 03 03 0e 2a 27 27 28 2a 2a 2f 42 5d 67 62 5f 5a 34 07 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 0e 28 3a 48 3f 3c 38 39 3c 4f 5b 5a 5c 3b 31 2c 26 05 03 03 02 03 03 14 31 2f 2f 2e 2f 32 34 36 3e 5a 71 75 72 65 2c 05 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 06 1f 31 3e 3d 3c 3b 38 3f 3f 4a 52 51 55 3b 32 2f 26 04 03 03 02 03 03 18 31 32 32 32 31 31 34 36 37 3a 45 60 70 6c 46 19 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 13 2a 3a 3e 3e 3c 3b 3b 3d 3e 48 49 42 44 37 31 31 26 04 03 03 02 03 03 1b 33 34 32 32 32 35 38 38 3b 3a 3a 3d 41 42 41 34 0c 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 07 22 34 3e 40 43 3a 3d 3e 3f 40 42 3e 3b 39 35 34 33 22 04 03 03 02 03 03 21 35 35 35 34 35 35 37 38 3a 3b 3a 3c 3a 39 3e 42 24 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 04 11 2a 3b 43 40 40 3a 3d 40 3f 41 40 3e 3b 38 38 35 32 1e 03 03 03 02 03 03 25 37 37 36 37 38 36 3b 3c 3d 3e 3f 3d 3b 3a 3f 43 3a 0b 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 05 1d 37 40 46 41 3f 3e 3e 40 3f 3f 3f 3a 3a 37 38 34 30 1a 03 03 03 02 03 03 26 36 38 39 39 39 38 3e 3e 3e 42 41 3f 3c 3e 41 45 44 23 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 0a 29 41 40 42 41 46 3e 41 42 40 3f 3f 3c 3b 38 36 34 2f 1a 03 03 03 02 03 03 2c 38 3c 3d 3d 3d 3d 41 42 44 44 43 44 40 41 43 46 45 39 08 03 03 03 02 03 03
  03 02 03 03 03 03 03 04 11 35 46 41 46 45 4a 44 46 44 42 3e 3f 3d 3b 39 36 35 31 1a 03 03 03 02 03 03 31 39 3d 3f 40 40 41 40 46 47 48 46 46 44 44 45 49 48 42 18 03 03 03 02 03 03
  03 02 03 03 03 03 03 05 1e 42 49 40 41 41 41 40 43 43 44 41 40 3f 3d 3b 37 37 32 18 03 03 03 02 03 04 36 3e 3f 40 3e 40 41 40 45 47 48 47 49 47 48 49 4a 49 45 2a 05 03 03 02 03 03
  03 02 03 03 03 03 03 09 2f 44 46 3f 42 41 40 42 43 44 42 41 41 3d 3b 39 38 37 33 16 03 03 03 02 03 06 3a 42 42 41 42 3f 40 40 42 47 47 47 48 48 4a 4b 4f 4f 4a 39 0d 03 03 02 03 03
  03 02 03 03 03 03 03 11 37 46 44 41 45 43 43 42 42 41 44 42 40 3d 3a 39 3b 38 35 14 03 03 03 02 03 08 49 4a 46 45 48 48 46 45 44 46 48 47 49 49 4b 4c 51 51 4f 3f 1e 03 03 02 03 03
  03 02 03 03 03 03 05 17 43 46 41 41 43 43 42 43 42 42 42 41 41 3d 3b 39 3b 39 36 12 03 03 03 02 03 0c 4d 57 54 55 53 54 4c 4c 46 47 48 49 49 4a 4c 4d 52 58 4d 45 2a 06 03 02 03 03
  03 02 03 03 03 03 07 1f 4a 46 44 43 46 45 44 44 43 42 45 43 40 3d 3c 3b 3e 3f 3c 13 03 03 03 02 03 11 4d 4e 4f 52 51 57 58 53 4f 4e 4d 4b 4c 4b 4f 53 5c 59 53 4b 38 0d 03 02 03 03
  03 02 03 03 03 03 0b 29 4f 49 47 47 47 45 46 44 44 44 45 43 43 41 43 47 47 45 46 15 03 03 03 02 03 17 50 4f 53 59 5e 5a 56 53 53 53 53 4e 4c 4c 58 77 7d 64 5a 4d 46 1b 03 02 03 03
  03 02 03 03 03 03 0b 3d 55 49 49 4a 4c 4a 48 45 45 47 46 44 46 4c 51 4b 49 49 46 12 03 03 03 02 03 1f 54 56 5a 62 6b 5d 56 56 58 5d 5c 56 50 4d 67 8f 85 6b 5f 4f 47 2d 07 03 03 03
  03 02 03 03 03 03 12 65 56 4d 4c 4f 4f 51 51 50 52 52 4f 4e 52 53 54 54 52 51 4d 10 03 03 03 02 03 25 5b 5d 5d 60 60 5d 5b 59 57 56 57 5f 57 57 62 71 67 61 5e 4f 49 39 12 02 03 03
  03 02 03 03 03 04 2b 78 55 51 52 53 5c 63 61 60 60 5d 5c 59 5a 59 59 5b 5a 59 53 0e 03 03 03 02 03 2e 63 60 62 62 62 61 5e 5c 5b 58 53 5b 5c 60 63 60 5c 5d 52 4a 46 40 2b 04 03 03
  03 02 03 03 03 06 43 7a 54 53 58 63 67 67 69 6d 72 74 74 6f 6f 6d 6d 6a 6c 6a 63 0d 03 03 03 02 03 44 7a 77 7b 7d 77 68 64 61 5e 5a 55 53 58 5d 63 63 57 5c 5d 4d 44 45 4b 09 03 03
  03 02 03 03 03 0b 4f 7f 58 5a 68 65 6a 79 84 86 86 8a 8f 91 8e 8e 8c 8c 8f 8c 7e 0b 03 03 03 02 03 56 84 7b 7d 7b 7b 72 6d 66 62 5f 5d 56 54 5d 69 70 62 5b 66 50 45 4c 52 12 03 03
  03 02 03 03 03 0e 4f 87 65 66 67 6c 84 8b 84 83 83 88 8a 8d 95 95 8f 8a 86 83 72 08 03 03 03 03 04 57 73 73 76 75 77 76 72 6d 68 64 60 5e 5d 57 5a 65 62 59 59 51 44 5a 56 14 03 03
  03 02 03 03 03 0e 4e 92 76 6b 70 7b 84 83 80 82 84 86 8d 92 9c 9d 96 8c 8b 89 78 07 03 03 03 03 07 63 78 79 7b 7e 7f 7e 7c 76 6d 6a 66 61 63 60 5c 63 64 5b 58 50 4a 6c 53 11 03 03
  03 02 03 03 03 0d 4b 95 76 72 7f 85 88 87 88 8a 8c 92 99 a1 ab a7 a1 9a 9f a2 80 05 04 03 03 04 0a 71 80 81 82 85 87 85 81 7a 76 72 6b 66 65 67 61 62 67 62 5d 53 50 70 52 11 03 03
  03 02 03 03 03 0a 44 93 76 7d 89 88 8d 91 92 93 96 99 9f ac b6 b3 b0 ac b7 bf 84 06 04 03 03 06 11 7b 8e 89 8b 8b 8e 8b 83 7e 79 76 6f 6b 68 67 6c 63 65 6d 65 59 57 72 4a 0c 03 03
  03 02 03 03 03 09 3b 91 7b 83 8a 89 92 98 9c 9f a0 a3 a3 ab b6 b9 b6 b4 bc c8 84 0a 06 04 03 08 1d 7d 95 98 95 96 98 90 89 83 7f 7d 77 71 6d 6b 70 70 69 6b 6d 6b 61 70 3f 09 03 03
  03 02 03 03 03 06 2d 85 81 86 8c 90 9a a0 a3 a5 a7 a8 ac aa b0 b3 b6 b3 b3 c2 85 17 0f 0a 0c 16 34 a5 ab 98 98 9f 9d 95 8e 88 87 85 81 7b 77 75 74 79 77 6f 6a 70 69 67 2d 05 03 03
  03 02 03 03 03 04 1d 75 7f 81 91 93 97 9f a3 a7 a8 ab ab a6 ad b1 b1 af ad b3 9d 3a 24 1f 23 30 58 c9 e1 a5 96 a7 a3 9a 96 91 90 8e 8a 89 85 80 7e 7c 7b 79 71 6d 70 5a 16 04 03 03
  03 02 03 03 03 03 0f 62 78 7f 8a 86 8c 94 9a a0 a4 a9 ab a8 a8 aa b7 a8 a6 ab bc 71 52 41 49 6b 81 d5 ea b3 97 a7 aa a2 9a 9a 97 96 97 97 93 8a 87 82 7b 7b 77 6e 69 49 09 03 03 03
  03 02 03 03 03 03 0a 59 77 7b 78 73 7d 86 8b 92 a2 aa ad ac aa a8 b2 ae a8 ac c9 c3 8f 7a 75 9b d2 fc df ae 9f a9 ad a7 a2 a2 a1 a1 a2 a4 a3 99 92 87 7f 78 76 6f 63 34 05 02 03 03
  03 02 03 03 03 03 0a 5f 7d 6f 69 6b 74 79 7e 88 9c ae b2 b1 b0 b0 bf c2 be c2 dc f9 ec de da f5 fe fb dc bb b8 b2 b3 b2 b0 ad aa ad ad b1 b1 a6 9d 90 83 7c 70 6d 6a 3b 03 03 03 03
  03 02 03 03 03 03 0b 64 88 69 68 6d 72 77 7b 88 a1 b5 bb b9 b7 c0 d4 d1 d5 dd e6 f1 fb ff ff ff ff fb e7 e7 e8 df d5 cd c4 b9 b9 ba b8 bc b3 a8 9e 91 7e 7a 73 6a 73 52 04 02 03 03
  03 02 03 03 03 03 07 47 93 6c 70 74 75 7d 84 99 b3 c6 d1 cd c8 cd d8 de de dc dc dd f4 ff ff ff ff ff fe fd fe fd fa f1 dc c9 c6 c5 c2 bd b6 a7 99 8f 83 73 6e 6a 7b 5c 07 02 03 03
  03 02 03 03 03 03 04 26 7f 89 76 79 7b 7c 84 92 aa ca d6 cf ca cf da de e3 e2 dd da eb fe ff ff ff ff ff fb f7 f5 ef eb e3 da d1 ce cb c8 c4 b5 a7 98 8d 7f 70 72 97 60 09 03 03 03
  03 02 03 03 03 03 03 0b 49 7d 72 78 7d 7b 7a 81 94 ab ac a0 a5 bb d2 e4 ee ea de db ea fe ff ff ff ff ff fe fc fa fa f5 f1 e8 e4 e0 dd de dc d3 c5 b4 9f 92 87 7d 9e 49 09 03 03 03
  03 02 03 03 03 03 03 04 1c 5b 61 77 86 8d 87 8e 94 90 90 8c 94 a5 bf d6 ee e8 dc de f5 ff ff ff ff ff ff ff fd fa f5 ea ea ea e9 e5 e7 eb ee e6 dc ce b6 a3 95 86 84 2c 04 02 03 03
  03 02 03 03 03 03 03 03 07 31 58 6b 84 92 96 96 9a 92 98 8e 91 9d b2 ce e3 e3 e1 ea fc ff ff ff ff ff ff ff ff f7 ea da d2 d5 db d9 df e3 ec ed ee ef e0 c7 a2 9e 70 1b 03 02 03 03
  03 02 03 03 03 03 03 03 04 10 44 76 7d 87 8a 91 9d 9e 9f 9a 92 9b b3 cd df e7 ee f9 ff ff ff ff ff fd fc fe ff fa e8 d7 c9 c7 d0 e7 f4 f1 f7 ef e8 f0 d6 ba bf af 3a 07 03 02 03 03
  03 02 03 03 03 03 03 03 03 04 22 67 7b 6d 6b 79 97 a0 a5 a3 9e a2 b6 ce e1 eb f7 fc fe ff ff fe f5 dd e0 f3 fe fe ec d5 cd d2 f5 fc f2 df f0 d8 d7 c5 a2 a2 ae 3f 0f 04 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 04 14 35 57 59 5e 6a 6d 85 98 a8 a7 b3 bf c7 d2 e6 ca c2 d9 e7 de c0 b8 b1 cb e7 e4 e4 d1 c7 ea fe f9 e9 e9 cd b3 ae 9f 82 90 48 0c 04 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 08 19 2d 3c 49 5d 66 7a 94 93 92 98 9a ad b3 9c 8f 93 a4 9f 9c aa a2 9c a6 a1 a2 9f a6 c6 f9 f6 ef ce a2 8f 87 69 4e 34 0a 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 07 18 2a 46 53 6f 76 75 7c 7f 77 79 78 76 7d 8a 98 99 a0 96 8f 85 7a 78 83 87 96 a8 c5 d0 cb ba 87 6f 52 31 14 04 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 04 0f 23 25 23 3a 48 56 64 67 6d 6e 6d 71 79 7a 7c 83 81 78 6e 68 5d 6b 72 8a a7 93 a8 bc 9b 6d 2a 10 06 04 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 04 06 05 0a 13 16 1f 2c 3b 48 4b 4d 57 5f 62 64 64 5c 52 4a 43 48 3e 41 45 3b 31 23 18 0d 05 03 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 03 03 03 03 04 05 0a 0c 12 21 30 2b 37 42 39 2c 27 1f 1c 16 14 0f 0e 0b 07 07 07 05 05 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 04 03 05 07 0d 10 0d 0e 0c 0a 06 04 06 03 03 03 05 03 03 04 03 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 03 03 03 03 02 03 03 03 02 03 03 03 03 03 03 03 03 02 03 03
  