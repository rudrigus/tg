-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "11/18/2015 21:55:21"
                                                            
-- Vhdl Test Bench template for design  :  ProcessadorImagemGMAW
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;
--use work.imagensteste.all;

ENTITY ProcessadorImagemGMAW_TB IS
END ProcessadorImagemGMAW_TB;
ARCHITECTURE ProcessadorImagemGMAW_arch OF ProcessadorImagemGMAW_TB IS
-- constants                                                 

  constant imagem_teste0 : MatrizImagem :=  ((X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"13", X"20", X"22", X"1a", X"13", X"0b", X"0f", X"10", X"13", X"06", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"1b", X"30", X"41", X"3a", X"38", X"34", X"31", X"3b", X"3d", X"3b", X"24", X"1b", X"19", X"15", X"0f", X"04", X"03", X"03", X"02", X"03", X"03", X"05", X"09", X"0b", X"0a", X"0b", X"0c", X"0e", X"1a", X"22", X"25", X"21", X"22", X"22", X"16", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"17", X"2e", X"4b", X"4d", X"3e", X"3b", X"38", X"3b", X"4f", X"56", X"55", X"4f", X"30", X"2d", X"29", X"24", X"05", X"03", X"03", X"02", X"03", X"03", X"0e", X"2a", X"27", X"27", X"28", X"2a", X"2a", X"2f", X"42", X"5d", X"67", X"62", X"5f", X"5a", X"34", X"07", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0e", X"28", X"3a", X"48", X"3f", X"3c", X"38", X"39", X"3c", X"4f", X"5b", X"5a", X"5c", X"3b", X"31", X"2c", X"26", X"05", X"03", X"03", X"02", X"03", X"03", X"14", X"31", X"2f", X"2f", X"2e", X"2f", X"32", X"34", X"36", X"3e", X"5a", X"71", X"75", X"72", X"65", X"2c", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"1f", X"31", X"3e", X"3d", X"3c", X"3b", X"38", X"3f", X"3f", X"4a", X"52", X"51", X"55", X"3b", X"32", X"2f", X"26", X"04", X"03", X"03", X"02", X"03", X"03", X"18", X"31", X"32", X"32", X"32", X"31", X"31", X"34", X"36", X"37", X"3a", X"45", X"60", X"70", X"6c", X"46", X"19", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"13", X"2a", X"3a", X"3e", X"3e", X"3c", X"3b", X"3b", X"3d", X"3e", X"48", X"49", X"42", X"44", X"37", X"31", X"31", X"26", X"04", X"03", X"03", X"02", X"03", X"03", X"1b", X"33", X"34", X"32", X"32", X"32", X"35", X"38", X"38", X"3b", X"3a", X"3a", X"3d", X"41", X"42", X"41", X"34", X"0c", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"22", X"34", X"3e", X"40", X"43", X"3a", X"3d", X"3e", X"3f", X"40", X"42", X"3e", X"3b", X"39", X"35", X"34", X"33", X"22", X"04", X"03", X"03", X"02", X"03", X"03", X"21", X"35", X"35", X"35", X"34", X"35", X"35", X"37", X"38", X"3a", X"3b", X"3a", X"3c", X"3a", X"39", X"3e", X"42", X"24", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"11", X"2a", X"3b", X"43", X"40", X"40", X"3a", X"3d", X"40", X"3f", X"41", X"40", X"3e", X"3b", X"38", X"38", X"35", X"32", X"1e", X"03", X"03", X"03", X"02", X"03", X"03", X"25", X"37", X"37", X"36", X"37", X"38", X"36", X"3b", X"3c", X"3d", X"3e", X"3f", X"3d", X"3b", X"3a", X"3f", X"43", X"3a", X"0b", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"05", X"1d", X"37", X"40", X"46", X"41", X"3f", X"3e", X"3e", X"40", X"3f", X"3f", X"3f", X"3a", X"3a", X"37", X"38", X"34", X"30", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"26", X"36", X"38", X"39", X"39", X"39", X"38", X"3e", X"3e", X"3e", X"42", X"41", X"3f", X"3c", X"3e", X"41", X"45", X"44", X"23", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0a", X"29", X"41", X"40", X"42", X"41", X"46", X"3e", X"41", X"42", X"40", X"3f", X"3f", X"3c", X"3b", X"38", X"36", X"34", X"2f", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"2c", X"38", X"3c", X"3d", X"3d", X"3d", X"3d", X"41", X"42", X"44", X"44", X"43", X"44", X"40", X"41", X"43", X"46", X"45", X"39", X"08", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"11", X"35", X"46", X"41", X"46", X"45", X"4a", X"44", X"46", X"44", X"42", X"3e", X"3f", X"3d", X"3b", X"39", X"36", X"35", X"31", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"31", X"39", X"3d", X"3f", X"40", X"40", X"41", X"40", X"46", X"47", X"48", X"46", X"46", X"44", X"44", X"45", X"49", X"48", X"42", X"18", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"05", X"1e", X"42", X"49", X"40", X"41", X"41", X"41", X"40", X"43", X"43", X"44", X"41", X"40", X"3f", X"3d", X"3b", X"37", X"37", X"32", X"18", X"03", X"03", X"03", X"02", X"03", X"04", X"36", X"3e", X"3f", X"40", X"3e", X"40", X"41", X"40", X"45", X"47", X"48", X"47", X"49", X"47", X"48", X"49", X"4a", X"49", X"45", X"2a", X"05", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"09", X"2f", X"44", X"46", X"3f", X"42", X"41", X"40", X"42", X"43", X"44", X"42", X"41", X"41", X"3d", X"3b", X"39", X"38", X"37", X"33", X"16", X"03", X"03", X"03", X"02", X"03", X"06", X"3a", X"42", X"42", X"41", X"42", X"3f", X"40", X"40", X"42", X"47", X"47", X"47", X"48", X"48", X"4a", X"4b", X"4f", X"4f", X"4a", X"39", X"0d", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"11", X"37", X"46", X"44", X"41", X"45", X"43", X"43", X"42", X"42", X"41", X"44", X"42", X"40", X"3d", X"3a", X"39", X"3b", X"38", X"35", X"14", X"03", X"03", X"03", X"02", X"03", X"08", X"49", X"4a", X"46", X"45", X"48", X"48", X"46", X"45", X"44", X"46", X"48", X"47", X"49", X"49", X"4b", X"4c", X"51", X"51", X"4f", X"3f", X"1e", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"17", X"43", X"46", X"41", X"41", X"43", X"43", X"42", X"43", X"42", X"42", X"42", X"41", X"41", X"3d", X"3b", X"39", X"3b", X"39", X"36", X"12", X"03", X"03", X"03", X"02", X"03", X"0c", X"4d", X"57", X"54", X"55", X"53", X"54", X"4c", X"4c", X"46", X"47", X"48", X"49", X"49", X"4a", X"4c", X"4d", X"52", X"58", X"4d", X"45", X"2a", X"06", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"07", X"1f", X"4a", X"46", X"44", X"43", X"46", X"45", X"44", X"44", X"43", X"42", X"45", X"43", X"40", X"3d", X"3c", X"3b", X"3e", X"3f", X"3c", X"13", X"03", X"03", X"03", X"02", X"03", X"11", X"4d", X"4e", X"4f", X"52", X"51", X"57", X"58", X"53", X"4f", X"4e", X"4d", X"4b", X"4c", X"4b", X"4f", X"53", X"5c", X"59", X"53", X"4b", X"38", X"0d", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"29", X"4f", X"49", X"47", X"47", X"47", X"45", X"46", X"44", X"44", X"44", X"45", X"43", X"43", X"41", X"43", X"47", X"47", X"45", X"46", X"15", X"03", X"03", X"03", X"02", X"03", X"17", X"50", X"4f", X"53", X"59", X"5e", X"5a", X"56", X"53", X"53", X"53", X"53", X"4e", X"4c", X"4c", X"58", X"77", X"7d", X"64", X"5a", X"4d", X"46", X"1b", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"3d", X"55", X"49", X"49", X"4a", X"4c", X"4a", X"48", X"45", X"45", X"47", X"46", X"44", X"46", X"4c", X"51", X"4b", X"49", X"49", X"46", X"12", X"03", X"03", X"03", X"02", X"03", X"1f", X"54", X"56", X"5a", X"62", X"6b", X"5d", X"56", X"56", X"58", X"5d", X"5c", X"56", X"50", X"4d", X"67", X"8f", X"85", X"6b", X"5f", X"4f", X"47", X"2d", X"07", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"12", X"65", X"56", X"4d", X"4c", X"4f", X"4f", X"51", X"51", X"50", X"52", X"52", X"4f", X"4e", X"52", X"53", X"54", X"54", X"52", X"51", X"4d", X"10", X"03", X"03", X"03", X"02", X"03", X"25", X"5b", X"5d", X"5d", X"60", X"60", X"5d", X"5b", X"59", X"57", X"56", X"57", X"5f", X"57", X"57", X"62", X"71", X"67", X"61", X"5e", X"4f", X"49", X"39", X"12", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"2b", X"78", X"55", X"51", X"52", X"53", X"5c", X"63", X"61", X"60", X"60", X"5d", X"5c", X"59", X"5a", X"59", X"59", X"5b", X"5a", X"59", X"53", X"0e", X"03", X"03", X"03", X"02", X"03", X"2e", X"63", X"60", X"62", X"62", X"62", X"61", X"5e", X"5c", X"5b", X"58", X"53", X"5b", X"5c", X"60", X"63", X"60", X"5c", X"5d", X"52", X"4a", X"46", X"40", X"2b", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"06", X"43", X"7a", X"54", X"53", X"58", X"63", X"67", X"67", X"69", X"6d", X"72", X"74", X"74", X"6f", X"6f", X"6d", X"6d", X"6a", X"6c", X"6a", X"63", X"0d", X"03", X"03", X"03", X"02", X"03", X"44", X"7a", X"77", X"7b", X"7d", X"77", X"68", X"64", X"61", X"5e", X"5a", X"55", X"53", X"58", X"5d", X"63", X"63", X"57", X"5c", X"5d", X"4d", X"44", X"45", X"4b", X"09", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0b", X"4f", X"7f", X"58", X"5a", X"68", X"65", X"6a", X"79", X"84", X"86", X"86", X"8a", X"8f", X"91", X"8e", X"8e", X"8c", X"8c", X"8f", X"8c", X"7e", X"0b", X"03", X"03", X"03", X"02", X"03", X"56", X"84", X"7b", X"7d", X"7b", X"7b", X"72", X"6d", X"66", X"62", X"5f", X"5d", X"56", X"54", X"5d", X"69", X"70", X"62", X"5b", X"66", X"50", X"45", X"4c", X"52", X"12", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0e", X"4f", X"87", X"65", X"66", X"67", X"6c", X"84", X"8b", X"84", X"83", X"83", X"88", X"8a", X"8d", X"95", X"95", X"8f", X"8a", X"86", X"83", X"72", X"08", X"03", X"03", X"03", X"03", X"04", X"57", X"73", X"73", X"76", X"75", X"77", X"76", X"72", X"6d", X"68", X"64", X"60", X"5e", X"5d", X"57", X"5a", X"65", X"62", X"59", X"59", X"51", X"44", X"5a", X"56", X"14", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0e", X"4e", X"92", X"76", X"6b", X"70", X"7b", X"84", X"83", X"80", X"82", X"84", X"86", X"8d", X"92", X"9c", X"9d", X"96", X"8c", X"8b", X"89", X"78", X"07", X"03", X"03", X"03", X"03", X"07", X"63", X"78", X"79", X"7b", X"7e", X"7f", X"7e", X"7c", X"76", X"6d", X"6a", X"66", X"61", X"63", X"60", X"5c", X"63", X"64", X"5b", X"58", X"50", X"4a", X"6c", X"53", X"11", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0d", X"4b", X"95", X"76", X"72", X"7f", X"85", X"88", X"87", X"88", X"8a", X"8c", X"92", X"99", X"a1", X"ab", X"a7", X"a1", X"9a", X"9f", X"a2", X"80", X"05", X"04", X"03", X"03", X"04", X"0a", X"71", X"80", X"81", X"82", X"85", X"87", X"85", X"81", X"7a", X"76", X"72", X"6b", X"66", X"65", X"67", X"61", X"62", X"67", X"62", X"5d", X"53", X"50", X"70", X"52", X"11", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0a", X"44", X"93", X"76", X"7d", X"89", X"88", X"8d", X"91", X"92", X"93", X"96", X"99", X"9f", X"ac", X"b6", X"b3", X"b0", X"ac", X"b7", X"bf", X"84", X"06", X"04", X"03", X"03", X"06", X"11", X"7b", X"8e", X"89", X"8b", X"8b", X"8e", X"8b", X"83", X"7e", X"79", X"76", X"6f", X"6b", X"68", X"67", X"6c", X"63", X"65", X"6d", X"65", X"59", X"57", X"72", X"4a", X"0c", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"09", X"3b", X"91", X"7b", X"83", X"8a", X"89", X"92", X"98", X"9c", X"9f", X"a0", X"a3", X"a3", X"ab", X"b6", X"b9", X"b6", X"b4", X"bc", X"c8", X"84", X"0a", X"06", X"04", X"03", X"08", X"1d", X"7d", X"95", X"98", X"95", X"96", X"98", X"90", X"89", X"83", X"7f", X"7d", X"77", X"71", X"6d", X"6b", X"70", X"70", X"69", X"6b", X"6d", X"6b", X"61", X"70", X"3f", X"09", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"06", X"2d", X"85", X"81", X"86", X"8c", X"90", X"9a", X"a0", X"a3", X"a5", X"a7", X"a8", X"ac", X"aa", X"b0", X"b3", X"b6", X"b3", X"b3", X"c2", X"85", X"17", X"0f", X"0a", X"0c", X"16", X"34", X"a5", X"ab", X"98", X"98", X"9f", X"9d", X"95", X"8e", X"88", X"87", X"85", X"81", X"7b", X"77", X"75", X"74", X"79", X"77", X"6f", X"6a", X"70", X"69", X"67", X"2d", X"05", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"1d", X"75", X"7f", X"81", X"91", X"93", X"97", X"9f", X"a3", X"a7", X"a8", X"ab", X"ab", X"a6", X"ad", X"b1", X"b1", X"af", X"ad", X"b3", X"9d", X"3a", X"24", X"1f", X"23", X"30", X"58", X"c9", X"e1", X"a5", X"96", X"a7", X"a3", X"9a", X"96", X"91", X"90", X"8e", X"8a", X"89", X"85", X"80", X"7e", X"7c", X"7b", X"79", X"71", X"6d", X"70", X"5a", X"16", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0f", X"62", X"78", X"7f", X"8a", X"86", X"8c", X"94", X"9a", X"a0", X"a4", X"a9", X"ab", X"a8", X"a8", X"aa", X"b7", X"a8", X"a6", X"ab", X"bc", X"71", X"52", X"41", X"49", X"6b", X"81", X"d5", X"ea", X"b3", X"97", X"a7", X"aa", X"a2", X"9a", X"9a", X"97", X"96", X"97", X"97", X"93", X"8a", X"87", X"82", X"7b", X"7b", X"77", X"6e", X"69", X"49", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0a", X"59", X"77", X"7b", X"78", X"73", X"7d", X"86", X"8b", X"92", X"a2", X"aa", X"ad", X"ac", X"aa", X"a8", X"b2", X"ae", X"a8", X"ac", X"c9", X"c3", X"8f", X"7a", X"75", X"9b", X"d2", X"fc", X"df", X"ae", X"9f", X"a9", X"ad", X"a7", X"a2", X"a2", X"a1", X"a1", X"a2", X"a4", X"a3", X"99", X"92", X"87", X"7f", X"78", X"76", X"6f", X"63", X"34", X"05", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0a", X"5f", X"7d", X"6f", X"69", X"6b", X"74", X"79", X"7e", X"88", X"9c", X"ae", X"b2", X"b1", X"b0", X"b0", X"bf", X"c2", X"be", X"c2", X"dc", X"f9", X"ec", X"de", X"da", X"f5", X"fe", X"fb", X"dc", X"bb", X"b8", X"b2", X"b3", X"b2", X"b0", X"ad", X"aa", X"ad", X"ad", X"b1", X"b1", X"a6", X"9d", X"90", X"83", X"7c", X"70", X"6d", X"6a", X"3b", X"03", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"64", X"88", X"69", X"68", X"6d", X"72", X"77", X"7b", X"88", X"a1", X"b5", X"bb", X"b9", X"b7", X"c0", X"d4", X"d1", X"d5", X"dd", X"e6", X"f1", X"fb", X"ff", X"ff", X"ff", X"ff", X"fb", X"e7", X"e7", X"e8", X"df", X"d5", X"cd", X"c4", X"b9", X"b9", X"ba", X"b8", X"bc", X"b3", X"a8", X"9e", X"91", X"7e", X"7a", X"73", X"6a", X"73", X"52", X"04", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"07", X"47", X"93", X"6c", X"70", X"74", X"75", X"7d", X"84", X"99", X"b3", X"c6", X"d1", X"cd", X"c8", X"cd", X"d8", X"de", X"de", X"dc", X"dc", X"dd", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fd", X"fe", X"fd", X"fa", X"f1", X"dc", X"c9", X"c6", X"c5", X"c2", X"bd", X"b6", X"a7", X"99", X"8f", X"83", X"73", X"6e", X"6a", X"7b", X"5c", X"07", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"26", X"7f", X"89", X"76", X"79", X"7b", X"7c", X"84", X"92", X"aa", X"ca", X"d6", X"cf", X"ca", X"cf", X"da", X"de", X"e3", X"e2", X"dd", X"da", X"eb", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f7", X"f5", X"ef", X"eb", X"e3", X"da", X"d1", X"ce", X"cb", X"c8", X"c4", X"b5", X"a7", X"98", X"8d", X"7f", X"70", X"72", X"97", X"60", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"0b", X"49", X"7d", X"72", X"78", X"7d", X"7b", X"7a", X"81", X"94", X"ab", X"ac", X"a0", X"a5", X"bb", X"d2", X"e4", X"ee", X"ea", X"de", X"db", X"ea", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fc", X"fa", X"fa", X"f5", X"f1", X"e8", X"e4", X"e0", X"dd", X"de", X"dc", X"d3", X"c5", X"b4", X"9f", X"92", X"87", X"7d", X"9e", X"49", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"1c", X"5b", X"61", X"77", X"86", X"8d", X"87", X"8e", X"94", X"90", X"90", X"8c", X"94", X"a5", X"bf", X"d6", X"ee", X"e8", X"dc", X"de", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fa", X"f5", X"ea", X"ea", X"ea", X"e9", X"e5", X"e7", X"eb", X"ee", X"e6", X"dc", X"ce", X"b6", X"a3", X"95", X"86", X"84", X"2c", X"04", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"31", X"58", X"6b", X"84", X"92", X"96", X"96", X"9a", X"92", X"98", X"8e", X"91", X"9d", X"b2", X"ce", X"e3", X"e3", X"e1", X"ea", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"ea", X"da", X"d2", X"d5", X"db", X"d9", X"df", X"e3", X"ec", X"ed", X"ee", X"ef", X"e0", X"c7", X"a2", X"9e", X"70", X"1b", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"10", X"44", X"76", X"7d", X"87", X"8a", X"91", X"9d", X"9e", X"9f", X"9a", X"92", X"9b", X"b3", X"cd", X"df", X"e7", X"ee", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fc", X"fe", X"ff", X"fa", X"e8", X"d7", X"c9", X"c7", X"d0", X"e7", X"f4", X"f1", X"f7", X"ef", X"e8", X"f0", X"d6", X"ba", X"bf", X"af", X"3a", X"07", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"22", X"67", X"7b", X"6d", X"6b", X"79", X"97", X"a0", X"a5", X"a3", X"9e", X"a2", X"b6", X"ce", X"e1", X"eb", X"f7", X"fc", X"fe", X"ff", X"ff", X"fe", X"f5", X"dd", X"e0", X"f3", X"fe", X"fe", X"ec", X"d5", X"cd", X"d2", X"f5", X"fc", X"f2", X"df", X"f0", X"d8", X"d7", X"c5", X"a2", X"a2", X"ae", X"3f", X"0f", X"04", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"14", X"35", X"57", X"59", X"5e", X"6a", X"6d", X"85", X"98", X"a8", X"a7", X"b3", X"bf", X"c7", X"d2", X"e6", X"ca", X"c2", X"d9", X"e7", X"de", X"c0", X"b8", X"b1", X"cb", X"e7", X"e4", X"e4", X"d1", X"c7", X"ea", X"fe", X"f9", X"e9", X"e9", X"cd", X"b3", X"ae", X"9f", X"82", X"90", X"48", X"0c", X"04", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"08", X"19", X"2d", X"3c", X"49", X"5d", X"66", X"7a", X"94", X"93", X"92", X"98", X"9a", X"ad", X"b3", X"9c", X"8f", X"93", X"a4", X"9f", X"9c", X"aa", X"a2", X"9c", X"a6", X"a1", X"a2", X"9f", X"a6", X"c6", X"f9", X"f6", X"ef", X"ce", X"a2", X"8f", X"87", X"69", X"4e", X"34", X"0a", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"18", X"2a", X"46", X"53", X"6f", X"76", X"75", X"7c", X"7f", X"77", X"79", X"78", X"76", X"7d", X"8a", X"98", X"99", X"a0", X"96", X"8f", X"85", X"7a", X"78", X"83", X"87", X"96", X"a8", X"c5", X"d0", X"cb", X"ba", X"87", X"6f", X"52", X"31", X"14", X"04", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"0f", X"23", X"25", X"23", X"3a", X"48", X"56", X"64", X"67", X"6d", X"6e", X"6d", X"71", X"79", X"7a", X"7c", X"83", X"81", X"78", X"6e", X"68", X"5d", X"6b", X"72", X"8a", X"a7", X"93", X"a8", X"bc", X"9b", X"6d", X"2a", X"10", X"06", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"04", X"06", X"05", X"0a", X"13", X"16", X"1f", X"2c", X"3b", X"48", X"4b", X"4d", X"57", X"5f", X"62", X"64", X"64", X"5c", X"52", X"4a", X"43", X"48", X"3e", X"41", X"45", X"3b", X"31", X"23", X"18", X"0d", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"0a", X"0c", X"12", X"21", X"30", X"2b", X"37", X"42", X"39", X"2c", X"27", X"1f", X"1c", X"16", X"14", X"0f", X"0e", X"0b", X"07", X"07", X"07", X"05", X"05", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"03", X"05", X"07", X"0d", X"10", X"0d", X"0e", X"0c", X"0a", X"06", X"04", X"06", X"03", X"03", X"03", X"05", X"03", X"03", X"04", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"));
  
  constant imagem_teste1 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

  constant imagem_teste2 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

  constant imagem_teste3 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
  (X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

-- signals                                                   
SIGNAL ENDSIM : STD_LOGIC := '0';
SIGNAL clk_count : natural := 0;
SIGNAL brilho_maximo : UNSIGNED(24 DOWNTO 0);
SIGNAL threshold1    : std_logic_vector(7 downto 0);
SIGNAL meioVert      : unsigned(7 downto 0);
SIGNAL meioImagem    : unsigned(7 downto 0);
SIGNAL in_clock : STD_LOGIC;
SIGNAL in_janela : STD_LOGIC;
SIGNAL pixel_entrada : STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
SIGNAL bloco_atual : natural range qtd_imagens downto 0 := 0;
SIGNAL linha : integer range 0 to numcols - 1 := 0;
SIGNAL coluna : integer range 0 to numlin - 1 := 0;
SIGNAL reset : STD_LOGIC;
SIGNAL start_stop :  STD_LOGIC;
SIGNAL contador12b : STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL qtd_imagens : UNSIGNED(1 DOWNTO 0) := "11";
--SIGNAL fim_imagem : STD_LOGIC := '0';
SIGNAL frequencia_camera : real := 150.000E6;


COMPONENT ProcessadorImagemGMAW
	PORT (
	brilho_maximo : IN UNSIGNED(24 DOWNTO 0);
  threshold1    : in STD_LOGIC_VECTOR(7 downto 0);
  meioVert      : in UNSIGNED(7 downto 0);
  meioImagem    : in UNSIGNED(7 downto 0);
	in_clock      : IN STD_LOGIC;
	in_janela     : IN STD_LOGIC;
	pixel_entrada : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
	);	
END COMPONENT;


-- Procedure for clock generation
  procedure clk_gen(signal clk : out std_logic; constant FREQ : real) is
    constant PERIOD    : time := 1 sec / FREQ;        -- Full period
    constant HIGH_TIME : time := PERIOD / 2;          -- High time
    constant LOW_TIME  : time := PERIOD - HIGH_TIME;  -- Low time; always >= HIGH_TIME
  begin
    -- Check the arguments
    assert (HIGH_TIME /= 0 fs) report "clk_plain: High time is zero; time resolution to large for frequency" severity FAILURE;
    -- Generate a clock cycle
    loop
      if (ENDSIM = '0') then
        clk <= '1';
        wait for HIGH_TIME;
        clk <= '0';
        wait for LOW_TIME;
      else
        wait;
      end if;
    end loop;
  end procedure;



BEGIN
  -- Clock generation with concurrent procedure call
  clk_gen(in_clock, frequencia_camera);  -- 166.667 MHz clock

  -- Time resolution show
  assert FALSE report "Time resolution: " & time'image(time'succ(0 fs)) severity NOTE;



	i1 : ProcessadorImagemGMAW
	PORT MAP (
-- list connections between master ports and signals
	brilho_maximo => brilho_maximo,
  threshold1 => threshold1,
  meioVert => meioVert,
  meioImagem => meioImagem,
	in_clock => in_clock,
	in_janela => in_janela,
	pixel_entrada => pixel_entrada
	);

brilho_maximo <= to_unsigned(720000,25) after 0 ns;
threshold1    <= "00001010" after 0 ns;
meioVert      <= to_unsigned(30,8) after 0 ns;
meioImagem    <= to_unsigned(31,8) after 0 ns;

in_janela <= '1' after 0 ns,
             '0' after 5 ns,
             '1' after (1 sec / frequencia_camera) * (numcols * numlin)- 1 ns,
             '0' after (1 sec / frequencia_camera) * (numcols * numlin + 1) - 1 ns,
             '1' after (1 sec / frequencia_camera) * 2 * (numcols * numlin) - 1 ns,
             '0' after (1 sec / frequencia_camera) * (2 *(numcols * numlin) + 1) - 1 ns,
             '1' after (1 sec / frequencia_camera) * 3 * (numcols * numlin) - 1 ns,
             '0' after (1 sec / frequencia_camera) * (3 *(numcols * numlin) + 1) - 1 ns;

IN_process: process (in_clock) begin
  if(rising_edge(in_clock)) then
    clk_count <= clk_count + 1;

    -- avanca as imagens
    case bloco_atual is
      when 0 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste0(linha, coluna));
      when 1 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste1(linha, coluna));
      when 2 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste2(linha, coluna));
      when 3 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste3(linha, coluna));
      when others => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste0(linha, coluna));
    end case;

    -- marcacao de linhas, colunas e parada na simulacao
    if (coluna = numcols - 1) then
      coluna <= 0;
      if (linha = numlin -1) then
        linha <= 0;
        --fim_imagem <= '1';
        bloco_atual <= bloco_atual + 1;
      else
        linha <= linha + 1;
      end if;    
    else
      coluna <= coluna + 1;
    end if;

    if (clk_count = 4 * (numlin * numcols)) then
      ENDSIM <= '1';
    end if;
  end if;
  

--when -label end_of_simulation {end_of_sim == '1'} {echo "End of simulation" ; stop ;}
end process;


END ProcessadorImagemGMAW_arch;
 