 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 1f 1a 13 11 0c 12 19 17 0d 13 14 12 16 0b 0f 1d 1c 1e 22 28 22 1e 1b 1a 23 16 23 27 2d 28 19 14 14 0f 0e 03 06 05 03 07 06 05 0d 09 14 24 20 24 1f 0f 11 06 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0d 06 0d 06 05 03 03 06 05 04 02 06 05 10 0f 1c 15 20 26 1d 16 24 1f 35 3b 2d 33 2a 2f 2b 2e 29 2c 2b 2f 31 2e 38 39 2f 37 2f 3b 3b 44 45 3d 36 34 29 2a 2d 30 1c 16 0f 05 07 1f 26 1c 1b 1f 29 30 29 2d 2f 25 19 1a 06 05 03 00 0b 1b 1c 1e 0b 06 06 05 06 05 03 00 0b 05 03 02 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 07 00 06 13 14 13 0d 05 0f 08 0a 0b 07 11 15 13 10 15 17 1a 16 20 28 2f 3b 46 45 4d 4f 4f 4d 53 57 57 55 4e 4d 60 5e 60 61 5e 5d 5b 52 5e 5f 50 4f 42 3b 44 39 34 3b 35 32 2f 1f 24 24 32 32 33 35 34 30 4a 4c 39 24 25 19 11 19 0e 0e 0a 11 25 21 25 12 09 07 09 06 13 12 16 10 05 03 00 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 04 06 06 05 10 0d 0b 13 0f 1a 19 17 15 19 21 19 1f 24 26 2a 2d 2e 2c 31 2a 32 3e 43 51 4d 5d 5d 5d 61 64 69 6a 6d 69 62 69 6e 68 6b 69 64 6d 65 6c 6b 6d 65 55 4b 4b 43 3e 3d 46 44 4e 54 53 5c 52 4b 4d 49 3d 38 3b 4c 50 37 34 2e 2e 32 29 22 23 2b 29 30 24 2b 27 1c 22 18 11 1d 18 1a 21 0e 0a 02 06 0c 07 0d 06 08 03 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 14 0b 06 07 0c 03 07 05 07 0f 1b 1e 25 31 2b 24 2a 2e 2d 2a 35 3a 30 31 41 38 30 34 38 37 3d 51 59 4e 58 67 6a 61 59 54 5d 67 60 6e 66 70 6a 69 66 6b 66 68 6d 5f 69 6e 61 65 5a 57 59 4d 5b 61 75 80 7b 6c 69 65 6f 69 64 60 56 52 54 4c 47 4c 4d 55 49 53 3f 3e 38 3c 3a 34 2b 2b 29 25 24 2a 1b 26 26 11 03 04 06 09 08 07 06 0b 10 14 11 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 06 01 07 10 0a 04 11 0b 0e 08 06 11 2a 27 39 36 42 4d 47 43 47 44 41 36 37 3c 36 45 44 4e 53 4f 46 41 4d 51 6c 60 66 6b 61 5b 5d 66 67 75 7a 75 7a 81 7c 6e 6c 65 65 68 6b 6f 6c 75 6d 74 71 6d 67 67 67 6c 70 8e 7f 76 6e 6d 70 74 7f 82 84 81 7c 6f 78 7f 7e 71 6d 68 55 60 4f 47 42 4d 37 3c 35 35 1b 2f 2e 2e 2d 19 14 10 0f 08 0b 05 0b 07 0c 17 12 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 0a 10 0b 0b 15 10 0b 15 18 24 25 29 35 36 43 43 4d 55 65 5d 5d 6e 6a 57 61 59 6e 71 74 7b 72 69 57 50 54 54 62 6c 6a 6a 57 5d 59 61 63 6d 71 7d 7b 7c 73 69 63 65 62 61 64 6b 67 65 65 68 64 66 65 68 5e 6c 6d 71 73 77 73 75 70 7b 81 80 94 95 95 8f 8b 8a 79 78 77 74 66 65 5c 57 5b 56 51 46 4f 4d 50 4a 38 2b 33 26 1e 1f 20 19 13 15 1a 15 14 1a 19 11 10 09 06 05 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 03 06 05 04 00 06 05 05 01 0c 06 0a 08 06 13 12 0b 0b 1e 2d 2b 2f 31 2a 2e 2f 2c 37 43 48 50 67 7b 84 73 74 93 96 95 8e 90 8a 94 9b 8b 86 6f 5b 58 58 56 5a 63 61 67 62 64 5b 65 62 69 6d 6e 6f 6d 6d 65 65 6d 62 65 64 5e 61 6a 6b 62 6f 5b 62 6c 64 70 6f 6b 74 75 74 75 74 76 76 7b 81 83 89 82 83 84 7c 75 71 72 6b 71 6f 6b 65 65 5f 57 58 5d 58 5e 5d 4d 45 40 36 32 35 30 2b 28 2e 21 1c 10 09 15 1d 0e 0f 09 0a 07 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 06 06 05 0a 06 06 07 0c 0f 16 19 13 25 2e 34 39 3f 3b 31 39 3a 36 44 4c 55 6c 80 99 9d 88 7c 6a 90 a4 ab 9c a1 a1 a0 99 86 7b 64 54 52 55 53 5b 58 5c 62 62 5f 5a 65 5d 61 61 64 5b 60 67 64 5c 63 5f 58 5e 65 64 62 6a 6b 64 69 60 61 68 6a 65 71 6a 76 6f 7a 79 6e 7b 7a 7b 7b 7b 7e 87 84 7f 7a 80 79 81 74 6d 76 6b 69 6a 67 68 6b 66 65 61 5d 54 4f 4a 44 4d 3e 3a 38 2b 30 2a 1a 28 1e 14 11 10 0e 14 0a 0a 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 0e 06 05 05 0d 07 05 11 09 15 16 24 2d 30 38 3f 4c 44 52 52 53 50 55 52 66 6f 76 86 91 9d aa ad 9b 74 67 6d 7e 9e af ad a6 a2 9d 8f 7b 62 5c 5d 52 5a 5c 5e 5f 4f 5e 60 60 66 62 62 62 5e 65 62 64 6a 60 62 5f 5c 65 5f 6c 67 65 70 67 6d 6c 6e 6c 6d 68 65 70 72 73 72 74 7e 74 7c 7a 7b 7f 7e 7f 8a 8b 80 82 7a 7e 7d 7a 7e 75 74 79 7a 70 69 78 6d 70 6c 6e 6d 59 5c 5c 55 5a 57 4b 39 44 2f 35 32 2f 29 1c 24 21 1b 20 1c 18 0e 04 09 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 01 06 07 05 05 0d 0d 0b 0b 10 0e 0f 1f 1f 38 40 4f 57 59 62 65 6a 6c 78 7f 83 81 8b 9c 95 aa b8 bc b7 b9 9b 7c 6f 64 6a 6e 75 8a 8d 90 84 79 77 63 5e 55 57 5c 5c 5b 57 5e 55 5e 67 63 61 68 5f 6c 67 66 62 6f 6b 61 61 65 62 64 6a 67 68 6f 76 78 76 72 76 6f 69 73 71 73 75 72 68 75 81 7b 7a 7e 77 81 85 8d 91 8d 8a 7f 81 7e 87 82 80 7c 74 79 7e 75 6f 73 71 78 70 6b 68 65 60 63 65 63 64 4a 57 4a 48 43 41 32 37 30 29 2e 2f 26 2e 2d 19 11 0a 05 06 04 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 0a 0c 0d 0d 19 1b 1a 24 31 40 4b 5a 61 6c 85 8f 93 8f 9e a4 a8 b0 ab b3 ba b9 c2 c4 c2 b8 a3 84 7b 70 6b 5f 6c 70 64 6a 71 6c 66 66 61 60 60 5d 5e 65 68 5f 5f 5c 5b 5f 5d 5f 59 5f 5d 61 61 6a 66 6a 5e 6b 68 6d 70 6b 70 6c 72 75 7a 73 77 78 74 6f 7b 76 76 7e 75 7d 75 7a 7d 7c 75 74 7c 82 80 8f 96 8a 85 81 81 84 84 82 83 7e 7e 79 6e 75 74 78 75 6e 6e 61 61 63 6a 67 62 64 64 63 5b 5e 55 53 54 4b 3e 3e 37 39 35 2e 2c 28 23 1a 0b 17 09 0b 06 0c 03 03 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 05 06 0b 06 10 14 1a 20 1a 22 25 34 45 57 6a 78 7e 8a 93 a7 aa ac b7 b8 c2 c8 c6 c8 ca bf b8 b5 a5 95 8a 7b 7c 6e 73 70 67 6f 6f 69 66 69 6e 6b 64 68 5d 64 5c 61 5f 60 5e 5c 67 60 5b 64 60 68 5f 69 68 68 67 6f 6d 6a 6b 67 6f 71 78 71 79 7e 81 7b 82 7b 81 7c 76 74 81 76 7d 79 81 71 7d 80 7f 81 7b 82 7d 83 84 94 88 81 82 85 8a 7b 87 83 7b 7c 7c 73 7a 6e 79 70 70 6d 73 74 6c 68 67 66 67 6f 67 65 65 58 58 56 55 54 4f 44 43 3e 45 34 26 25 22 18 14 0f 03 0d 0b 10 09 08 0a 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 08 0a 0a 06 0c 1a 12 22 2c 31 39 3e 46 45 53 5b 63 6e 72 75 7b 7e 8a 8f 9c ad ae b1 b6 b5 b9 ad 9e 9a 89 87 76 7a 75 6f 76 6c 71 6e 73 6f 70 6d 71 73 6d 71 71 6b 6b 5e 5c 5d 6a 64 69 62 64 66 67 66 69 62 70 63 6e 75 6a 6d 68 6d 73 7c 76 75 7b 86 76 84 7f 87 8e 80 7e 81 81 7d 7f 80 76 7e 77 7e 89 7c 81 80 82 81 81 89 92 84 85 8d 88 89 82 7c 85 7f 80 7b 6f 7b 71 72 75 74 6c 70 76 69 70 6d 6b 6d 72 68 60 62 62 61 63 60 59 59 64 55 4e 5f 4a 39 2e 1a 17 0c 11 15 0c 15 0e 06 09 12 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 06 08 0b 06 0e 0e 19 1e 26 2a 37 42 4a 54 53 61 62 57 5d 5c 61 6a 69 69 6c 6a 70 74 79 7a 7c 88 8a 89 84 79 75 77 6e 71 71 75 72 6d 72 6d 71 76 74 71 71 80 74 72 6f 6d 6e 75 70 6e 6d 6d 6f 6a 63 64 64 64 63 6d 74 6c 70 6a 72 71 74 78 83 7b 7f 7d 7d 81 81 89 83 8d 90 8c 94 84 87 83 7f 84 84 83 84 83 87 80 80 83 82 7b 7f 7b 8e 97 86 81 86 84 88 88 7e 82 88 7b 7d 79 76 75 71 76 7b 73 79 75 72 71 74 6f 74 6f 65 63 6e 5e 64 5f 5b 5c 5c 64 6a 74 7f 71 4b 33 2a 13 15 17 15 14 18 17 0f 0e 0c 05 0b 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 03 06 05 03 02 06 05 0a 08 09 11 12 1b 21 2e 3f 44 4f 51 59 5f 6c 61 64 63 63 65 66 69 67 66 6f 6a 70 72 73 68 6e 74 74 6c 76 6f 79 76 6b 76 78 78 7c 74 77 7e 82 7a 7c 70 6e 7c 74 74 7b 7e 7a 70 76 6f 7b 72 7b 73 65 68 70 6f 6c 6e 68 74 6d 73 76 7f 7c 7a 7b 82 87 8a 80 8c 8d 8b 8d 92 96 9b 95 9a 85 90 8e 8b 92 8b 83 84 84 87 84 7d 8d 86 83 84 86 8c 8f 89 84 87 7f 86 87 8b 82 83 81 7e 80 75 83 80 74 7d 79 7e 81 7b 7e 72 70 75 77 67 6c 67 71 65 67 5d 64 64 69 69 7c 95 85 64 61 50 42 36 22 12 1b 1b 13 18 15 10 03 02 06 06 05 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 03 0d 11 0d 1a 17 26 26 35 44 45 51 5f 5e 64 64 67 70 6d 6e 64 6a 6c 6d 77 64 6c 65 6c 66 7b 69 75 70 7b 73 6d 75 6c 75 71 7b 7b 75 75 78 74 82 75 83 78 7b 86 7f 83 88 83 85 7d 80 7b 79 79 7a 76 77 79 7d 74 73 73 73 6f 6c 72 78 71 7a 7d 80 89 85 8a 87 91 8d 91 99 96 98 9d a2 9a 9c 9a 94 9b 92 95 90 8e 88 96 8a 8d 89 89 85 83 86 7e 8f 94 8f 80 8a 83 87 8d 8f 86 8d 84 82 87 7e 82 84 82 81 84 77 7b 77 84 7f 7d 83 7a 7c 77 76 6a 6a 72 6d 65 62 6b 68 66 6e 74 72 88 86 71 5b 47 33 41 3a 2a 1a 19 0c 05 08 0d 06 0a 06 05 0a 0d 08 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0c 0e 07 18 18 23 35 32 3f 43 4f 59 58 5d 65 6f 6b 68 66 78 75 6d 79 75 70 6d 69 69 72 6f 6f 71 71 6a 6f 70 76 73 73 70 6e 76 72 75 78 72 7a 77 7a 75 84 77 84 83 79 88 7f 8e 8a 8b 8c 7e 7b 82 88 7b 84 82 83 78 7f 7d 78 7a 74 72 82 7d 75 7b 84 7f 8b 91 84 94 95 93 9c 9c a1 9e a5 a0 a0 a0 9c 9b 9c 9c 97 94 90 8f 95 94 90 88 8b 83 84 83 84 88 9d 8f 8b 87 8a 84 8d 8a 8b 8f 8d 87 89 89 8a 8b 81 87 88 8c 84 89 86 7a 85 7c 81 85 7f 76 78 6e 68 69 72 70 67 66 66 68 6e 6c 84 96 92 7d 69 63 5e 4f 43 26 1b 11 10 12 12 09 0b 03 0f 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05
 03 07 06 0c 18 22 2d 39 3e 43 49 5a 57 62 65 6b 6c 66 70 6d 75 76 76 6a 6d 72 76 78 70 6e 70 6c 70 74 7b 70 6b 6f 74 73 73 76 75 76 75 72 74 78 77 76 7c 83 81 88 86 86 8e 88 8e 8b 8b 8e 91 91 90 89 85 86 87 89 85 88 81 81 7e 78 84 78 7b 7c 7e 83 83 8e 93 95 8f 9a 99 a1 9d 9e 9a a4 a7 a1 a8 a4 a5 a3 a3 99 a3 9f 9a 97 9b 93 91 91 89 90 80 8d 81 8e 97 93 8f 85 8b 90 90 8e 8e 94 97 91 92 91 89 8d 8d 90 89 94 90 8c 98 84 91 8b 8f 8d 93 80 81 7b 7a 74 72 6a 6e 6a 6d 69 66 69 6b 75 89 91 8a 88 7d 6b 63 52 34 26 1a 10 0c 0f 0e 0d 10 10 0e 10 03 06 09 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0c 16 18 19 2b 2e 41 43 52 58 5f 62 61 63 68 6d 6e 73 76 77 79 7a 76 79 76 78 79 7c 70 70 71 75 6f 70 6f 75 75 74 79 76 6d 77 6f 7b 7f 78 7a 7b 77 79 7d 83 8b 80 88 8b 8d 94 8b 87 92 8e 93 9d 93 9a 8f 8e 98 97 8c 91 8c 88 8e 8c 90 8a 89 8b 88 8c 89 94 94 9e a1 a0 a7 a9 a6 af a8 ab a0 ac b5 ad af ad a8 a9 ab a6 a5 a2 a3 96 9c 91 8f 87 8c 90 89 89 8c 91 94 8b 8c 90 91 92 98 9b 97 99 a0 99 9b 94 93 99 9a 9a 96 9d 90 9b 95 93 96 95 95 8c 8f 88 87 78 71 78 75 6d 74 71 70 6a 71 64 6d 7d 85 8e 8a 88 82 73 65 59 3c 35 1f 13 18 17 0d 15 10 0f 14 0d 0d 07 05 03 02 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 01 0a 0e 29 2c 35 36 47 50 60 6c 73 6f 67 5c 62 64 71 6c 74 6b 71 78 73 77 77 78 77 77 76 7a 77 71 71 6e 6b 6d 74 75 7d 74 77 78 73 79 77 76 77 7b 80 7f 7f 82 84 7e 90 8b 89 92 8f 8f 95 94 93 98 93 98 9b 90 9f 99 9a 9a 99 9f 9b a0 9b 9d a0 a1 a1 a1 a7 a8 a7 a7 b3 a8 b5 b4 b2 b8 af b9 bc b5 b9 b4 b4 b4 ac ae a9 ac ab a2 9d a1 96 94 97 8d 91 8f 91 91 89 8c 91 96 8d 84 8e 89 93 98 96 9b 93 a1 96 9d 99 a3 a2 98 a1 a2 a4 a0 a5 9a 9e 9a 9e 99 96 8d 84 89 7d 7a 7b 75 6f 73 70 6f 69 65 66 62 65 65 6a 73 7c 7e 75 70 6e 6a 4f 32 29 1f 17 1d 0e 12 0b 11 11 07 08 0e 06 0d 06 05 03 01 08 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0d 0b 15 25 30
 32 35 3c 48 58 74 75 6f 64 66 65 64 67 67 67 71 74 70 7a 7e 7c 7e 7d 7c 7b 7c 71 77 71 6d 6d 79 78 7a 7a 82 78 7a 76 80 82 7f 7b 7e 75 80 7c 7c 82 7e 87 84 8c 8f 94 90 90 9c 9d 98 9f 9c a0 9c a2 a9 a5 9a a1 a0 ac b6 b0 b0 ba b5 bd ba ba be b5 bb bf bb b6 c3 bf c3 be bc b8 b8 bb b9 bb b8 b5 b5 b2 b0 aa af ab a6 9d a0 9c 9a 92 96 94 90 9a 94 8f 88 8f 8d 91 8e 91 94 96 a3 a2 a1 9e a3 a3 a0 a5 a2 a6 a4 a2 a4 9d a4 a1 a1 a6 9f 9e 9e 9a 9a 8c 8b 7f 7a 7a 79 6f 68 6b 6c 58 66 63 5d 60 63 63 65 5f 69 63 68 67 70 74 6a 49 30 25 1f 23 1f 18 17 15 14 0a 0a 0a 06 08 05 03 06 08 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 07 06 08 0e 1d 27 35 31 31 42 5a 73 73 6f 69 6b 66 6b 64 5e 63 65 6f 7d 77 75 79 79 78 83 82 80 87 87 83 7c 7c 7b 75 79 7a 78 80 80 77 7c 7c 87 88 82 8d 81 85 82 8c 7b 8a 89 8e 92 89 90 89 9d 94 98 aa a4 a6 99 a2 a1 a0 a6 ad aa b2 bf c0 c5 c7 cd d2 d4 db d9 d8 d6 d4 d4 d6 d0 cd d1 d0 d4 c9 d2 cd c8 c7 c4 bd b9 b7 b8 ba b7 b1 b7 ad ab aa a7 9b 9e 97 9e 98 99 89 93 94 90 91 91 99 93 91 9d 9a 9c a5 a7 af a8 a9 af a7 ab b1 a4 ab a8 af ae aa a2 9e a5 a1 a3 9f 9c 89 85 83 86 7d 7a 74 74 6c 65 61 66 5d 61 5f 5b 5d 50 5b 58 57 5e 67 6f 85 88 69 61 3b 29 22 29 1b 14 17 16 1b 0e 19 12 14 07 0d 0a 06 0d 0a 06 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0b 0f 25 2a 2b 37 2e 51 67 6f 80 6b 62 66 64 63 67 61 5e 67 66 76 78 76 7d 78 82 78 85 85 84 86 82 7c 80 78 79 7f 75 7e 7d 83 80 7f 7f 84 85 7d 86 89 87 8a 88 88 90 89 8e 93 94 8e 9b 96 9b a4 a0 a9 a5 a5 a4 a3 ab ad ad b2 b6 c4 d6 e1 ec e3 ea f1 e9 f3 ea ec e9 f0 e6 e8 e5 e0 e6 df e1 e2 d6 d4 d0 ce cc c4 c0 be c1 b9 b5 af ab b2 af ac a0 9c a0 99 9d 95 94 94 91 92 97 93 96 93 91 96 a2 a8 a6 a4 ab af af b0 b0 a5 a8 ab b7 b8 b3 b8 a5 b1 ad a8 9f aa 98 a1 95 92 8e 83 84 76 77 6e 71 6c 69 6e 5f 61 60 5f 5f 5d 5e 52 59 56 51 62 6f 96 93 7e 76 61 54 3e 36 1c 25 20 1f 20 1f 2b 1b 16 09 05 05 0f 0b 0c 07 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 03 02 06 0b 11 19 1c 27 2f 34 39 5d
 6f 77 76 6b 5f 61 64 5f 59 64 61 68 69 69 70 6f 70 76 77 84 85 87 81 84 84 84 81 7e 82 80 74 7d 7e 7b 7a 83 85 82 8a 88 90 92 8d 91 89 94 95 90 94 8f 95 96 92 9d a0 9f a4 a6 a6 a7 ae ae ac b0 a9 b3 b9 bd d8 e3 f3 fa ff ff ff ff ff ff ff ff ff fc f9 fc f4 fa f9 e8 ec ee df e2 d6 d6 d3 c1 c6 bb c0 b9 ac b1 ae b7 a5 ad a0 9f 96 98 99 8a 94 92 8b 8c 97 90 90 9d 9c a2 9e a1 ae ae b1 b4 ad b0 ac a7 b4 b6 b8 b0 ad b1 b4 ae ae af ac a2 a5 9e 85 8a 81 7c 80 75 72 6f 62 64 63 65 68 5f 56 5a 54 5b 57 54 4a 4b 59 64 85 8e 89 83 7b 83 64 4e 40 40 3e 3b 39 32 25 1f 19 0b 0a 04 0b 07 0b 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 0b 08 13 1b 20 32 46 49 6c 7b 6f 69 65 5f 67 66 60 69 63 6b 6a 65 6e 74 6b 71 79 79 80 86 7d 89 8f 91 8e 89 86 8b 8a 82 84 84 84 7f 81 89 89 86 80 8e 94 9b 9e 9c 9a 9e 9b 9d 98 9f a1 9f 9e a2 a1 9f a7 ab a9 af ae b1 b7 b3 b5 c4 c4 d5 e2 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 f6 ea e4 e4 e4 db ce ca bf b6 b0 b5 ba b1 a8 ad a1 9d 9c 9a a3 93 97 91 93 92 92 9e 98 98 9c a7 b0 b4 b9 b8 b1 b3 b7 b7 b0 bb bc b5 bd bc b3 b8 b2 b1 af b0 ab a9 87 9a 8d 8d 85 7f 7e 79 75 74 68 61 6c 70 64 62 64 54 5a 54 55 5b 5a 4f 55 5a 62 75 72 7e 8b 8f 87 80 78 6f 5c 54 51 3d 38 2f 1c 0e 14 11 15 13 10 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 06 07 0e 19 20 26 31 4f 5c 6f 88 7f 68 61 5e 60 60 64 66 67 69 67 6f 6a 72 6b 6e 73 78 7a 80 8c 85 8c 8e 8b 9d 8c 93 89 89 8e 86 88 88 90 89 96 95 90 97 9d 9c 96 9e a1 a7 aa a2 a7 ac a9 a3 ae 9e a9 ad a6 b4 ab b1 b1 ad b4 b9 b5 b0 c6 d1 e4 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd f8 f2 f0 f2 e4 de d6 cb c6 bb b8 bb b1 b7 ab a6 ac a0 a0 9b 9a 94 94 9b 97 9b 97 94 a0 a6 a9 b6 b4 b9 b6 bb bb ba b6 b4 b7 bc c0 bf bb ba ba bb b1 af ba a9 a6 ac 97 99 8e 85 7d 7e 78 7b 7b 72 72 71 66 65 69 5c 58 58 52 57 51 57 50 51 54 54 57 62 71 7f 8b 8f 8e 95 82 72 63 51 4f 46 35 22 1e 19 18 15 0b 17 06 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 02 06 0c 0f 0c 14 14 25 38 4e 72 84 85 83 6c
 64 5e 5b 64 62 62 66 68 6e 72 68 77 65 70 73 76 76 73 84 88 8b 87 95 97 95 8c 93 91 92 8e 90 8c 8e 8d 91 94 8e 96 92 a0 a3 a2 ac a7 a9 ad a6 ae ab ad b2 b6 aa ab b1 b5 b2 b3 b1 b3 b7 ab b3 b7 c0 cc e8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fa f3 ee dd d0 c3 bd ba c1 b9 ae b3 a7 ac 9c aa a6 99 98 9a 99 9a 93 9c a0 ab b1 b4 ba ba b7 bd be c7 c3 c3 c2 be bc bf c2 bc b8 b8 b9 ba af b1 b4 a5 ab 9f 99 96 8c 85 79 7d 73 74 6f 6f 6b 6b 66 6b 5d 5c 55 4d 4d 5b 53 52 50 56 56 56 4e 5b 64 7b 87 96 a1 96 84 75 63 5d 55 4e 48 2f 26 0e 0c 13 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 0b 0a 06 07 12 1a 1e 28 3e 60 7f 92 88 7a 79 69 5b 64 63 5c 60 66 62 69 67 6f 69 6e 6a 6d 74 76 7f 7e 80 92 8b 91 91 97 99 91 93 98 96 a0 97 8c 97 94 98 9e 94 9a a3 a3 ae ac b1 b5 b7 b0 b0 ba bb bc b7 c0 bb ba bc c2 c0 b7 bf bb b9 be be bd cf d9 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f1 e6 c5 c1 b8 bc c0 ba b4 ae af a9 a9 a6 a5 a3 a1 a0 a1 9a a0 a9 ad b2 bb bf c3 c2 c4 c0 c5 c4 c5 bf c0 bd be c4 bf c0 c1 c1 b9 b6 af b2 b0 a4 9c 9b 97 92 89 85 7b 7f 7d 77 75 76 71 6b 5d 65 60 5a 64 59 59 60 54 5b 5d 59 5c 60 56 62 64 6b 7e a6 a5 90 8f 7c 72 62 5f 4d 35 1c 12 0c 12 0d 0b 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 06 07 06 04 09 16 09 17 24 20 3c 63 85 97 93 7a 62 6a 72 6d 6a 64 65 64 69 5e 73 64 6f 70 71 72 71 79 75 7d 7d 88 86 92 9a 9e 93 a2 98 9a a4 9d 99 9b a3 9c 97 a0 9f a4 aa ab ad a6 b0 b2 b5 ba bb b4 c0 c0 c3 c3 c3 bd ba cb c2 c1 c6 c5 c3 c2 c4 c9 ca da ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f8 d7 bd c5 bd c5 ba c1 b9 b0 b2 b2 ad a8 a6 ac a2 a7 ac a8 a9 b8 c0 be c2 c5 c8 cf c1 cc c5 c7 cc c8 c7 c8 c6 c1 be bc bf b4 b6 b6 b2 ae aa a8 a0 a5 91 8d 84 86 7d 80 80 7b 73 6b 68 71 64 5d 5c 5b 5e 55 62 62 5e 5c 63 5d 5f 60 5a 5e 64 71 8c a4 a5 9e 8b 81 6e 60 43 33 25 17 11 15 0f 06 11 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 09 14 19 17 1a 25 2e 32 5d 7e 85 81 7a 6c 67 67 67
 72 6c 68 60 5e 63 6a 67 62 6e 70 6b 72 78 78 7e 79 88 82 89 99 8f 9c 98 9d 9d 9b 9b 9f 9b 9d a2 9f 9f 9e a6 a1 a6 ae b0 b3 be be b8 c2 c1 bf c3 c9 c4 cc cb c5 cd cf ca d0 cb cc c5 c7 ca c7 d2 e5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e1 c5 cb c0 ca c0 c1 b8 bc b2 b4 b3 a9 ad ac a8 ae a8 af ac b5 c1 c0 ca cc cc d3 d0 d1 ce c7 c8 c8 c2 ca ba c6 c6 c2 c4 b8 b3 b5 b5 b7 b2 a0 aa a0 98 93 96 87 8c 85 7e 7f 73 78 6c 70 66 65 5e 5e 5f 5e 5b 64 62 60 64 64 5b 5f 59 64 61 62 7b 95 a0 a0 93 82 6e 60 5d 40 2b 25 1a 1b 11 19 17 0f 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 06 06 05 04 06 06 0f 12 1b 17 14 1d 32 52 84 9a 8b 76 67 54 63 60 63 65 66 70 71 69 63 68 6b 68 6e 76 6d 7a 6e 77 77 8a 8a 90 8a 98 9b a3 a4 a7 a7 9e a9 a0 a3 a3 a7 ad a5 aa ad af b1 b8 b3 b9 ba c7 c0 bb be bf c9 cd c2 c7 c9 cb d0 d6 cf d6 db d6 d1 cc cf d0 df ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea d3 cf c6 c2 c0 c3 bf c2 b8 bb be b0 ad b3 b3 b7 bb b5 c1 c5 ca d4 ca d2 d6 d5 d6 d1 d9 cf c2 cd ce c8 c9 c5 c9 c8 c9 c4 b7 b8 be ad b8 af a9 a6 99 9b 9b 96 93 87 89 84 80 87 78 71 74 66 69 71 69 6b 65 65 6f 67 61 61 5d 64 5d 65 61 60 6c 7d 86 94 8b 88 78 6b 67 57 3f 2b 2d 25 29 1f 20 1a 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 05 0a 02 07 05 08 08 16 1b 1c 23 27 20 2e 3e 66 8b ab 9e 77 60 5f 5b 5e 5f 6a 6f 6e 71 6e 6e 74 69 6c 71 74 6f 75 80 7e 86 81 84 86 8d 9c 9f a6 a9 a5 a9 ab ac a4 a8 a5 b3 b5 aa b0 b4 b2 b9 b2 b7 c4 c3 c6 c1 c7 c8 c9 c2 d2 d3 d3 d1 d2 d4 d3 da d8 d5 dd d9 d9 d9 d8 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 d5 d7 cd cf cd c7 c4 cb c0 c9 be c0 bc c4 c0 c1 c3 c6 c9 d2 d6 d3 d7 df dd de d7 da cc d0 d0 ce cd cc cf c8 c7 cd cc c2 bb b3 b9 be bf b2 af ad a4 a1 9e a5 98 95 8e 8f 87 7e 80 7c 72 74 75 73 6a 6d 70 64 6d 6f 6b 66 64 63 66 69 62 6c 67 6e 73 78 7d 75 79 69 64 61 61 50 40 3b 33 21 27 1d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 04 06 0c 0e 18 13 1c 1d 27 34 3c 4a 60 81 92 a1 a6 7f 5f 58 55 60 65
 6a 69 6d 74 73 72 70 6b 6c 71 6d 78 77 70 84 7e 7c 84 8f 8d 99 9d a7 ae af a4 b3 a8 b1 ae ad aa b7 b8 b8 b3 b7 c5 b8 c5 bf c5 c8 c9 c5 c8 c6 ce d4 d0 d6 d2 cf d9 dd da d9 dd e6 db e0 df e4 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e2 d6 cb d4 d7 d1 c4 d0 c9 c5 ca c8 c7 cc c6 c8 c9 d1 d1 d4 dc d6 d6 e0 e2 dc da d4 d0 d2 d3 d3 cd c8 d3 ca c1 c9 ca c5 c2 c0 b5 bd ba b4 b1 b4 ae a6 ac a4 a0 a2 93 90 87 84 7b 84 7d 79 77 79 70 74 78 71 79 71 71 67 69 69 60 65 65 66 6d 6c 6c 72 68 6b 6c 61 6c 76 76 62 4b 40 3c 30 25 14 11 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 04 0b 06 09 10 0a 09 10 12 1e 16 23 24 3f 49 66 7d 7b 88 94 95 95 77 5f 5a 57 61 64 65 65 6a 67 70 76 7a 75 6e 72 6e 78 78 77 76 7b 86 89 87 95 97 a2 a8 a6 ae af af b4 b1 b4 b8 b6 ba b9 bd c2 c5 be be c0 cd c4 c7 d7 d5 ca ce d2 d2 c7 d5 d4 d3 e1 e2 df df e2 e3 db db e1 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 df da db d2 d7 d5 d4 d5 d2 ce c9 ce ca cd d8 de d6 d6 e1 dc e0 e5 e1 e0 da dd d8 d6 d0 cf d4 d9 d1 d2 d1 c8 c3 c6 c5 c6 bc b8 be c0 b2 b5 b6 b2 a7 ad a6 a6 a0 9a 92 8f 89 8a 89 84 82 85 82 7b 7a 77 7a 75 77 74 68 6b 63 5d 75 70 71 67 69 67 71 6c 6c 67 6d 68 74 84 70 5a 52 45 30 21 15 10 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 0a 0e 0c 09 14 11 15 10 0f 19 18 1c 24 35 45 66 74 86 8f 8f 9e a5 9a 94 77 5a 57 60 5b 63 6d 6c 69 6f 73 70 7c 7f 76 78 76 71 7a 76 7e 85 83 86 91 99 9b 9e ab a6 b1 b0 bb bc be b9 bb be c2 c0 c7 c7 c7 ca c5 c9 cc cc cc da d7 d0 d2 d7 d9 d6 dc d9 dc de e7 e6 e3 e9 ec f0 eb e6 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e3 e4 de d9 de e1 d7 d9 db d7 d9 de df d8 e2 da db e1 e6 ee e5 e6 e5 e0 e0 dd e0 de df d5 d2 dd d4 d0 d1 d3 d0 cf c0 c5 bf c2 c2 c2 bf bb b8 ad af b0 a9 a5 a8 a6 9d 97 92 90 90 92 8d 8c 88 7f 84 7c 80 79 78 79 76 6c 76 6d 78 6b 73 75 6d 65 68 68 65 69 69 7b 94 8c 72 61 4c 4b 37 29 22 18 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 05 06 0f 10 1a 16 0e 11 18 1b 1d 2c 45 63 79 90 8d 9a 9e a0 a7 a4 88 6a 50 53 58 5e 5d
 69 60 6a 6f 6c 6c 78 7e 7f 81 7d 78 73 84 7f 8c 88 86 92 96 9b a5 ad ac ba b4 b8 ba be b8 c4 c4 c4 c0 c8 c7 ca d0 c9 d2 d2 d0 d2 e1 d0 d6 d5 d5 e0 d7 da dd d9 e1 e4 e4 e3 e0 e8 e5 ee ee fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e7 dc e5 e5 dd d5 df d8 d9 e3 d7 dd e3 e7 e7 e5 e5 e8 eb ee e7 e5 e5 e2 e2 e2 de dc dc d5 da d2 d9 d5 d7 d5 d0 cc c8 c6 c5 c7 c1 bf bc be bd b3 b5 b2 ab ae a3 a5 a0 a4 98 98 96 9a 92 92 8c 88 8d 87 81 7c 78 78 7b 6c 77 70 76 6d 6f 70 72 63 6c 64 66 6a 74 8a 9c 8c 76 6b 60 44 2d 2d 23 29 17 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0a 08 09 16 13 1f 1f 18 1b 15 29 26 35 5a 7e 8f 98 a2 9b a0 a0 aa 9f 7d 5c 54 56 5f 61 61 62 67 6e 69 6d 6d 72 74 84 86 7e 80 78 74 81 82 88 8c 92 9b a1 a2 ac aa b6 b3 bd c1 c3 c9 c7 c4 c3 c6 c4 c7 cb d2 d0 d1 d6 d9 d1 d1 be be dd d8 d7 df d9 d9 e1 df e1 da e8 e6 e7 eb e8 f2 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ea e9 e5 e7 e1 e0 e0 dd de e1 da e5 e3 da e0 dc e9 e6 e4 f0 ef ea eb ec e5 df e2 dd dd e1 d2 da d1 d3 d2 d4 d2 cb d1 c5 c7 c1 c5 cc b8 bc bf b3 b7 bb b5 ae aa a6 a8 a5 a2 9e a3 98 9a 9d 94 89 8f 7f 82 83 7e 81 76 75 6f 6c 68 71 70 64 6e 69 6c 64 67 6c 74 8a 98 89 73 65 56 45 33 2f 2f 25 1e 07 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 13 14 12 1e 24 20 28 38 37 29 27 2a 34 48 69 89 9b a7 a9 a2 ab a7 ad 9d 6f 50 53 52 51 62 69 62 66 6b 68 6e 76 79 7c 7c 84 7f 84 87 8a 81 8c 86 89 93 97 a0 a4 ab b0 af b7 bc c5 c2 c2 ce cb d1 cb d1 d4 cf d5 dc d8 db de db e3 dd dd db e3 e3 e2 e0 e7 da dd df e8 df e5 e4 ec e6 eb f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f6 ff ef f8 f7 fd f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e4 ed e2 e6 ed e5 dd e5 e4 e1 e4 df e5 dd e4 e4 ec ed e9 f5 f2 e6 f3 ef ef eb e9 e0 df de d5 da e0 d5 d0 d8 cf d0 d3 ce c7 c6 c6 bf c7 bb b5 bf c1 be ab ad ae b1 a7 9c a1 9d a9 98 95 97 96 90 90 8d 8a 85 80 77 77 73 75 77 6f 70 6f 6b 6e 69 68 66 60 66 77 9c 91 8e 78 5d 4b 48 39 41 37 28 1f 07 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 09 0d 0d 15 17 20 26 35 3c 45 4d 39 30 32 3f 53 7b 80 9c b6 b7 a5 a4 95 86 82 59 55 63 59 5e 5d 5b
 69 68 69 64 70 72 78 80 80 82 85 8a 8f 8e 8d 91 8f 8d 9b a5 98 a7 a8 ad b8 b8 bc c6 c7 cd d0 ce d8 d8 da d8 d6 df dc dc df d8 e1 e5 dc de e2 d8 e6 e3 e2 e3 e9 e6 e3 de e1 ea eb f0 e9 ee ea ff ff ff ff ff ff ff ff ff ff ff ff f7 f6 ee ee ed f3 f4 ed ec f0 f3 fa f4 ff ff ff ff ff ff ff ff ff ff ff fd eb ea e8 e5 e0 e3 e0 e0 dc e2 dd e5 e7 e3 ec f2 eb ea f2 ee f5 f6 ee f2 f3 ee eb ea e1 e4 e2 e3 dd d7 de dc d3 d6 d3 d1 c9 cd ca ce cf bd ca c4 c1 c2 c1 b9 b2 ab a9 ad a8 aa a2 ac a3 9e 9d 99 90 90 92 8a 87 82 7d 79 81 75 73 70 6b 6d 6d 72 68 6e 61 5a 67 7e 99 9a 8d 7a 6d 63 5e 57 4c 43 2a 19 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 0e 0b 19 1c 26 36 42 54 55 5b 53 4d 4b 44 5f 7c 95 a2 a8 a7 a9 8f 7a 6d 5b 63 5d 59 5d 65 60 63 62 6d 6b 6f 74 69 73 79 7e 7e 89 86 92 90 89 92 98 93 91 a3 a9 9f ad b1 b3 bb c0 c0 cb d1 d0 d1 d8 d9 d6 dd d8 e1 de d7 e4 d5 e3 e3 e5 df dd e7 da e0 e5 e4 e2 e3 e7 e4 db e8 e5 ec ea ea eb f3 ff ff ff ff ff ff ff ff ef fa f2 f3 ee e4 e9 e5 ec ef ec ed ee f3 fa fc fc ff ff ff ff ff ff ff ff fa f1 f0 e7 e6 e7 e6 e6 e4 e5 e3 da e0 e1 de e4 e1 e8 ee eb f1 f5 ef ef f5 f7 ec f3 ea e9 e4 ed e6 e5 de e2 df d6 da d6 d6 d2 d1 d3 d0 c8 cd c8 c8 c7 c5 bc c1 bc b4 b4 ad ae ae aa aa a8 9d a3 9f 97 9b 92 8f 89 8a 8a 88 7b 77 7b 7d 7a 6e 6d 74 72 66 68 6c 5b 5f 63 75 89 98 89 7c 6f 67 6a 5f 4d 3f 31 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 0b 14 16 1c 1f 2e 43 45 4f 54 64 65 70 6b 70 66 80 7c 97 9b a6 a6 a5 86 6d 68 66 5f 60 67 5f 60 66 5c 66 72 6f 68 6a 77 76 80 8b 7c 87 87 90 96 96 90 96 9a 9f 9d a2 a6 ad b1 b3 b3 bb c5 bf ca d2 d5 d9 e1 de e1 dd e2 de df e0 e0 e3 e0 db e3 e6 e4 e8 e4 e4 e7 e4 eb e9 e6 e8 e4 ea ea e8 ea ed ee fe ff fa fe ff f9 f4 f9 f0 f1 f0 e7 ef f0 e5 e9 ef ee f0 f0 f3 f6 f6 fb ff fa fd ff ff ff fd f4 f8 f2 f5 ed e3 e6 e6 e4 e3 c8 df e2 e3 e6 e7 e0 ea e3 e3 e2 e9 eb f1 ee f2 f9 f2 f9 ed f2 ec e6 e2 e6 ea e3 e5 de e1 df d7 d4 d2 d6 d0 cf ca c8 d2 ce cb c4 be bd c1 c0 ba ad aa a7 af a9 ab ab a0 a0 a1 9f 96 96 8f 8c 84 85 7e 7c 76 79 6f 7c 74 7d 6e 75 5e 62 63 64 64 6a 80 94 8e 7f 6f 6f 6f 60 4f 37 20 1f 17 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0d 10 1c 18 26 2a 31 3e 48 4d 5d 5d 6b 73 76 7f 80 87 80 8d 90 9f a1 a0 93 7a 65 5e 61 63 63 6d 65 5e 68 6c
 68 6b 6b 6e 73 74 79 77 83 88 86 8f 8e 9f 8a 95 9f a0 a7 a6 aa ae aa b6 c2 b9 bd ca cc d2 cd df e0 de e3 e4 e4 e8 e9 de e9 e4 e6 ea ea ea e9 e1 e5 e1 eb e2 f1 eb f0 ed ee ea ed ef eb f1 f2 ec f2 ed f7 f5 fb f1 f0 ec ea ef f2 ef ef ef f0 f0 ee f7 f2 f5 f2 f8 fb ff ff fd ff fc fe ff f9 f7 f3 e9 ea e8 e1 e2 e6 e4 e0 eb df df d8 e0 dc de e2 e9 ec eb ea ea f7 f4 f8 f7 f5 f5 f6 ee ea f2 f0 e1 e5 de e3 e2 e0 dd dc d5 db cf d3 da cf d1 cf cb c8 c4 c6 c0 bc c3 b9 b0 b3 b5 b3 ad ad ab a6 a7 9c 9a 97 92 92 8d 85 83 82 76 7d 79 7e 7a 75 6c 6f 68 6c 60 65 58 67 61 70 7d 7d 75 74 6b 6f 60 4d 28 20 16 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0e 15 20 28 34 38 40 46 44 59 5e 6c 79 78 81 85 8f 8b 8b 8b 99 a3 9a 90 83 6a 61 5b 60 5d 61 6a 5f 64 67 69 6e 70 6f 72 7d 75 82 7c 81 89 8f 87 93 96 9e 9a a3 a4 9c a5 a8 b5 b7 b9 ba be c6 c7 c7 cd d0 dd df da e5 e3 ed e8 e4 eb ee e4 ec ec ec ee ec ea ec f1 ed e8 ef ee e9 e5 f4 ea ec f2 ec f2 ee ee f6 f0 f4 f3 f4 ef f5 f2 f0 f0 ee eb f0 ed f1 f8 f8 f9 f8 ff fc fe ff ff ff ff ff ff ff fd f6 f3 f3 ea e3 ec e3 e0 ea e0 e8 e1 dc e2 dc e1 e0 d9 e3 ee f0 ee ef f2 f7 f2 f7 f0 fa fb f7 f9 f3 f3 ee e7 eb e7 ec e2 e2 dd df dd dd cf cf ca d1 d4 d6 ca cd c4 c4 b7 c7 b6 ba b5 b0 b2 a8 a1 a6 a6 a8 a0 a8 97 96 92 8b 8f 8e 87 85 7c 7c 78 7f 76 77 6c 6c 70 66 62 5f 64 5e 58 5e 68 6a 61 6a 6c 6c 62 42 29 16 12 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 11 25 20 2e 3a 45 58 5b 5f 60 6e 76 78 7e 89 84 8f 98 89 8c 8e 8e 8a 86 73 65 64 65 66 63 64 6d 68 64 71 67 70 75 74 77 72 7c 84 88 88 96 91 93 98 99 9e a3 a5 a5 ac aa af b3 bd bb c4 c0 c4 c2 d1 cd d6 de ea e4 e8 f2 f1 e9 ec f5 f2 f9 f9 fa f5 f1 f5 f3 f0 f0 ed ec f5 f7 f6 f2 f4 f0 fb f7 fa f9 f2 ee fb f0 f3 f5 f8 f0 f6 f5 f3 f1 e8 ef f1 fb f7 ff fb fc f7 fe ff ff ff ff ff ff ff fe ff fb f7 fb f2 ea e6 e0 df e0 e0 e6 e6 e4 e0 ec e2 e0 da e4 e7 e9 ed f2 de f1 ee f5 fc f5 fc ff f9 fa f2 ef f5 f1 ee e6 e9 e4 e1 df e5 dd d3 e3 d7 d0 da d6 d6 c7 cf c4 c0 bc c2 b5 b8 b5 b7 b7 b0 aa a6 a8 a0 9e 9a 9c 95 98 8d 87 8b 88 7e 86 7d 7f 78 7a 77 70 72 75 67 64 64 63 5d 60 59 6c 69 62 62 6b 70 51 42 30 1e 14 0b 05 05 02 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 0b 0e 1e 21 31 37 42 53 61 62 6d 6f 76 76 7b 84 89 8e 8e 95 88 89 87 8c 7d 71 5d 5f 66 64 65 6a 68 70 6f 70 6e 71
 72 6e 71 7b 7d 84 8e 8c 8c 8f 8b 9c 9e 9e aa a2 a9 ab ae b3 ba be b9 c2 c7 c5 c8 c9 d4 cd d9 e2 dd eb ee fb f5 f3 fa f9 fe fa ff ff ff fc ff fd fa f6 f6 f9 ff fd ef f5 fb f4 f5 f7 fa f6 f7 fa fd fd fb fc f5 f2 f6 fb f4 fb f6 f8 fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f0 eb e6 e5 da e4 de e3 e6 e0 d9 e1 dd e3 e8 e4 e3 e8 e8 ed f3 ee f7 f5 f5 f5 ff f9 fd f2 f1 fb f0 ee ee eb ee ef ea e2 dd e0 e3 db e0 d9 db d9 df d0 ce d1 c6 c6 c6 c4 c4 ad b6 b9 ae b0 af a5 a5 a1 98 96 98 94 8c 94 8a 89 80 78 7a 85 76 78 79 75 76 73 60 70 68 68 69 65 66 60 63 61 64 68 64 57 43 27 24 13 07 08 04 00 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 09 1a 1c 22 34 3f 4b 5d 6e 72 71 7c 7f 7b 84 8a 90 88 86 8a 85 79 74 6c 6a 60 5b 5f 6a 62 61 67 6b 71 6b 76 6d 6a 75 76 78 7f 7d 82 89 8e 8a 92 92 9a 97 9b 9f a7 b3 aa b0 b5 b9 c1 bb c0 c8 cd d2 cf cf d6 d6 e1 e1 ed ed f1 f7 f6 f6 ff ff fe ff ff ff ff ff ff ff fd fb fd f6 f8 ff ff fe ff ff ff ff ff ff ff ff f3 f9 f6 fb f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec ec eb e3 e1 e2 e2 e5 df df df e0 dc df e1 e3 e7 ee f1 f3 f6 f1 f5 f6 f9 ef fe fc f4 fa f5 f4 ef f1 f6 ee f3 ec ed eb e1 e8 e2 d9 dc de d9 d3 d7 d1 d1 d1 c7 c8 ca c2 c3 af b0 a6 a5 ac a9 a6 a0 9b 9b 8f 88 93 8b 8d 83 82 84 82 79 78 82 7a 6f 70 69 6a 6f 67 68 6b 6e 6c 71 65 62 65 69 5f 5b 4f 35 24 18 11 0f 07 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0b 14 1f 23 30 2e 4a 59 66 77 77 72 7f 82 7d 8b 8b 91 89 80 7b 78 6a 66 6a 68 5e 66 6c 6a 6b 59 6d 6c 72 70 6f 76 77 79 75 77 7e 81 7b 8e 8a 8b 93 95 95 9e a2 a4 a9 b0 ac b5 b4 bb c2 c4 c6 d3 ce db d8 df d6 e1 e3 e1 e8 ed fb f3 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 fe f1 ef ea e1 e0 eb db e2 df dc e1 e4 e3 e3 eb ed e9 f4 f6 f4 f6 f6 f5 f3 f5 f9 fa f9 fc f7 f4 f1 ed ee e8 ea ec ec ea e3 e4 e5 e8 e0 dd dc dd de d4 d0 d6 bd c7 c2 c1 bd ba ab ac ae ae a3 a7 a0 93 94 91 87 8e 8e 8a 84 82 84 84 79 7d 74 71 79 6f 75 70 79 76 71 79 75 79 79 71 66 69 60 67 63 55 3b 2f 1b 1a 0b 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 14 1b 29 28 38 33 56 68 72 82 79 7e 7b 77 82 82 82 84 84 76 76 65 6f 61 64 68 61 67 6f 6b 70 6a 73 67 7f 7f 76 7f 7e
 71 79 83 7f 84 81 87 7e 86 9c 98 97 a2 9d a3 a6 b0 b8 b2 bf b4 bc d2 d2 ce d3 dc e3 e7 e5 eb e7 f3 ef f1 f4 fa fe ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fb f0 e0 e1 e6 e2 de e5 e0 e4 df e1 e1 e8 e7 f2 eb f4 fa f2 f3 f1 f9 f5 f7 f7 ee f5 f5 fc ee f5 f6 ed f4 f0 f2 ef ee e4 e3 e2 e9 e4 de d9 de d6 ca cd cc c7 c2 bf b8 b4 b1 a9 ac a7 a5 a3 94 94 98 90 8b 8f 8d 80 8c 81 82 79 79 7b 79 78 77 76 74 7c 7e 7d 82 83 80 86 84 80 71 6d 68 67 62 56 3a 33 30 1a 14 05 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 11 24 23 33 3e 4a 5a 64 77 7f 82 7d 7d 76 72 77 77 7b 78 6c 68 68 60 66 64 66 6f 66 6d 66 71 6c 73 70 73 6f 77 7d 76 7d 7d 7a 7f 7e 82 82 85 8c 87 8a 96 99 9d a0 a3 a7 a9 b4 b2 bb c9 c1 ca d5 d4 de e6 f1 ef f9 f9 f9 fd fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef e6 ea e5 e3 e9 e4 e3 dc e1 e5 e8 ea ef ef f0 f1 f8 f0 fe f9 f4 f1 f5 f7 ed f5 f2 f6 f4 f9 f5 f1 f6 f0 ef ef f3 eb eb eb eb e1 df d5 e3 d7 cf cd c7 c5 c5 ba b8 ad ac a5 a1 9f a5 9b 97 93 92 94 89 87 89 8a 86 80 86 7b 77 71 76 7a 79 7b 83 82 90 8f 98 98 9c 98 93 85 7c 74 69 65 64 5a 4a 42 33 18 0b 0c 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 1b 22 30 38 42 55 5c 67 7c 7b 84 73 78 71 6d 70 76 7e 69 60 67 60 61 61 65 66 65 6a 65 72 78 78 76 74 7f 78 7c 84 80 86 80 86 7d 7c 86 83 81 7c 98 8a 92 97 91 93 a0 a7 a4 b3 b1 b7 bf ca c5 cd cf d1 df ef f4 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fd ef eb e9 e6 eb e4 e0 e6 e1 e8 ea e5 e3 f0 f0 f2 f1 f1 ef f6 f3 f1 f2 f0 f2 f8 f0 f3 f4 f2 f5 eb ef f8 f3 f1 ec ea ec e4 e5 ea e2 e5 e3 db d5 cb c5 c6 c4 b7 af ac a3 aa 97 97 99 96 98 8f 99 93 80 89 80 8e 8a 7c 7c 81 75 71 76 79 7f 89 90 9b a6 a6 a3 b0 b1 b2 af a0 85 76 70 66 70 60 57 4b 33 29 17 0f 05 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 17 22 25 3c 45 4f 60 62 74 85 8b 83 70 6f 6a 74 74 77 6d 66 56 64 64 64 5c 69 6a 67 69 69 75 7b 75 7e 83 80 7f 80 7b 80
 8c 84 86 8b 82 87 86 81 8a 88 8d 91 92 9f a0 9f ac a1 a6 b8 ba bf c6 cb cc d9 df ed f4 f2 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 f8 ed f3 e6 e6 e5 e5 e9 eb ed ea ec ef f1 eb eb ee f3 e9 e9 f0 fa f7 ef f6 e8 ed f8 f8 f4 f4 fb f5 f2 f5 f1 f4 ed ed e7 e6 eb df df db cf ca cd bf bb b7 b9 af a0 a4 9a 9c 9d a1 9a 93 8e 94 8e 8f 8c 84 84 7b 84 84 81 89 76 7f 84 99 a5 c1 c9 c6 cd d4 d7 cb c6 a7 95 86 6e 6e 74 79 65 54 44 2b 17 13 10 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0f 1b 20 2c 31 44 54 67 73 86 8f 8a 86 6e 75 6d 75 76 6a 61 5e 5d 65 65 61 63 63 65 60 68 6c 70 7a 7b 79 78 83 86 88 86 8f 8d 89 87 8b 92 86 86 8e 91 95 90 94 92 96 98 a1 a7 a7 aa ba b7 c5 c1 c8 d1 de eb f0 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f5 f3 f8 ef e4 ec e4 e4 ea ea e8 f2 e7 ef e6 e9 f4 e8 f8 e9 f3 f4 ef ee ee f6 f7 fb fc f3 f3 f2 f6 f9 f5 f2 f5 f5 e7 ec e7 dc df d5 ce c8 c7 ba bb b6 b1 ac a7 99 9e 9c 99 98 91 93 93 8e 8b 87 87 83 83 80 80 81 79 7c 6f 86 87 a5 c0 e0 eb e8 e9 f0 e2 d6 cf b4 97 7d 75 77 7e 81 6c 5e 42 32 1f 1b 13 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 00 06 10 15 25 33 44 4b 5e 66 77 7f 8d 90 7e 75 7c 77 6e 61 5e 59 57 58 62 5e 60 65 62 67 64 65 68 72 74 7a 79 7a 7e 7d 87 8b 8a 92 8d 89 8c 8b 8a 8e 92 91 8f 8b 95 97 9e a1 a5 a6 ae b2 b2 b6 c3 c9 cf de e6 f3 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f8 f5 f5 f5 ed ef f1 e6 eb e1 ea e7 ec e7 ec e7 e6 f1 e9 ed f2 ec f1 f1 f3 f3 f2 ee f2 f3 fc f7 f6 f0 f2 eb ef f5 e2 e6 df d9 d1 d2 c8 c0 bb b6 b4 a3 a6 a6 9b 99 9d 99 9b 98 90 90 8a 8e 89 89 84 7c 86 7f 77 77 74 79 87 93 b7 d2 e6 ff fb ff ff f9 df cb ab 8f 7e 75 72 80 7b 6d 5d 3c 2e 2b 19 14 0b 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 15 1e 24 33 3e 52 5e 71 82 8f 9b 9a 86 84 78 74 67 64 5b 58 52 5e 5d 62 5e 65 66 64 5f 67 69 72 70 6d 76 7e 7c 83 85 8e 85
 8d 91 90 93 95 9a 91 96 9a 9c 98 9e a2 a6 a7 a5 a8 a4 af b7 b6 bf c2 d0 d9 e6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 fa f3 f7 f1 f0 ed e7 e9 e8 e4 e6 e5 e9 e6 e4 ed ec ed f6 f5 f8 f5 f8 f2 f9 f4 f4 fa f6 f9 f1 f0 f1 ed e4 ef e8 e6 de db d3 d1 c7 c1 bb b3 b2 b0 a6 a5 a0 99 98 95 97 94 8d 8f 94 85 89 85 86 77 80 81 76 77 78 7e 83 93 b4 c7 ec fd ff ff ff f8 e1 d1 a7 8d 76 6f 6e 84 87 80 67 55 3f 2b 21 14 0a 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0d 19 28 2f 3c 41 50 5a 76 81 8f 95 a1 89 84 7a 65 5d 5c 5d 57 56 5a 5d 5d 64 59 5e 60 6b 63 6a 6a 74 74 75 7b 7e 84 85 8a 8c 8e 96 92 98 9b 9a 9b 9b 9b a0 9b 97 a3 a9 a9 a6 a4 ae b4 b8 c3 c4 ca d3 e9 e8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fb ed fa f7 ed f1 e2 e3 e5 e1 de de e0 e5 ea ea e8 ea ee eb f0 f8 ec f4 f5 f0 f5 f5 eb eb ee ef e9 f1 e6 e5 da df e3 dc d1 c7 c7 c5 ba ba ae b3 b0 a5 a6 a0 9a 98 99 95 94 93 8a 83 89 7f 82 85 7e 7d 73 76 7a 86 8b 97 aa c5 eb f7 fc ff ff fb e9 d0 a4 8a 74 6e 71 84 8e 7a 64 51 3d 2e 2c 1f 12 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 0e 22 28 38 4e 4a 66 76 8d 96 9e 91 7b 76 67 5d 54 5a 57 5a 5e 55 59 5f 5e 5e 6b 67 5c 6d 6a 6a 6f 6c 7b 77 80 85 7b 87 87 94 8c 9b 98 a0 9a 9a 99 a3 a2 a2 a6 a5 a9 ae b2 b3 b2 bb b9 c3 cb d1 d1 da e8 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc f8 f5 f5 ed f0 e9 e0 db dc d8 df de e0 e1 e5 eb ec e9 ee f0 ee e5 ea ef ed e7 e8 e9 ec e9 ea e7 e9 e8 e5 df de dc db d6 d0 c6 c1 b4 be b5 ae ac a2 a7 a0 97 9b 92 97 92 90 8d 90 88 81 88 8a 7c 83 7f 75 72 75 83 7f 83 a0 b6 ce d8 ea f5 fd ff ef cd a3 7d 6f 6d 70 84 8d 76 6d 4c 47 38 2e 21 11 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 11 1b 23 31 42 4f 5b 69 80 89 97 99 8d 72 6b 5f 52 5a 5c 61 5d 59 5f 5b 60 60 64 5f 69 5e 5e 65 6d 73 73 77 75 7c 77 81 85 84
 92 98 90 9b a1 9f 9b a2 a5 ac a9 ab b4 af b8 b4 ba b1 c2 ca cb cc d6 d8 da e3 f3 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef f5 e5 ed e7 e1 e4 df db dd dc dd d9 e2 e6 e8 e8 e1 df e9 e8 e7 e0 e7 e9 e4 e7 e2 e8 e9 de e0 dd e5 e1 e2 df db d9 dc de cd c9 c1 b6 bc bc b2 b1 9f a3 9b 9c 99 9a 9e 9a 93 8d 90 81 7c 85 86 87 88 7e 75 70 7a 7b 78 8a 93 a4 b8 c3 d8 ed f5 fe ef c6 a0 88 6a 66 72 85 90 85 6f 60 4c 3d 2c 21 10 0b 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 09 17 28 2b 45 51 62 6d 83 91 9d 92 87 75 67 58 56 5d 5f 61 58 59 59 60 62 61 60 62 5f 63 63 64 72 70 73 75 7a 7b 80 86 85 8a 8c 93 8c 8f 97 9f 9f a4 a4 ac b3 ae b4 bc b0 c1 bf b9 c6 ca ca d6 d5 db da df f2 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f7 f4 ed e4 e6 da da dd d9 db e4 db e6 e3 e0 e4 e3 dd e1 e4 df d7 de da df dc df db e1 e2 de db de df e4 d7 d7 d7 e0 d3 d2 be c2 c1 ba b4 ae ad aa a4 99 9f a0 99 9d 9b 91 95 85 88 81 8a 85 81 81 7f 81 84 78 7a 83 77 7c 8d 8d a4 ab c7 ec ef f3 da bf a4 7e 73 67 6f 87 8d 83 79 61 51 37 32 24 10 0a 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 09 10 24 31 3e 56 68 77 81 93 9c 8d 7e 68 5a 57 57 5e 59 59 55 56 5b 60 62 5d 60 60 60 67 69 6f 6d 72 73 75 75 82 86 7e 7a 89 8c 8d 8e 90 92 9e 97 a5 a9 a2 af ae ae b6 b5 b6 c1 bd cb c8 ce d0 d6 d4 de e6 ec f4 f4 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 e9 e3 df e2 d2 da d3 db d5 dc d4 e0 da d7 d3 d1 db d6 d5 d5 d5 d6 d7 ce d2 d0 d2 ce d8 dc d9 d4 d4 cf d4 d6 ce d2 cb cb d0 c1 c1 b8 b6 b1 ac af a1 a0 9b 9c 95 9b 8d 96 8a 8f 85 81 82 83 84 80 7f 83 81 80 7e 79 78 79 7b 87 82 92 9c b4 c2 d9 d8 ce ad 98 7c 68 62 6c 89 8d 7f 76 5c 47 3a 33 21 18 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0f 18 22 31 49 55 6b 83 92 96 9c 88 71 62 54 5f 56 5e 68 5a 61 61 55 5e 54 60 66 5c 6d 66 5d 69 70 75 76 76 7f 7f 7f 82 85 88
 8b 8d 8d 8e a2 97 9c a4 a1 ad b1 af b9 bd bb c6 c3 c6 cc c9 d3 db d9 d4 e4 e2 e9 f3 f3 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 e7 dc e3 d5 d3 d0 d4 d7 d1 d3 d7 d9 d0 cb ca d1 d1 d0 d4 d4 c9 ce d4 d1 d1 d6 d3 cd d0 d0 d1 cf d4 ca d0 c8 cd cf cb cf d0 b9 c3 b8 ad ae b6 af a6 a6 a3 a1 98 95 99 9c 89 8f 8d 89 84 87 88 7c 81 82 83 80 7d 84 79 80 75 79 75 82 8e 98 a7 af b4 a8 99 88 6d 63 6e 6d 8d 90 87 76 5c 58 44 30 26 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 05 09 08 1c 29 28 40 54 6c 83 8f a2 99 78 6b 65 62 5f 62 60 5f 5e 57 60 5d 6b 5f 6b 62 67 6c 63 67 6c 73 72 72 75 7b 81 7d 85 7a 8d 8e 8c 8b 8e 99 94 9d 97 a6 a7 b0 ac bc bd c1 c5 c8 c7 ce cf d7 de e1 dd e5 ec ed f9 fc fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 dc d8 cc d0 cf d5 cc d1 d1 cb cf c6 c7 cc cd cb c8 d0 ce d4 cc c4 cb cd ce ce d0 c8 c6 c4 c9 c7 c1 c6 c6 c7 ca cf c3 c2 cb b9 ba ba ae a9 ad a9 a9 a9 96 97 9a 91 94 8e 94 8c 87 8b 89 81 83 8b 84 78 84 81 80 81 7a 73 74 7a 7b 80 7d 8a 8e 93 95 8f 7c 75 6b 63 62 73 8c 9d 85 79 62 45 3d 35 1d 11 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 10 11 20 2f 43 60 6b 88 98 95 89 72 61 60 62 67 62 5c 61 65 60 64 62 6a 62 60 69 5f 65 64 67 74 6c 78 75 72 7a 77 87 80 82 89 89 87 90 98 97 94 9c a2 a4 9f ad b5 b6 be bd cf cb c5 c8 cc d8 de da db e1 ed f7 ec f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef da ce c0 c1 d0 ca c7 cf cf c8 c9 ca c8 cd c4 c2 c4 c9 cb c5 c8 be c1 ca c9 c6 c3 c0 c5 c1 c2 c2 c2 c2 c0 c6 c3 bb c6 c3 b8 b6 b3 b9 a5 af a7 a4 9e 9e a0 9a 97 99 92 92 91 8b 93 89 80 7f 82 81 8f 80 81 83 78 7e 7d 7a 75 77 72 6f 76 7b 80 7d 81 6f 6c 6b 66 67 62 7a 90 97 88 7b 5e 4f 3b 26 1b 10 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 07 0d 29 33 43 58 71 8d 98 93 84 6d 65 63 5d 68 67 62 6b 5e 68 65 60 68 6b 62 62 65 6f 70 6a 6d 69 76 75 73 73 6f 7f 7d 88 8d
 93 90 90 93 9d 9d a1 9d a8 a9 a9 bf bc b6 c5 cb c6 cb d0 d3 db db da e3 f0 ec f5 f7 f8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb cb ce bd c3 c8 c6 c7 c3 c5 c7 c0 c6 b9 c6 cd c6 c3 c5 ca c4 c3 c1 bc c6 bf be bb c3 c3 be c7 ba c1 bf bb b8 c1 b5 c5 b8 bb b1 b3 b1 a7 aa a7 9f 96 9c 92 9d 93 95 90 97 99 93 8e 91 89 8a 83 80 87 7b 85 77 72 7c 7a 78 6b 78 6d 76 71 70 6f 76 6b 64 67 63 58 5f 67 6e 92 8e 8b 73 68 58 3f 3b 1f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0a 18 2a 33 48 65 74 91 9a 88 70 62 63 67 63 6f 69 63 66 61 63 69 61 66 68 67 65 6b 6c 6f 73 72 71 79 78 73 80 81 81 81 89 7f 89 92 8c 89 9d 97 9d a9 b0 a1 b6 b8 bc b8 be bf c5 cd ca dd de df e6 e9 e8 f1 f5 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa c6 c7 b6 c0 c3 bc b8 bd c2 cb c8 c6 bc bd bb ba bd be ba bd c4 b9 b7 be c2 c6 bb c0 bc be bd b8 bf be bd ba b6 b6 b6 b4 b2 a7 b1 a7 a1 ab a0 a4 a2 94 99 90 94 90 96 99 8a 93 8b 8d 88 81 89 8e 8b 88 80 7f 71 77 73 78 7d 67 6e 6f 67 69 67 69 66 65 63 6d 56 5e 65 6b 87 9c 87 83 5e 4e 46 2f 20 18 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 09 13 22 2d 3d 5e 75 88 97 84 6e 63 62 5b 66 62 68 62 6a 68 67 67 68 5c 62 63 6d 71 6d 65 6e 76 74 76 75 75 77 80 7c 88 89 87 8e 8a 8f 90 9d 9e a0 a8 aa a4 aa b5 b9 c1 be c2 be cf cd d3 dd e0 de e5 e9 e9 f4 fb ff fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa fa f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c2 c0 b7 bc bd c6 b7 b0 bb b4 be bf b6 c1 b7 b4 bb b3 b4 bd b9 b3 b6 c1 b4 b8 c1 b9 ba b9 be af b8 b9 b3 b3 ae b4 aa b5 b2 a9 b2 aa a0 a5 9e a4 9b 96 97 94 95 97 95 8e 91 96 92 89 87 86 87 83 84 85 7e 7f 75 75 6f 70 69 6f 6b 64 5f 5d 5a 63 5b 64 59 5a 58 5b 67 75 8b 95 8a 80 5e 4e 48 26 21 0c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 13 21 2a 42 55 76 8c 8a 72 65 6a 6b 62 65 6d 6a 69 61 69 69 67 67 6c 61 64 6d 6f 72 6e 66 70 72 7b 7a 7f 80 82 82 85 8e 88
 91 8c 91 9b 97 9c 9b a5 9e aa b0 b5 bd be c7 c0 cf cf c8 d9 d8 d9 e8 e4 ef f0 f3 f3 fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f5 fc f8 e8 f5 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c3 b5 b6 b6 b9 b6 bc b7 bc b4 b2 bb b5 bb b4 b8 b5 bc af c2 b8 b0 b2 af b7 b5 ae b1 af b0 be ae ac af ae b0 b5 b6 ac b5 a9 ab ab a8 a3 a0 a4 a1 98 95 9d 98 94 98 95 8c 8f 97 8b 8f 8c 89 87 8b 86 81 7d 79 6c 70 6c 67 6d 66 5e 67 64 5f 5e 63 59 60 5e 62 60 60 60 6e 89 8a 87 7b 68 53 3a 34 1a 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 0e 23 37 43 5e 76 8d 87 74 69 63 63 64 62 63 64 6d 75 6d 6b 6f 68 6c 69 69 67 75 73 6b 69 76 76 7a 79 7c 7a 7a 7f 89 91 93 8f 8f 94 9f a2 9d 9e a7 aa a9 a9 af b7 be c9 c2 cb d0 d5 d4 d6 d9 e2 e2 e8 f2 ef f1 f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fe fc f6 f9 ee f1 eb e6 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f2 fd ff ff ff ff ff ff ff ff ff ff c3 bb af bb b8 b6 b9 ae b5 b7 ae b5 bb b1 b8 b0 b3 b5 a7 b4 b2 ac ad ae ae b1 b7 ab b4 ab b2 ad ac ab aa b1 af a5 b3 ac af aa a1 a6 a1 a4 9f a6 95 9c a0 94 8e 94 8e 94 8d 89 87 88 91 87 89 82 7d 79 76 70 70 6d 68 6b 6c 6e 62 68 61 65 5f 63 5d 5f 5f 5b 57 62 66 6e 80 94 87 82 64 5b 39 34 27 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0f 1f 2f 45 60 7e 90 8a 70 6f 66 63 65 62 66 65 6e 6f 73 6f 67 6a 6d 70 6a 69 74 6f 75 73 6e 74 7d 74 7e 85 84 87 85 86 86 9b 8c 98 97 a3 95 a2 a4 a9 b3 b6 b5 b9 b8 bb c9 ca ce d2 d0 d8 d8 df e2 ee ef e9 f6 f5 f6 fd ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff fc ff f6 f8 f6 f3 ea ef ea ea e4 eb f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 e5 e9 ed f6 fe ff ff ff ff ff ff ff ff c9 bf af ae b3 b3 af af b5 b8 a9 ad b5 af aa a9 a9 af ac ae aa ae a5 b0 a8 b0 a7 af ae ad aa ab a5 a1 a4 a7 a5 ab a9 a6 ab a7 a5 a5 9a a2 9c 9d 96 95 96 99 92 97 8b 97 8c 8b 93 91 88 87 85 7f 78 7a 77 78 74 6f 6b 68 68 69 6a 67 61 65 5e 60 61 5a 60 60 5d 5e 52 62 81 90 8b 7e 5e 51 35 35 18 0d 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0b 06 16 2a 34 45 5f 72 86 85 74 67 69 68 64 69 6d 6f 72 6d 70 75 76 77 70 74 71 6d 6e 6e 70 7a 75 82 81 81 7f 8c 86 84 8e 8f 89
 8e 91 95 98 93 a5 98 a4 a7 ae ab b5 b2 ba be c2 c2 c6 cd d4 dc dd db df e5 ea e7 f1 f1 ef f1 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ff fb ff f5 ee ee e1 e9 ec df e2 da e0 e8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fb f7 ff f6 e6 d4 d8 d9 df e5 f1 fd ff ff ff ff ff ff c4 ad a6 ae ac ad ac ae ab a7 af aa a9 ab ad a4 ab a9 9c a6 ab a3 a6 a8 a4 ad a4 a6 a2 a1 a3 aa a4 a5 a0 a3 a9 a4 a5 9f a6 a5 a0 a5 9f 98 99 98 9a 94 95 93 92 8c 90 8f 8f 90 95 8f 86 7f 87 78 7b 6e 6b 6b 66 6e 66 67 65 6d 69 65 5a 5e 5d 60 64 60 63 61 5d 60 63 63 80 8f 89 75 66 51 42 30 1a 05 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 10 25 30 4c 57 79 7f 7b 76 6d 6b 68 60 63 6a 70 72 72 6f 71 74 7c 76 72 72 72 75 75 78 72 79 7a 84 84 84 88 89 8b 8d 92 8e 8e 90 99 92 a0 97 9d a3 a9 a4 ac af b5 b3 b2 c2 c3 ca ca d1 ce d9 de e7 df e4 e7 f2 f3 f6 f3 fb fb f8 ff ff ff ff f7 ff ff ff ff ff fe fd f2 f9 f7 f8 f5 f5 ef ea e7 e9 de e0 e0 e0 df e7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 de e4 e5 e4 db d6 ce c8 c9 d0 d4 d3 df f5 ff ff ff ff ff c8 a8 a9 a2 a5 b1 a8 ac ac b1 a7 ad a7 a3 a5 a0 a6 a5 a2 a7 a3 9f a5 a3 a0 a9 9f a5 a3 a9 a3 a5 a4 a2 99 a5 99 a0 a3 98 a9 9f 99 a0 9f 99 96 9b 93 99 99 8c 96 8b 89 90 90 8f 8f 81 86 7f 84 75 7a 73 76 71 70 6e 71 65 64 6b 5d 68 62 65 5e 53 63 61 67 63 5f 5f 5e 64 7e 86 82 7e 66 50 47 34 19 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 06 00 09 19 26 2d 42 5a 69 77 78 74 69 73 71 6b 6c 68 6d 68 6d 76 6f 71 77 7c 79 75 71 6e 6e 79 76 77 84 80 82 7e 85 89 83 88 92 94 95 90 94 9a a0 99 a1 9d a1 af a3 aa b3 b5 bb bf c6 ce cd d1 ce d7 d7 e1 e5 e9 e9 f0 f6 f1 f6 fb ff f9 f7 fd fe ff f8 f8 fa fb fa fc f1 ef f2 ef f5 f0 ed f1 eb ed ea e5 db d8 da d2 dc e6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dc c4 be c5 ca c7 b4 b6 b4 bb bc c2 c1 cb d9 ea f1 ff ff ff cb ad 97 a2 a0 a6 a9 a1 a3 a0 a1 a4 9b 9f 9b 9d a2 9f a1 9e 9e ab a0 a2 9f a5 99 9c 9c a0 98 9b 98 a0 a1 9f 9d 95 94 9b a4 90 9c 9c 94 96 98 95 91 97 8e 94 93 90 8e 8e 95 89 8e 84 7c 77 73 70 75 6e 6f 6e 63 70 63 63 69 67 67 68 5a 69 6b 62 62 5f 60 5c 5e 62 5e 68 6d 90 88 79 68 58 3c 28 1c 0d 07 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 10 22 34 3d 55 64 7d 7b 6e 71 68 6f 68 6a 70 6d 6d 6e 6c 73 76 73 6f 7a 7c 71 79 7a 70 7c 72 81 7e 7a 81 7d 89 8c 8a 88 93
 90 8e 94 92 97 9b 95 9c a1 9d a4 ac af b5 b8 ba c1 c0 d0 cf d2 da de dd e6 ee e6 e4 ee ef ea eb f1 ea f6 f1 f1 f5 f3 f1 f4 f0 f5 f5 ef e9 e8 ef e3 e6 e6 e4 ed e6 de cf d7 d0 d5 cd d9 e2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ff ff f1 cc b6 a1 a4 a3 a9 a5 ab a9 ad ac ac a6 af bc d3 da fc ff fd c4 a9 9a 9d a3 a0 9b 98 9e 9d 9d 99 9a 93 96 a0 97 9b 93 96 99 98 a3 9b 99 9d 97 92 91 9a 8f 98 92 96 95 99 9d 99 9a 8f 9b 91 93 99 8c 96 94 8e 93 90 8a 91 8f 90 8d 89 8e 81 7f 81 7e 75 79 77 75 6c 6a 69 66 6d 71 65 6e 6a 65 60 67 64 5f 5b 5f 5a 55 5a 5b 53 59 64 6f 83 87 7c 6a 50 35 22 10 0f 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 07 13 2a 2b 3e 55 64 75 77 70 6f 6f 71 73 68 6a 6c 72 6b 73 6f 6d 77 78 76 7b 7e 7f 7e 81 7e 7d 84 78 7f 81 86 87 8a 86 8c 8d 91 93 8d 94 99 92 98 9c 9d 9f a6 a6 af af b4 c3 c4 c5 d2 d4 d3 df e5 df ea de ea e1 ec ed ea eb f1 ea ef f1 e7 ef ee ec f6 ec ee ec e8 e6 dc e2 e2 db d8 da da e1 d9 d6 d8 c6 ca cd cd da ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 ef e8 e0 d0 d3 c8 b8 ae a1 95 9b 95 9a 96 99 9a 98 96 95 95 9d aa bb cf de ff f5 c1 a1 96 a0 97 98 a0 98 92 9b 9a 98 96 9c 95 91 92 9d 97 96 95 9e a1 95 92 9f 96 95 94 95 9b 96 8e 92 97 97 90 92 94 90 8d 98 96 95 91 94 8a 8d 98 94 8d 94 8d 8a 87 84 89 81 82 82 7e 76 7c 6f 75 6f 75 75 6a 74 66 68 62 6c 67 67 6b 66 63 5f 5c 5f 58 5d 5c 55 5a 63 6e 84 83 7b 65 50 3b 30 11 11 0a 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 05 06 17 23 2f 41 4b 61 77 72 7b 68 6a 78 73 6c 71 71 68 73 72 6a 70 70 72 73 75 7b 7a 83 7a 7e 81 79 7e 82 85 84 8d 84 86 85 89 92 91 8d 90 8f 95 94 91 96 a0 9e a6 ad b8 b7 c2 c0 bc d0 d5 d1 d5 dc de e9 e6 e1 e8 e8 e8 eb e5 e5 ee e7 eb dd e5 eb e3 ea eb eb eb e8 e4 e7 e3 dd da db d9 d7 d1 d9 d0 ce cf c6 c8 cb d9 ff ff ff ff ff ff ff ff ff ff ff f1 e5 df d0 cd bf b8 b6 ab 9f 9d 96 90 8a 83 80 81 7e 7e 8b 8c 86 86 83 8d 9e a5 b4 cc eb ed bd 94 8c 94 94 90 9c 8d 8f 94 8e 94 92 99 9a 96 93 8f 93 99 8f 91 8c 96 8e 92 90 8b 91 8e 94 95 91 93 93 95 94 93 8e 91 99 93 91 95 92 94 96 8d 95 8c 89 8e 87 84 88 84 87 7f 81 89 77 74 78 78 78 6e 6e 72 6f 70 73 6e 6c 67 65 65 64 64 68 67 59 60 61 61 63 64 55 5f 6e 81 84 7e 66 51 34 20 19 0e 07 05 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 17 1c 2f 39 4d 64 6e 78 67 6f 6b 65 69 6d 73 68 6c 6d 6a 6c 67 72 71 7a 75 73 7c 82 7d 85 7e 7d 84 85 7e 82 85 87 89 87 86
 94 8b 90 89 88 92 8d 97 9c 9f a6 a7 b3 af b6 bf bd c5 cf ce d1 dd db e1 dc e1 e6 e4 dd e8 e8 e3 e0 e4 e5 e0 e1 df e3 e0 e5 dd dc e1 dc df d8 dd d3 d8 d6 d4 d3 cf d0 be ca c6 b7 c2 bd d1 ff ff ff ff ff ff ff ff ff ff ea d8 c9 c4 bf b2 a6 9b 9a 95 8e 89 7b 77 71 76 61 69 6b 64 6c 73 6c 6d 77 7a 81 95 9b b7 d4 d9 ad 8f 85 84 88 8b 95 94 91 8e 90 89 8e 8b 8a 8d 91 8c 8a 93 8f 8c 8a 8f 91 8d 90 8b 8d 8e 8e 8a 8a 86 8e 90 8e 89 94 93 8f 8e 8f 8e 88 8f 8f 88 98 8e 83 88 85 85 80 83 85 7d 7d 7c 73 79 72 75 7a 76 72 71 65 69 71 67 6e 66 68 6a 60 68 5a 61 62 61 60 54 62 61 5d 58 6b 79 7f 74 5f 4d 37 2c 20 12 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 11 20 2a 46 4f 60 6e 76 6b 6d 6e 68 6f 73 74 6e 6f 70 6e 73 6a 72 71 6e 75 71 74 7a 76 7d 7f 7d 7f 85 7f 84 8d 84 8f 92 8a 8e 8a 8f 8d 8c 8f 94 97 9a 9b a5 aa a9 b0 b0 bd c9 c3 cd cd d0 d9 e0 db df dd dd e4 e7 e2 dd da e1 e4 dc e1 da d5 d8 d2 db d6 d0 dc d5 db d6 d0 d5 db d2 d1 c4 c3 c1 c1 b9 b9 ba b5 bf c6 e9 ff ff ff ff ff ff ff ff e3 cf c3 b8 a7 a4 94 92 87 78 71 6c 69 55 60 58 59 5c 56 54 56 59 66 6b 64 62 6b 6f 81 8f a6 cc cb a7 8a 82 83 84 95 8d 8e 8c 8f 8f 99 94 98 92 8e 93 8d 8c 8a 87 91 87 8c 88 89 83 8d 92 8d 8a 89 81 87 8c 86 91 85 81 93 93 8a 96 8e 8f 8a 91 95 88 8d 87 7e 81 81 81 7e 81 71 79 7f 73 79 79 72 78 70 76 74 6a 6e 6d 6a 6a 67 64 68 63 5f 66 5e 64 5d 58 65 5b 5e 5b 63 6d 71 83 77 62 51 3d 26 25 12 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 05 00 0c 10 22 2e 43 4a 5e 6b 72 72 67 69 6d 69 72 73 73 72 76 74 70 68 70 72 71 72 75 76 7c 82 7f 83 79 7d 79 7e 83 87 8b 8a 89 8b 94 8d 8f 8c 8e 8d 90 96 9c 9f a0 a8 aa b4 b6 b5 be bb c8 cc d0 d1 d8 dc d4 db e1 d1 d8 de d2 e5 e1 dd d9 e0 d7 d7 d6 d5 d9 d4 d7 d5 cc d0 cd d6 cd c4 ca c3 c8 c6 be b3 b7 af b1 ab b1 b9 de ff ff ff ff ff ff ff ed cf ba a9 96 82 82 74 76 6d 5f 5e 55 57 4f 47 44 4b 40 4b 48 4c 47 50 53 57 57 64 6e 7f 7f 91 b4 c2 9f 8b 85 88 89 85 8e 85 8b 97 95 95 92 94 96 89 8b 86 87 90 8a 8e 8f 91 7e 8c 80 78 80 83 82 89 85 8b 8b 8b 8a 8f 90 8e 96 8e 91 91 91 90 91 8b 8a 89 85 84 7f 78 83 7a 7e 82 7e 89 7b 75 77 7d 73 7e 76 73 6f 74 6e 71 68 6a 68 6b 62 63 64 56 5c 63 5b 61 68 5f 60 60 68 70 7f 78 62 55 3a 29 16 14 0e 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 12 06 12 24 2a 3a 49 5e 6e 6c 6b 64 62 6d 66 6e 6c 6e 75 78 74 71 71 6a 6f 74 71 76 7e 75 7a 7c 7f 81 7e 7b 82 85 84 82 7e 89 7e
 8f 8c 85 8a 8e 8e 95 93 92 9c 9b 9c a3 a9 ad b3 bf c0 c1 c4 d0 cd d6 d4 dc db d1 d5 d3 d1 d3 d2 d0 cf d2 dc d5 d2 d5 cd ca cd c9 d4 cc c2 c9 c6 c4 c9 cd c2 bc bd b7 b2 ae ae a6 a9 a1 ac d0 ff ff ff ff ff ff f2 d4 b5 a9 8e 7e 6f 6f 67 58 55 48 47 3d 40 3c 41 3b 3d 37 39 3c 40 44 37 3e 3f 4a 57 64 64 78 81 a9 b7 95 84 86 82 88 87 8d 95 95 93 90 8e 93 8a 92 84 83 8d 87 83 88 87 84 85 84 84 83 7c 7c 83 7f 84 86 87 83 87 85 8a 99 91 98 90 90 95 92 90 95 8a 89 88 85 85 81 7c 7e 7c 78 7e 76 76 76 75 7d 6b 73 70 77 75 6b 70 6d 64 67 6c 6d 68 68 5f 63 60 62 64 65 60 5a 5b 61 5d 67 71 7f 76 5f 49 39 1f 1c 11 08 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0d 0a 1a 1f 36 39 4c 5a 6d 74 72 64 5e 64 6e 6e 74 74 70 73 77 77 76 70 76 72 71 6d 78 72 76 70 78 7c 7c 7f 7f 81 84 81 88 94 8b 8c 88 86 83 8e 8b 88 8f 93 91 95 a5 a2 a4 ab b4 bb c1 b5 c5 bb c6 cf cb d5 d1 c9 cc d4 d1 d3 cd d8 ce d3 d0 d3 cd ce c8 c8 c5 c7 c0 c9 c9 bb c5 ba b5 bf b9 b7 b9 bb b0 ab a7 9f 9d 9b a6 c2 ff ff ff ff ff ff db be a6 88 72 61 62 51 47 47 45 44 3b 34 37 35 30 2f 2e 33 32 3b 32 32 3b 3c 3b 42 3f 4f 5e 69 7e 97 a9 91 90 85 8a 8d 90 a4 99 a0 9f 9f 96 8f 91 87 89 89 87 89 83 80 85 7f 7c 78 8a 81 82 79 7a 7c 7c 88 8c 87 90 8c 8b 8b 8d 98 90 91 92 95 90 8d 8a 90 8a 85 8b 84 8b 7d 84 7e 79 7c 76 76 79 7b 7b 7e 6c 72 71 6b 6f 6a 6b 6e 6b 66 69 6f 66 60 65 60 60 64 63 5a 63 5f 6b 67 76 7b 7a 5b 51 39 27 21 1c 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 03 0d 11 1b 25 29 41 49 5a 6f 77 6b 5c 62 66 64 6d 74 6f 76 76 7b 7b 6f 6f 72 6d 76 79 75 79 79 75 78 82 7f 7b 7e 86 84 7d 8b 88 84 83 86 8b 89 8c 8a 91 9a 92 93 9d 9a 9c a1 a8 aa b0 ba bd c0 c2 c5 cd c6 cc c5 cd cd d3 cc cb d3 c8 d0 cb c9 ce c0 bf c3 cb c4 c2 c7 c4 c0 ba b6 bb b3 b2 b9 b7 b3 af aa ae a0 9b 95 92 9c af f6 ff ff ff ff f3 d0 a8 8e 7a 73 4e 49 40 3c 3e 3c 33 37 35 39 32 31 2d 2b 30 2d 2d 2e 2c 28 33 41 40 3a 45 51 62 6f 96 a5 91 94 87 85 8f 9b a0 9c 9e a1 a1 94 8f 8f 88 87 87 8a 85 87 81 7d 7e 80 83 80 82 7a 80 79 81 86 83 8b 86 88 91 8a 85 93 93 8c 8b 97 90 8f 87 85 88 8d 8d 88 87 85 83 7f 79 7e 82 80 73 81 78 78 77 7b 7a 75 79 6b 6d 6f 6e 67 6d 66 60 66 69 62 61 60 6a 66 65 64 69 65 6d 7d 85 7f 63 4e 3e 2e 2c 10 07 05 03 03 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0b 21 2d 33 39 4a 5b 74 70 69 66 62 62 64 6e 6c 74 6a 72 7b 7d 76 77 70 70 76 73 6e 78 76 6d 6f 7d 79 7b 7f 7f 84 86 81 88 87
 8f 86 85 8a 8a 89 85 8f 90 98 9b a3 9d a3 a1 aa ae ab b0 b9 be bb c2 c7 c6 bc c7 cd c9 cb d1 c2 c8 c2 be ca c3 bc ba bd b9 b8 ba b5 af b0 b0 b0 ab ae a6 a8 ab ae a9 a6 a3 9b 9b 9b 93 96 9b ca ff ff ff ff f0 cb 94 71 66 5a 49 3e 2d 30 25 2c 2b 2e 25 2e 29 1f 21 28 23 24 2a 1c 2b 2c 2d 30 2c 2e 3a 4c 57 69 93 9c 8e 89 87 88 8a a0 9d 9c 97 98 93 99 90 8d 89 84 86 80 80 8d 7f 80 7f 77 86 87 89 79 80 87 7d 89 77 80 85 85 83 89 84 87 87 81 85 83 89 89 80 84 89 8b 8b 86 89 87 85 83 7c 79 7e 79 74 78 7f 7f 73 76 78 74 76 69 71 69 6a 64 69 6e 63 69 60 65 67 6b 63 68 64 64 65 62 6e 7e 7f 7e 64 53 41 2e 20 0e 15 05 03 05 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 0e 0d 18 2b 27 40 50 58 6e 6f 68 64 59 61 67 6d 74 76 76 80 7f 84 84 7a 72 72 71 75 75 75 77 78 75 7a 77 7a 7a 80 8f 7d 84 88 82 89 84 86 86 8c 89 92 97 97 90 9a 96 a1 9a a1 aa a6 aa ab b5 b9 b9 b9 b2 c2 c3 ba c1 bc c2 bc c5 c5 bf bd be bb b3 b0 b9 b9 b1 b4 b6 ab ac a9 a6 a3 a4 9d a7 a2 9f a6 9e 9f 92 9b 97 91 8c 95 aa ff ff ff ff ec e0 97 6b 59 4e 3a 30 29 30 25 27 27 1e 1f 23 20 20 1c 1c 17 1b 18 1d 1b 1f 22 1c 2f 2f 33 3a 4d 65 8c a0 8e 83 82 8c 88 91 96 94 98 92 90 88 90 89 81 8a 80 8c 80 86 7e 80 80 85 88 7e 7e 83 80 85 82 8b 85 7f 86 82 7a 7d 81 84 81 79 84 74 78 7d 77 7a 78 84 84 85 8a 8d 89 81 81 78 82 83 85 86 85 80 73 86 70 7b 6c 72 75 70 76 67 6a 6a 6a 66 67 63 65 5d 65 66 64 63 68 6c 6a 79 81 76 62 57 3f 2f 22 19 08 05 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 07 18 1c 24 36 3e 48 5e 6a 75 72 66 5e 64 64 68 6e 75 6e 80 8a 8d 8b 7e 77 75 74 6d 70 73 75 75 6d 73 74 76 77 78 84 7c 7b 82 84 86 81 8e 8e 84 8a 89 95 9e 92 94 93 95 90 a1 a3 ab a5 a8 ae b1 ab b5 ba b8 bc bc bd be c1 be bc c0 ba b9 bb ba af b5 ae b1 b0 b3 a1 a7 a0 9d a1 9e 9f 99 9a 98 9f a1 99 99 90 90 8f 8c 8c 87 9b e3 ff ff fa d6 b0 87 5f 46 43 35 2f 27 1d 20 21 23 20 16 19 1d 1c 18 1e 19 17 15 1c 1a 20 25 2e 24 28 25 3e 46 66 95 98 87 83 79 83 7e 85 90 87 87 89 85 94 80 81 83 7c 7e 83 87 84 87 83 83 83 80 81 82 8a 85 7a 7b 7d 7c 75 76 7d 6f 72 77 73 7f 72 6e 78 78 70 71 79 75 74 7c 7d 7a 85 85 84 86 80 8a 84 83 85 7b 7d 7e 78 7d 82 70 7f 70 6d 70 74 74 6c 61 6a 69 6a 6c 62 69 6a 6a 65 68 6c 78 7f 83 7d 62 5f 43 34 29 13 13 09 03 08 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 11 11 29 33 39 56 63 6c 78 6f 62 5f 62 64 67 6e 70 75 7c 81 84 86 82 81 78 77 78 71 6f 72 6f 75 76 72 75 7c 78 80 78 7e 7d 85
 83 81 85 87 85 8f 90 89 93 90 95 93 98 96 97 9b 9c 99 aa ae ac ab ab ae b5 b7 be b5 bb ba a9 b6 b8 b4 ab b3 a8 ac a6 aa b3 a4 a8 9e a0 91 a0 9d 9b 99 9a 94 94 90 91 94 90 8d 85 85 84 83 87 88 b4 ff ff de b0 8c 67 4b 36 2f 21 22 1f 1c 1a 19 12 1e 1a 09 17 0b 0f 0d 13 16 0a 0e 10 19 14 26 20 1c 20 35 4f 62 89 84 7a 76 78 77 75 81 7d 7e 7a 8c 81 81 87 80 7b 7f 7f 78 7e 82 7f 7e 7b 84 84 81 7a 7e 7c 7d 76 7e 79 7a 75 75 73 75 77 77 70 75 7a 70 69 72 6f 73 79 75 72 80 70 7c 79 83 8b 83 80 84 82 87 81 78 7c 7a 7c 79 79 70 73 6e 6d 6b 70 65 6c 66 67 66 6d 69 66 6e 69 65 64 62 72 81 88 80 68 5b 4a 36 1d 19 0c 05 03 00 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0c 20 29 34 3d 51 5b 66 7c 77 66 64 60 63 67 67 67 6b 79 7c 78 80 80 7a 7d 7d 78 73 7b 75 6c 76 76 78 75 71 72 78 80 71 7a 81 81 7c 86 87 85 89 90 85 8d 89 93 94 8d 97 99 96 9a 9c a2 a6 a9 a6 a9 ad b5 a4 af b2 b3 a9 ac b4 a9 aa a4 af a9 a7 a2 a6 a2 95 97 92 a1 94 92 8e 9b 92 8f 8a 85 8a 89 86 86 85 85 89 7d 89 82 81 8d ce fc be 86 60 48 35 28 22 26 1c 1a 11 15 10 10 10 0f 0c 0c 0c 0b 09 09 0e 0f 0f 13 0d 12 17 1d 17 1b 30 50 76 84 7f 7a 76 76 7a 71 76 77 7f 7b 81 7e 7b 78 72 80 78 7a 7d 7b 7e 87 77 7d 75 74 79 7b 7e 78 72 73 6f 72 7a 73 77 72 71 70 77 75 6d 71 74 6a 6c 70 6f 68 6c 75 72 78 72 75 7b 7d 78 85 89 85 82 7f 79 76 74 74 6e 73 74 6e 6b 68 6c 68 6d 6b 66 5e 65 68 62 6a 64 5a 5f 5f 6d 72 73 85 79 6c 5f 3e 33 27 0d 10 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 07 0b 1e 21 35 49 4a 5f 6a 76 7d 65 61 5d 66 66 69 66 6b 68 79 79 7b 7f 80 7e 7d 7c 78 79 7c 7d 77 77 78 7e 79 75 75 7c 7c 84 89 86 82 81 88 8c 89 82 8d 8a 8f 90 93 90 94 94 97 a1 9f 95 9c 9f a6 a5 a7 ad ab a8 aa aa a0 aa ab a7 a5 a7 aa a1 9a a0 9f a6 9b 96 88 96 9b 8e 92 92 86 88 86 85 7f 80 8a 79 82 7e 75 76 7f 7a 78 88 a8 de b5 70 4b 3c 2d 2a 1a 15 11 10 0e 13 15 0f 0c 11 0c 0e 0f 0d 05 08 0c 0e 0f 06 02 0c 19 1c 1b 25 28 52 6d 77 79 73 71 75 76 6f 76 73 7b 71 74 80 79 6c 72 75 77 76 75 73 82 6e 73 7a 7d 77 70 7b 6e 6d 72 70 75 71 74 6d 71 72 66 6f 6a 69 6f 74 6d 76 65 67 6f 72 6f 72 76 72 75 73 74 7d 7a 80 7d 88 85 89 84 74 76 72 78 6f 75 73 74 70 6f 5a 68 61 62 6a 65 64 68 66 64 62 5c 5e 66 6f 7c 85 83 6e 60 45 34 2b 1f 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 08 0e 1a 27 2f 3f 54 63 76 76 7d 6c 65 64 61 60 69 65 70 73 6f 74 78 77 7b 78 7e 7f 78 7e 77 7b 79 74 7d 7f 77 7b 85 7d 80 80 85
 85 88 8a 88 8b 86 86 8b 90 93 91 8f 91 90 8e 91 91 97 96 9f 9e 9f a5 a2 a1 a9 a2 9e a3 9e 9f 9f a1 a2 9e 9f 93 99 9a 91 9e 94 95 92 8b 8c 8b 7e 89 7e 83 89 7d 80 81 7b 7d 82 78 79 79 73 73 71 75 84 c0 ac 70 4c 35 24 18 1a 1a 12 14 0b 0a 13 05 05 06 06 07 13 10 0c 05 06 06 08 12 11 0f 16 12 15 18 2a 51 6b 77 6d 72 6f 6c 6c 73 70 78 74 74 7a 71 77 78 72 7d 74 73 72 76 78 71 73 70 79 69 72 6f 6e 70 6f 6e 73 72 75 6e 65 6c 60 6e 73 6f 69 72 6b 71 67 74 66 6e 6d 71 6b 73 76 6b 7a 73 73 7f 80 7e 84 7d 77 74 7d 74 70 70 74 73 70 70 73 6b 6e 63 69 65 68 6b 60 66 65 65 66 61 63 73 7c 84 83 6b 5e 4c 47 2c 17 0e 05 05 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 18 29 34 4f 52 60 63 77 78 68 66 64 63 66 5f 63 64 6f 6c 71 7c 6e 70 74 74 7b 74 70 76 73 75 7d 78 7b 73 6f 79 76 7c 7e 82 7b 7a 7e 84 86 84 87 84 7b 84 82 8d 80 8a 94 8b 91 92 8f 97 97 97 9b 9f a0 99 a2 9e a0 9f 9e 99 a5 93 92 91 91 8d 94 94 91 9a 8c 89 87 8f 7e 84 81 82 76 7b 78 80 73 80 76 73 73 7a 70 82 72 74 76 71 8c a2 67 44 30 1c 12 12 12 09 05 0a 06 09 05 00 08 09 05 04 06 09 04 0a 06 05 09 02 06 05 0c 12 15 2a 4d 63 6f 6b 6a 6b 70 74 76 6e 73 70 70 74 76 79 71 73 6e 6d 70 6f 73 73 6a 6f 71 6e 71 6f 65 6b 69 6f 71 64 6b 69 73 6f 64 60 68 68 6a 6f 6c 74 66 67 65 72 71 69 6a 63 6c 71 72 77 71 71 7d 74 7d 75 7e 7a 76 7a 71 78 72 68 71 67 6a 6e 6e 6c 6b 67 67 66 61 5c 66 5e 64 5a 62 63 77 7b 85 78 6c 67 4d 44 28 1a 0f 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 07 15 16 2b 38 41 51 5c 70 77 84 71 6a 67 67 5f 64 68 6d 6b 76 6c 71 6c 75 75 7b 73 78 76 77 74 70 74 6f 7c 77 72 7b 74 7c 7b 79 85 80 7a 80 82 84 86 87 85 8c 82 85 86 88 8c 89 93 90 88 94 93 90 95 97 9c 9a 93 9f 9c 9c 97 97 98 8e 91 92 91 8a 90 8b 8a 94 81 84 81 78 85 80 7a 82 7b 7a 75 75 72 73 71 73 79 69 6d 6e 6c 6b 6d 6a 6b 84 6b 44 28 22 12 10 10 07 0e 0b 0d 05 04 00 06 08 03 04 06 05 04 06 0b 08 03 06 09 05 0d 14 0f 25 43 62 70 62 71 73 6d 75 70 72 75 75 74 6e 72 6d 6e 6c 74 74 70 75 6d 65 77 68 6f 72 72 74 65 6a 6e 65 66 6a 6c 6f 6a 6e 67 66 6a 6c 79 70 6c 72 64 6a 6e 72 6c 70 72 6f 70 70 75 6d 6b 6a 72 7d 7c 7b 7b 77 71 71 71 73 76 70 74 66 68 66 68 6c 6b 67 63 64 65 61 5f 65 66 5f 67 64 71 7d 85 7b 6f 5f 4e 43 30 21 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 0d 18 23 38 46 58 5e 75 74 7a 7d 63 5e 61 60 6e 67 6a 6a 6c 77 6d 6a 71 79 76 7d 75 76 7b 70 70 72 75 79 71 79 7a 70 77 7d 77
 80 7f 7f 7d 82 7d 83 83 7e 8c 7d 80 87 8f 8a 8f 86 91 88 8f 8e 95 97 96 99 90 91 96 91 8c 95 97 88 90 8b 8f 8a 89 84 84 8f 7d 86 83 7b 80 75 75 7c 7f 71 71 77 71 6d 74 6c 69 6f 65 6c 6f 6c 71 66 67 6c 6a 5b 41 28 15 15 12 09 05 03 0d 0e 05 03 00 06 05 09 00 06 05 03 00 06 08 03 05 08 0b 10 0a 0f 21 43 65 71 70 67 67 69 6b 70 73 75 73 6a 79 6f 74 76 72 6d 76 6d 77 74 70 6a 6d 69 6d 6e 6b 65 64 6d 67 66 64 68 69 6b 6b 66 6c 6b 71 71 67 70 71 61 68 6b 6c 6f 6f 6b 74 73 6f 73 72 73 74 74 7c 79 73 7c 6f 6c 6e 73 7e 6f 69 6b 6c 6d 6d 66 69 67 5f 5f 69 64 5f 64 60 5d 5e 5f 64 77 86 85 7b 71 62 55 3d 38 16 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 1e 29 39 4b 56 65 66 79 7b 7d 61 61 64 5d 68 66 67 73 6e 75 6d 6c 6d 6e 7a 79 76 77 74 71 73 6a 6e 69 70 71 6c 70 69 76 6f 79 7b 84 7a 76 79 81 7e 84 89 7f 84 8c 85 89 89 84 8a 88 87 83 8f 8f 94 90 8f 8f 8b 85 87 8d 88 8e 88 82 89 84 80 83 80 7d 83 7b 7d 76 78 76 7a 77 74 71 72 6a 6b 73 70 6e 5f 6c 6b 66 6a 62 63 5f 66 5c 66 56 3a 26 0e 13 09 06 05 07 02 06 05 03 00 06 05 03 00 06 05 03 05 06 05 04 0a 06 08 0d 0a 12 16 36 5d 68 6e 6a 6f 60 6e 65 70 75 74 6c 70 6b 6c 6e 70 68 65 72 6b 6c 6f 63 65 6b 62 64 67 63 6a 6d 66 64 64 63 60 66 65 69 67 6b 6d 65 6e 66 68 6c 6a 63 6a 65 6d 70 71 66 64 63 76 6a 6f 7b 74 74 72 70 73 72 73 74 74 64 66 65 61 6c 66 65 71 60 63 66 5e 5e 60 5a 5e 64 5a 6c 63 76 83 85 84 66 5f 58 44 2c 1d 16 05 04 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0c 13 26 3a 4a 54 62 72 7b 80 79 6a 5a 5d 64 62 69 66 70 6e 70 72 70 6d 71 6d 73 71 72 77 6b 71 70 72 78 73 77 75 6d 70 72 75 75 71 74 7a 76 80 7d 7f 7a 7a 81 80 82 86 85 81 84 85 8e 90 88 8a 91 84 97 8a 8c 8b 89 89 82 87 80 81 88 80 84 7f 79 7d 7d 7c 82 7b 79 71 75 75 73 6c 71 6f 6b 69 66 60 62 6c 65 64 5d 64 69 64 58 60 5b 5a 52 41 2a 14 0a 05 06 07 07 04 06 06 05 02 06 05 06 00 06 05 04 02 06 06 03 06 07 05 03 04 0b 1c 3d 5e 65 6b 68 6b 63 6b 6a 6b 6a 67 72 70 69 67 66 6c 6a 73 68 66 5e 6b 70 61 66 66 62 60 5b 64 5c 66 66 67 64 60 66 67 6a 5e 64 6a 66 61 6e 64 5e 66 71 64 72 74 6d 6b 66 6b 77 66 67 67 6e 75 76 74 75 70 66 6b 72 73 70 66 72 60 6a 65 6b 66 62 64 65 6b 63 62 55 57 5d 62 62 65 71 7b 87 79 69 63 50 4b 37 22 16 05 03 01 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 09 0b 1f 28 35 4a 5f 63 71 7b 83 76 72 62 61 61 62 6f 68 68 73 6f 6f 6d 6f 74 76 76 70 76 74 6d 70 70 70 6f 72 79 71 79 6a 70 75
 73 73 78 79 7f 70 7f 77 7b 7d 80 80 7d 88 79 84 83 85 90 86 87 91 8f 85 89 89 83 83 85 8d 80 87 81 7e 7d 83 7b 7c 81 7c 7d 78 7d 74 73 72 75 74 77 69 71 6a 67 6e 66 6f 67 64 68 65 57 5d 64 62 5b 61 61 51 50 44 33 0f 08 03 06 07 03 01 06 06 05 00 06 05 03 01 06 05 03 00 06 05 0a 00 0b 08 04 08 06 15 34 53 65 71 6a 6a 63 6b 6c 6b 6f 6f 6f 6f 65 64 6f 70 6c 6b 65 68 67 6a 6a 66 65 64 69 5f 69 62 64 62 67 64 63 66 66 64 63 66 67 6d 6d 74 6e 71 69 64 70 66 72 6c 65 6b 6a 75 72 73 72 6e 77 79 75 6d 71 73 62 78 6b 6f 6f 6f 63 68 65 6e 65 67 62 66 5b 59 59 5e 5c 5c 5b 56 64 5d 6e 79 7d 77 6e 5f 5b 4e 3d 24 0a 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 07 06 15 27 33 47 58 61 6b 7a 77 78 75 5c 5a 59 5b 63 68 66 66 69 64 5e 62 6e 72 7a 70 6d 6c 6a 6c 69 6a 6b 66 75 70 67 71 6b 70 71 74 7a 74 72 75 75 79 83 78 83 80 7b 7a 79 86 7d 82 82 84 7e 88 89 80 83 7c 83 7f 87 7b 77 7d 7f 7b 7d 76 7b 6c 69 76 71 73 7b 76 73 6a 74 71 6a 6c 6a 69 5c 67 5e 56 5d 5b 5e 57 61 61 62 5f 65 66 5d 56 4d 44 2b 0b 0f 0b 08 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 08 06 06 08 12 2c 58 70 6f 6a 68 67 6a 6a 69 68 68 62 6c 6a 65 69 61 68 6b 6b 67 63 66 64 62 66 66 68 64 67 5a 5e 66 66 63 59 61 62 5b 5a 67 60 68 68 66 63 6c 63 66 6b 67 6b 6d 6d 6a 6b 68 75 66 6c 70 71 71 70 74 6f 64 6d 6b 75 73 65 6e 5f 69 68 64 6d 60 5b 5f 5e 5f 5c 5b 60 5e 5c 57 56 64 6e 7a 79 76 69 5e 56 47 3a 21 1d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0d 16 2d 3b 52 5c 69 70 7e 83 7e 7b 62 59 5b 60 66 64 66 69 63 71 64 66 69 6a 6e 68 73 6f 6a 6e 71 72 6f 6a 6f 6e 6b 70 70 6c 72 70 71 6b 78 78 73 76 77 79 7d 7b 75 7c 78 80 7e 7e 83 83 7f 81 88 84 7e 79 7d 7d 73 74 7a 82 7f 7a 79 79 71 73 6a 76 72 70 69 70 69 6e 6f 6b 70 64 67 69 62 5f 5a 61 5a 5e 60 60 5c 5b 5c 56 5c 5b 56 5b 50 4d 39 15 0d 09 06 05 03 01 06 07 03 00 06 05 03 00 06 05 03 01 06 05 03 0a 06 05 0e 09 0b 10 30 55 67 6e 68 6b 62 69 62 70 6c 67 66 66 66 6e 64 68 62 66 64 64 65 68 66 64 69 67 5f 64 61 5a 5e 5e 5f 66 5d 5e 67 60 64 64 6a 6c 72 62 66 6e 63 60 69 69 6f 6a 65 6b 5f 6b 66 6d 6d 6b 76 72 6d 6d 6d 6c 6a 67 67 6c 6a 6c 6b 68 6f 69 67 5f 5f 5b 58 57 5a 5f 57 5d 55 52 5b 60 6a 6f 7f 6f 5f 5f 4f 4f 39 27 19 11 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 0a 0f 1f 2c 41 43 54 70 72 74 84 86 74 6f 58 58 5e 65 62 67 69 63 66 6a 69 6d 6e 6d 65 70 6a 69 61 6f 6e 6c 6c 6d 71 6c 69 6e 6f
 6c 71 72 6e 76 70 74 7f 73 7d 7c 77 7a 81 85 83 81 7b 83 82 80 7b 79 7b 79 75 7c 75 6b 79 71 77 78 70 73 72 6a 6e 6b 6c 6a 6a 69 6c 70 6b 62 64 67 69 67 64 5f 5b 5a 54 5b 5d 5c 5e 58 61 5a 5d 61 58 5a 58 57 4d 32 12 0d 07 06 05 03 04 08 05 03 00 06 05 03 00 06 05 03 03 06 05 03 01 06 05 06 0b 0f 10 33 56 5c 68 5f 63 5d 6e 62 6f 6f 63 6d 66 6b 64 6a 68 63 69 62 5e 64 68 60 64 60 62 5b 61 65 5d 58 5f 61 6b 5f 60 5b 63 60 62 6b 67 71 61 63 64 5e 6d 63 64 66 6b 6b 66 65 6e 69 6b 69 6e 71 77 69 71 71 72 6b 6f 69 6f 67 6e 6f 69 60 60 68 6d 62 5d 5a 5b 60 5b 58 59 62 57 5e 54 61 6f 74 7a 64 5f 4d 53 43 2f 20 0e 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 17 14 2c 3c 4c 57 69 71 6f 81 80 82 72 5e 54 5d 5d 60 67 63 5e 65 66 65 69 6e 6c 60 69 68 66 6c 6e 6e 61 5f 6d 67 6e 70 6c 66 6f 69 78 6a 70 70 78 73 6d 74 6d 73 7b 7b 79 7e 78 77 83 7e 7e 76 7d 72 73 75 7a 6c 72 70 74 7e 78 79 69 76 70 6b 64 66 69 69 62 68 5d 67 65 6d 67 64 66 64 5b 54 5c 5c 57 5a 58 5b 57 5f 58 54 5e 59 54 58 4b 4e 2c 11 06 06 06 05 07 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 06 04 06 11 2e 47 65 5b 5d 65 5d 6c 68 5f 65 6c 6a 6f 65 69 61 64 6c 64 60 61 5f 67 61 67 62 64 61 60 5f 62 61 60 57 5a 62 5a 62 64 5d 61 6c 63 61 65 67 6b 62 67 6d 6a 69 6b 6b 66 6d 67 65 6d 6b 71 71 6f 71 6b 6c 64 68 6d 6a 74 69 69 63 68 5d 63 69 5f 5b 5f 5a 5a 56 57 55 5c 58 50 55 57 5f 69 72 6d 65 5d 56 4e 3d 2d 1e 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0b 1d 26 48 57 60 69 68 70 7a 7e 77 68 5f 4f 56 5c 60 66 6c 60 65 59 60 62 61 66 64 62 60 61 5e 65 64 64 69 61 6e 6d 6c 6a 6c 65 69 6b 68 6e 78 71 75 73 75 74 6e 76 78 7a 7d 71 7d 75 7d 6d 79 7c 79 7e 77 6a 6d 6d 6f 6b 67 73 73 6b 66 61 63 6a 5f 6b 69 61 5d 61 62 63 64 6b 65 61 57 59 59 56 58 57 54 57 5a 58 55 5f 5b 53 55 54 57 51 4f 34 14 08 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 2a 4d 60 67 5e 5e 5a 61 61 61 62 66 64 65 6d 6b 56 61 66 62 65 5f 60 5c 62 5a 5e 64 64 61 61 63 64 61 63 5e 5d 66 61 61 60 64 6a 68 68 67 64 60 61 69 65 66 65 60 68 6e 69 69 69 6c 67 67 66 72 69 6e 75 6d 65 62 65 6e 6f 73 69 66 62 64 61 60 5c 52 5d 59 58 50 57 57 55 57 4f 56 50 66 6e 69 64 5b 59 49 45 26 20 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 0b 13 1e 2a 3c 52 62 69 70 7c 84 7e 75 76 5d 55 5b 55 67 5d 65 66 66 67 66 65 62 62 68 66 65 5a 5d 59 61 65 6b 6f 78 73 70 68 67
 6d 6c 69 72 64 6c 75 6d 70 6e 70 73 72 73 73 77 7c 75 7b 78 73 74 7c 77 76 6e 6d 6b 73 68 6a 6a 6f 6c 70 74 6f 60 63 5e 69 5f 61 59 5c 5f 59 5e 68 5d 61 5b 5d 4f 5f 62 53 52 54 55 5b 5f 4f 51 4e 56 51 4a 50 49 37 10 03 03 06 05 03 01 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 07 06 09 0a 2b 4e 59 62 5b 62 5d 64 5f 6b 6a 67 6a 5d 64 64 6f 60 69 62 66 64 5d 63 65 63 61 6c 62 6c 6c 65 61 60 65 5c 61 5c 60 5d 65 65 67 65 64 6a 6d 6e 6c 60 66 63 6b 67 5e 6e 67 69 5f 66 6a 6d 6d 6e 6a 72 6c 65 67 6c 71 77 69 6e 70 68 74 63 67 60 5b 60 5d 55 5b 53 52 59 5d 58 57 48 4e 61 6e 65 60 5e 53 45 46 32 1d 13 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 15 1b 33 42 4a 67 61 70 79 77 7b 7e 76 5b 57 53 51 5f 62 5e 65 6a 60 67 66 65 62 64 60 64 60 66 5b 63 5f 5d 6b 71 6d 6b 65 68 6c 6b 6d 69 66 6a 67 71 6c 71 77 71 6b 74 6d 74 79 75 7a 6f 73 6e 73 68 73 6e 69 70 5f 65 6b 6d 6d 6c 66 64 67 5f 65 65 66 62 5d 5a 5d 5a 5b 5c 5d 58 57 55 56 5b 5a 5f 54 55 58 5a 4e 50 4b 4f 4f 53 55 4c 51 45 3a 0e 05 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 14 20 55 54 5e 59 66 5d 64 61 65 61 5f 67 69 68 6b 67 69 68 65 65 5d 5f 62 5d 60 56 6a 62 65 66 60 67 6a 66 68 5f 66 65 63 5e 60 64 65 68 64 6a 68 68 65 67 65 5d 61 63 6d 5f 62 60 64 60 62 68 68 69 6a 68 68 6b 6c 69 6e 70 69 70 6b 6f 5f 5a 64 53 59 5a 57 52 52 53 54 4c 4c 4a 49 4e 53 66 60 5b 5e 54 4a 47 2f 25 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0e 10 22 36 46 51 58 61 6f 6e 75 85 7d 76 58 49 55 55 5b 61 60 6c 5d 67 6d 66 65 63 61 5e 5b 57 5b 5a 61 5d 66 6e 73 65 6c 68 6a 69 62 6a 65 64 64 5d 6d 71 6c 63 6f 6a 6b 71 6e 73 6f 71 74 6f 71 6d 75 73 73 63 6e 66 66 6d 69 64 65 64 6d 63 66 5d 5f 65 58 5f 58 52 5c 58 5d 52 57 54 59 5d 5c 54 5e 52 55 4e 58 56 56 56 49 55 4f 45 54 42 44 30 14 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0a 0b 2a 51 5a 64 5c 5f 58 61 5a 65 5b 5d 61 6f 68 6b 64 6b 6c 6b 6a 5f 61 63 65 63 62 64 5e 5e 63 5e 61 5c 60 64 66 66 5f 6b 65 5f 62 56 66 60 65 63 68 68 68 5f 59 6c 64 63 5d 63 65 63 66 5d 6a 69 67 6a 64 68 63 68 69 68 69 75 6f 67 6a 62 67 5c 5e 58 5b 50 59 52 55 50 49 4b 42 3f 43 49 5b 67 63 5b 50 4e 44 3a 20 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 18 28 30 3e 58 5f 65 6c 6b 72 76 72 77 5a 4c 52 4c 57 5b 67 68 66 67 66 5e 62 5d 5f 60 59 64 5a 59 59 62 5d 65 6b 64 67 5f 65
 64 60 61 66 66 68 6f 67 65 6d 6e 6e 6f 6b 6e 73 69 63 6a 74 69 6d 74 61 6c 67 6a 66 68 61 63 68 64 63 66 60 5d 61 60 66 63 5b 5d 5b 52 62 55 58 5b 50 55 5c 51 55 4f 50 49 55 55 51 51 50 4a 4a 45 4d 54 47 49 48 32 10 0b 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 02 08 05 1e 49 5b 5e 65 5f 59 64 63 60 62 61 62 6b 68 70 63 69 65 69 65 65 6b 59 64 65 61 63 5b 5e 57 5c 62 66 64 65 64 6a 6d 67 63 64 68 69 71 5e 69 6c 62 67 64 6a 64 66 67 67 5e 63 62 63 65 60 66 60 5f 65 6f 6d 68 67 64 71 70 6f 6d 68 68 5f 5c 64 57 53 50 4f 58 50 4d 47 48 3d 4b 3f 46 49 5d 5f 5d 60 5a 4a 46 32 1e 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 03 12 1d 2a 38 3a 53 66 5b 6c 73 78 75 6f 64 57 4c 4e 52 4f 58 5e 5a 59 5f 65 60 66 56 54 5e 57 52 5a 58 5b 65 64 66 68 64 5e 5f 6c 67 6a 68 60 66 6b 6c 63 77 6e 62 6a 6e 6b 70 73 66 6c 6d 6f 6b 6d 6c 69 6b 62 61 64 62 64 65 62 63 62 5b 64 60 62 5d 5b 63 68 5b 5e 59 56 4e 55 57 52 55 4f 51 53 48 50 51 4c 52 4f 52 50 50 50 54 4f 46 50 42 3c 34 11 03 04 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 09 1e 4d 55 54 57 58 59 62 57 61 60 68 66 70 6a 64 64 68 5f 69 64 68 66 68 5e 5b 68 61 62 61 5e 61 5f 5b 5e 59 65 61 64 6a 65 6c 69 63 66 60 6b 63 57 5a 67 67 65 63 5d 64 66 58 5c 65 63 64 5f 62 62 69 66 6a 6b 62 6c 6c 69 6c 6d 66 63 60 62 58 57 5c 5c 4f 53 57 4a 53 4e 41 49 46 3f 45 49 64 5d 5f 58 4e 4a 38 20 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 05 13 1e 25 2e 4c 59 60 6d 6e 72 77 71 66 55 4e 47 53 49 54 57 4f 60 62 60 62 56 64 57 56 53 5a 5b 56 5a 59 52 5e 5f 64 5c 5d 62 5a 61 64 5a 66 69 62 62 65 66 6b 65 69 6a 6b 6b 66 65 70 66 6c 6b 6c 70 6a 6b 62 60 62 5d 60 63 5d 62 5f 5e 65 52 5f 60 5d 5e 5d 53 5a 52 57 51 59 57 57 51 50 44 46 4e 51 5b 50 52 49 50 4e 4b 47 4c 4f 49 4a 46 46 37 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 19 4a 55 5a 5c 5c 58 5b 57 60 66 60 62 6d 67 6c 68 69 70 66 5e 65 68 66 60 65 62 64 62 65 65 65 60 62 61 60 67 62 64 6b 68 64 65 64 6c 5d 65 65 5d 5c 62 62 62 64 5c 5e 5e 5d 60 64 56 57 5f 64 65 65 6a 64 62 65 65 65 60 65 66 60 61 50 57 5a 58 53 54 54 5e 4c 50 54 47 45 41 42 35 44 48 54 60 58 55 4b 3f 3a 1b 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 19 1b 29 3d 42 52 5d 62 6f 75 76 74 71 57 49 3f 52 4e 5d 52 58 5e 53 5f 5d 5c 5c 5b 58 57 58 50 53 5c 54 5a 60 5e 5a 63 5a 65 60
 60 62 5e 61 69 6b 64 6c 65 62 6a 6b 6b 6a 69 69 62 6b 70 62 68 70 6c 67 63 65 64 64 66 64 62 61 5c 63 60 5d 58 5b 5a 57 5c 60 59 57 58 55 4b 56 57 4f 4c 4e 43 4c 4d 46 4b 43 52 4e 4e 4b 4b 4b 4e 49 4a 5d 46 3c 38 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 05 06 05 03 00 0c 08 16 45 4f 53 56 5b 5e 5a 5d 65 66 67 66 6b 61 69 62 71 69 6b 68 65 66 68 61 64 5f 64 66 68 65 64 64 5f 6b 62 69 64 60 66 67 66 6b 64 6b 60 5b 6b 64 5d 5b 5d 64 5c 6a 65 59 5a 5c 67 59 5f 62 5e 62 6b 6c 63 68 6d 6d 67 63 60 62 65 5a 61 54 5b 56 54 5d 55 61 57 56 4a 45 42 48 3a 3f 3f 50 59 57 5f 57 46 42 31 17 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 14 18 1f 2d 36 40 4e 64 6a 70 71 76 6c 63 5f 4a 4b 49 47 54 58 54 5a 4b 53 61 59 60 58 52 59 52 54 58 51 52 60 55 5f 5b 54 59 60 60 5d 64 62 63 66 5e 5e 64 6e 69 66 69 6a 63 68 6a 63 6c 65 71 68 66 66 62 65 5f 67 63 5a 65 61 60 63 58 5b 60 59 60 5b 5f 63 5d 57 5a 4d 5a 54 4c 48 46 47 50 46 4b 4f 49 46 4a 4e 4a 4a 4d 46 53 4a 47 4c 4f 41 3a 32 18 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 06 14 44 61 5c 5a 5b 5b 5d 5c 69 61 65 67 71 69 6e 69 6c 75 6b 69 66 65 6a 5e 67 69 65 5d 67 62 5b 66 60 68 63 5e 64 67 6a 6e 67 6a 61 66 5f 60 62 5b 5c 62 62 5b 5f 61 60 60 5f 61 61 5c 5b 62 65 65 65 61 67 65 6e 66 6c 62 6e 5d 62 5a 53 56 58 57 58 5f 5a 58 56 47 49 47 41 48 35 38 39 40 54 5d 5a 56 4e 41 30 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 08 1f 22 26 3b 48 5d 61 65 6f 75 7a 75 65 50 4d 44 4a 4e 46 5b 56 4f 55 51 5f 60 60 5f 57 5d 55 4f 4e 59 61 4f 5b 59 5a 4e 55 65 62 5e 64 64 5d 60 63 65 5a 68 63 63 63 65 6a 6b 64 65 63 6b 67 65 6a 5c 66 65 66 64 62 58 50 5a 59 5d 5b 54 5f 55 52 61 5b 5c 60 57 52 58 49 50 53 4e 4c 4a 4a 48 4a 45 46 41 4a 4d 4c 4f 4a 47 42 48 4a 48 43 3b 39 2f 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 12 3c 51 59 5b 5b 5b 5d 58 5c 62 6b 69 67 6f 6d 65 6c 67 65 69 62 63 64 62 64 61 67 5d 61 5e 5e 5c 65 5b 5e 62 5f 5e 5b 5f 5d 5b 66 57 5f 5c 63 59 5e 63 56 58 5d 57 5e 5a 5a 5e 5e 5b 5d 63 5b 5d 69 65 6b 71 67 6a 6c 64 68 59 5c 57 5b 52 51 4d 55 5d 5a 56 57 4e 42 42 45 3d 40 3e 3f 40 52 56 5a 5a 4b 3d 29 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 04 0a 0a 0c 1f 23 2a 3b 45 52 5e 64 70 75 7d 7a 63 55 46 37 43 45 4e 56 52 54 56 55 59 58 5d 5e 5d 60 53 4d 51 54 56 4f 55 4d 5d 5b 5d 69 58
 5b 60 5e 58 6a 5d 67 64 65 71 5f 63 70 6b 6c 63 65 6a 66 66 64 60 66 5c 62 60 65 67 5e 62 5b 54 5c 59 5a 5c 57 59 5b 54 67 63 63 5c 5a 52 47 48 49 51 4d 48 46 3e 40 48 49 45 56 47 48 47 43 47 53 4c 46 41 49 3b 3a 13 06 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 11 3a 56 56 66 59 5a 5e 5e 63 6f 60 6b 6e 73 6a 6d 62 67 6c 67 6f 66 64 6a 5d 5c 61 63 5b 64 62 5e 5e 5d 64 67 64 64 60 65 61 59 61 59 5c 62 5e 5d 56 5b 64 5e 58 5d 5c 5d 5f 64 58 65 5e 5b 60 5d 67 66 6d 69 6a 64 64 5d 5a 5e 54 57 51 54 5f 56 59 5a 4c 57 4c 50 48 46 48 40 41 3a 34 43 51 59 59 55 48 3c 22 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 08 0b 0a 16 26 3a 3f 44 57 5e 67 6f 79 78 78 67 55 45 46 49 4b 44 51 4f 5a 5c 54 5b 59 59 60 56 51 56 57 4f 5a 56 5c 54 54 5b 58 57 5f 5d 5f 62 61 60 5c 62 5c 62 66 64 69 67 66 69 67 64 6a 6d 6f 64 61 62 5a 61 60 5e 64 5f 60 57 59 57 5a 5b 5b 5a 52 56 5b 5d 64 5e 68 5e 4f 51 4c 49 4e 3d 4e 44 55 4b 46 46 4c 49 4a 47 4a 4c 4a 4f 4f 51 4a 47 40 3e 31 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 14 38 60 63 5f 64 65 5f 5b 65 6a 64 68 6f 62 74 66 6a 6c 63 6c 6e 62 67 5f 6a 62 63 62 60 69 64 61 65 63 64 61 5f 66 5f 66 61 5b 5f 60 58 5a 60 51 4f 5d 58 57 5e 5b 5c 61 5f 5e 6a 65 61 64 64 69 64 6b 6d 67 6e 68 5d 64 69 55 5a 53 59 4b 52 50 59 5d 55 50 4d 56 52 43 41 3d 3b 3e 37 42 45 55 57 4d 44 39 2f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 09 11 14 2c 2d 40 51 55 61 6f 6a 71 72 74 6b 50 3d 46 46 4a 51 50 51 4f 5c 52 4a 5b 57 54 5d 56 54 52 52 50 51 51 53 57 5c 5c 51 58 62 5d 5c 5d 60 5d 62 5e 67 5f 63 6a 65 65 66 6b 66 6b 63 60 65 60 67 5e 56 5d 59 58 56 55 5b 5a 5d 57 51 52 54 55 54 50 56 64 58 60 5b 4b 50 4a 4e 4f 49 44 4a 45 44 48 46 46 47 4a 46 48 44 44 43 43 4b 48 46 40 40 31 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 30 64 5a 67 58 55 5a 55 65 65 66 6c 6c 6c 63 67 66 66 6d 64 5f 5f 5b 62 64 60 64 60 5d 5e 5f 5e 5c 61 64 5f 58 64 64 5c 5e 64 55 5c 56 50 5d 54 5b 5b 5a 58 57 5a 5f 56 69 5e 5f 62 5e 63 60 5e 6a 66 6d 64 67 69 67 5f 5f 55 51 55 53 54 4f 4f 57 51 4a 49 4b 4b 4c 40 41 3b 3a 32 36 3f 48 52 50 47 3a 2c 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0c 06 0d 1d 23 34 3b 45 55 62 6b 69 6d 77 7a 6a 62 49 45 4a 44 4a 5b 4f 53 52 50 4e 56 52 60 5a 52 55 52 57 51 55 4e 51 4c 55 52 5f 61 5b
 5d 62 62 61 68 5b 65 5d 60 67 61 62 68 62 5f 68 67 61 6b 62 6c 64 5e 5a 5d 5c 59 5f 55 5d 5e 5f 58 55 56 57 56 53 55 5c 62 61 5e 59 52 4b 46 46 49 50 4a 44 41 4b 41 44 43 45 50 46 45 4b 40 3c 3c 46 42 40 50 39 36 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 0d 33 5c 65 5f 56 55 63 5c 6d 65 66 6a 68 6a 6e 65 5f 65 5b 65 67 63 64 64 60 5c 62 65 5c 65 65 5c 64 66 5a 64 61 65 5b 5e 58 5b 55 57 54 58 5a 56 52 54 55 56 57 51 5e 62 64 5d 65 62 6b 65 60 62 69 65 60 65 65 63 5e 56 5e 56 55 54 54 4f 50 4f 50 4e 50 50 45 4e 4a 47 42 3c 36 37 30 3d 47 4d 4b 3e 3a 2b 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0e 14 1d 29 41 40 4d 5c 6b 65 72 70 7b 7d 76 59 49 3e 46 45 4c 56 50 54 58 57 4e 50 57 57 56 4f 53 4a 50 5e 54 4e 5b 57 5d 59 5f 64 64 5b 5f 64 5c 66 63 5e 60 5f 62 67 62 66 60 67 65 6c 64 63 63 58 62 61 5d 5e 5c 56 5c 59 4f 54 5a 51 4b 55 59 52 4f 57 5a 64 66 5e 5c 52 56 47 49 4d 4b 52 47 47 4b 44 49 50 44 4d 4a 4a 47 44 45 51 46 3e 47 40 39 29 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 0b 0f 2f 56 5e 69 62 5e 5a 5d 65 67 64 6c 73 74 71 6a 62 66 6a 63 62 5f 5e 62 65 6b 5e 62 63 61 66 58 63 62 64 67 62 66 62 5b 5a 5b 5e 59 55 59 5c 54 58 57 5b 51 53 61 58 5e 5a 61 5f 68 6b 68 6b 6b 6b 71 67 62 67 65 59 57 58 50 53 57 51 4f 51 50 52 4f 4f 53 4f 4f 4f 45 42 3d 36 34 36 3b 4a 3d 3c 38 28 20 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 0d 17 16 34 30 3f 51 56 67 70 73 7c 7b 80 77 5a 4f 43 4f 4a 52 56 53 56 5b 54 4f 55 52 55 56 54 4b 4d 4f 54 59 53 57 58 5b 53 5b 61 5d 58 6a 5e 5b 63 68 5e 65 69 67 5b 59 61 61 5f 62 66 5f 59 62 5f 5f 5d 63 5d 57 56 58 55 58 57 4f 51 58 4f 55 53 50 53 5d 5e 57 54 55 55 49 52 4e 52 4c 49 3d 45 4b 45 49 4b 46 4b 47 3e 47 4d 4d 3e 43 45 3e 4e 38 28 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0d 0a 26 56 62 61 61 5f 65 66 6d 69 67 6d 6d 6b 6a 67 6d 69 64 6f 69 5e 60 5b 60 65 62 66 66 62 5e 65 64 66 64 5d 65 59 60 5d 56 5e 55 53 4c 50 5b 53 56 57 47 4d 52 55 5f 51 56 5a 62 5d 70 62 68 62 64 6e 68 62 5e 5e 5a 53 53 47 4f 4b 52 4d 4c 50 4e 52 4f 4b 49 4b 49 44 42 37 39 35 37 36 3f 2e 2b 2c 25 1b 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 08 0a 13 22 2a 3a 4e 56 5c 69 62 6f 78 83 7d 78 65 4e 49 49 4a 51 55 53 52 4d 53 59 5b 54 56 51 50 50 57 51 55 55 54 55 59 56 59 5b 54 5f
 5c 5c 61 5f 5c 60 5d 61 62 60 61 5a 62 64 63 66 64 57 5c 66 5a 60 5e 50 60 4f 5b 4e 54 54 50 4d 57 53 51 52 47 4f 5b 58 58 62 5d 62 52 57 51 46 54 4f 51 52 55 53 53 4c 48 4a 47 47 4d 42 4a 49 48 47 45 44 45 3a 31 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 24 55 5d 69 62 59 63 65 6e 63 64 65 6a 72 6c 6c 61 6b 6c 62 5c 65 6a 61 66 56 64 5e 63 60 60 68 5b 60 62 63 65 61 65 5e 5a 55 5f 51 54 54 54 53 4a 4f 51 52 5b 4d 59 57 5c 5d 67 66 63 6f 6e 68 6b 6d 65 65 5d 54 56 4c 54 4f 4e 50 4d 53 47 55 3f 47 52 49 41 4c 41 36 3f 41 31 35 33 35 32 26 31 2a 20 10 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0d 11 20 28 35 4f 4f 68 6f 6f 6e 75 83 7c 7d 5d 4e 49 45 51 4f 4c 52 54 57 4d 56 5b 53 53 52 53 53 50 56 55 54 53 54 58 55 53 5c 5d 5b 5e 62 62 5c 65 67 6c 5f 63 62 64 63 61 64 59 5b 5e 6a 66 61 5a 5c 59 64 57 5b 5c 52 52 57 52 55 4e 54 56 54 52 58 5a 5c 60 5e 64 5c 5c 5d 51 54 5a 50 56 55 58 5e 51 51 51 52 4d 4b 49 44 45 47 43 44 45 42 40 3b 34 10 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 29 4a 59 63 64 62 63 64 6f 6b 6b 6b 6a 6a 73 64 69 67 65 66 60 63 61 5e 61 5e 69 61 60 64 5c 64 67 66 5f 5f 60 59 60 5d 60 5a 5c 5c 56 57 51 4f 52 53 49 54 4d 5e 56 55 5f 5b 62 61 6d 77 77 72 68 6f 65 68 67 5c 5a 49 56 50 4f 48 4b 48 4a 48 47 4a 4d 4b 4d 46 47 45 47 46 3b 3a 30 35 2d 2a 25 1a 1a 14 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0f 15 1d 33 3e 4c 53 5f 6a 6d 79 7b 81 77 7d 63 58 42 4a 49 4f 56 56 54 53 51 52 57 56 58 51 53 55 55 4f 55 52 54 5c 53 57 58 51 57 59 59 58 61 5d 5a 64 5a 60 65 6a 64 5e 5f 60 63 5d 61 5d 60 5e 57 5c 5c 60 53 4c 56 4f 4f 49 50 54 56 55 4c 52 4f 5f 51 64 61 5d 5a 5b 59 5a 58 58 59 55 58 4e 50 51 51 53 4d 48 4e 47 47 50 44 42 41 46 49 44 40 40 2a 11 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 01 06 05 03 16 52 5d 64 5f 62 64 62 67 66 6a 6c 6e 71 6c 6a 63 64 68 64 61 63 66 65 65 5b 68 5e 6a 66 56 65 5f 65 67 63 5f 5b 62 5c 5c 5a 4d 59 53 59 51 4f 50 4f 50 56 4f 51 49 50 5b 5d 61 63 6f 7c 77 6a 63 62 68 5e 58 5a 53 53 4c 54 4c 4e 4b 4b 51 46 4d 4f 4a 49 49 48 43 45 41 40 3a 38 31 2e 31 2c 26 1e 14 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0e 18 1f 36 38 48 58 60 66 68 79 75 80 81 77 6a 4e 4b 50 3f 47 4e 4e 4d 55 59 57 4c 55 4e 49 5c 4d 52 4b 4f 54 53 59 55 59 5c 56 53 58
 57 65 5e 5f 55 5e 5b 56 5f 5b 5c 62 61 53 63 60 5a 5f 60 66 5a 5b 5e 56 56 5c 50 4a 52 50 4d 50 50 4c 52 52 4d 58 5c 58 5e 5c 5d 61 4f 58 50 54 4a 46 52 52 47 4f 52 46 4b 4d 4f 4d 46 4a 44 43 45 42 42 44 3a 40 32 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 1a 4d 5e 68 66 68 65 6a 5e 63 6a 6c 71 6e 6b 6a 72 67 68 60 69 5c 66 5a 6a 5f 65 5c 64 69 60 69 63 61 68 57 60 63 5b 62 52 5d 57 55 55 5b 50 4e 4e 50 54 52 53 4c 53 52 5a 5c 68 62 65 74 75 6a 66 5a 59 5e 5b 5a 53 4c 4f 4b 47 50 51 46 47 43 48 49 4a 46 4e 43 3f 41 3e 39 3c 36 33 26 2e 1f 24 14 09 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 10 23 32 3c 4c 54 64 70 6d 7d 7b 82 86 84 63 4e 48 41 49 4f 50 4e 58 4f 5c 52 4f 4c 4f 55 57 51 53 53 46 58 51 4d 5b 57 55 55 59 61 57 62 5c 59 5e 5f 64 5e 58 5a 5b 59 5d 68 5f 61 58 5e 5d 5b 5a 56 58 51 5a 56 4d 55 51 4e 50 55 51 58 4b 4b 4a 58 5a 5e 61 59 5c 60 48 4d 4f 42 4c 4e 4e 45 48 43 47 4c 4d 45 4e 42 51 45 4a 46 48 4b 4a 49 48 41 2c 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 15 3f 62 65 68 65 68 6a 6a 6b 64 6c 6a 6d 70 66 65 62 64 68 63 62 6d 61 6f 68 64 67 64 64 64 5d 62 60 64 57 5d 61 5b 58 60 53 5e 60 55 54 56 51 53 55 4e 4f 57 52 57 5c 5c 57 59 61 6e 6f 74 61 5d 5a 60 5f 5b 5d 51 4d 4c 4f 4e 4c 55 43 52 49 48 4e 45 4d 49 41 49 44 48 3f 42 3e 32 2e 28 25 1d 10 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0d 1d 20 35 54 5a 69 71 6c 79 7a 87 88 81 66 59 4b 4c 4f 4f 55 5b 5c 4f 53 52 4d 58 57 53 50 4c 51 53 50 54 57 4b 4e 51 5b 58 5d 57 57 5b 5e 61 5a 5a 5d 61 5e 61 59 57 60 5b 5f 5e 5a 60 5b 5b 56 55 5f 4e 56 56 4f 54 51 48 53 54 4e 53 53 50 4b 56 5d 59 57 4f 55 55 58 50 4d 4c 48 46 4a 53 4c 4f 4d 53 49 43 52 44 41 4c 52 4e 4a 45 47 42 40 43 32 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 49 60 63 6e 64 68 62 67 6f 69 6e 65 6f 69 70 6f 6e 6b 5f 64 62 64 67 60 63 64 65 66 62 5d 5f 5d 5a 5f 69 60 64 5f 5c 55 56 4b 58 53 50 5d 45 54 4e 4d 54 53 52 55 53 54 5d 60 64 6b 71 67 60 5f 60 58 54 57 57 4b 48 54 4c 47 4b 52 4a 47 45 4a 4e 41 4b 49 43 47 41 43 3d 3f 3e 2f 30 28 18 1c 0d 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 07 10 1c 21 3a 40 4f 62 6a 65 70 7c 84 82 78 6c 4c 41 4c 48 4a 48 58 55 52 5a 4f 51 54 4d 54 4b 4c 4e 47 50 50 54 57 51 52 5b 58 58 58
 5e 59 56 58 55 5b 5a 5d 57 5c 53 63 59 58 58 5f 55 56 5a 58 56 53 58 5a 5e 56 4b 50 4f 51 50 51 4d 49 43 56 54 53 55 58 61 44 5a 49 44 4f 43 4b 46 41 4a 48 42 4b 48 46 4d 47 4a 48 46 47 3e 47 49 49 43 44 3e 40 2a 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 40 5b 64 61 5d 64 62 6b 69 6c 6d 6e 6d 6c 66 70 68 6a 6a 6d 61 68 69 6a 5d 5c 63 64 5f 5d 5e 65 68 64 5f 5b 5e 5b 53 59 54 56 51 4b 50 4f 4c 4f 52 52 4c 52 56 54 51 5a 5b 5c 63 60 64 6c 57 52 58 57 5a 51 47 4d 45 4d 47 4e 47 4f 43 53 3a 48 43 43 48 4e 44 48 3f 42 40 3d 34 2c 2f 2d 14 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 1b 26 36 3e 50 5f 68 69 7a 79 80 86 83 65 55 42 4d 44 4f 4b 50 57 59 4f 55 54 54 55 4d 48 47 4b 4c 4e 54 50 50 4e 55 56 59 5a 5d 57 5f 4f 5b 60 54 62 5a 5d 59 56 5b 58 59 62 5c 52 5a 56 54 52 51 52 55 52 54 59 51 51 4e 45 4d 4f 4f 54 53 52 56 59 52 56 52 4e 4a 44 50 50 4c 4b 4b 42 51 4e 42 4c 4d 45 47 46 49 3e 48 47 4f 44 43 49 46 44 46 35 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 46 5d 6b 6a 67 6a 6a 6c 68 63 62 6a 69 70 6e 68 68 67 66 62 63 67 69 6c 65 69 5d 63 5b 64 5f 5e 5b 64 67 62 62 51 54 5d 54 52 56 51 54 51 46 49 4a 50 55 54 4d 55 5a 5b 5d 62 62 60 64 64 66 5b 5e 54 52 4f 53 54 4e 49 50 4e 46 45 52 4a 3f 44 45 4a 4d 46 4a 48 3d 3d 3c 34 34 2d 2e 24 1e 12 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0e 13 23 33 31 47 5d 62 64 72 72 80 7c 7d 6e 53 4a 48 46 45 4e 48 4d 4f 4c 51 4d 4f 51 4f 50 4c 46 4f 50 50 56 55 50 53 56 50 55 55 58 5c 5f 54 52 58 59 51 52 5b 55 55 5b 5f 5a 54 58 5a 59 57 55 54 57 52 4f 52 51 4c 46 49 52 4e 53 4b 51 50 54 5a 5e 5b 56 4e 4d 49 45 4a 43 44 4a 47 4a 46 46 4c 4d 50 48 49 4a 48 44 4f 4b 49 44 46 49 43 40 42 31 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 45 57 62 70 62 67 60 60 66 6c 69 6f 6a 6f 65 65 6d 6a 62 6c 6b 70 6a 69 66 64 5c 61 59 62 62 5e 57 63 6d 69 68 5c 54 50 54 51 52 4f 52 48 56 50 4c 52 50 52 57 52 5c 60 61 61 5f 5d 61 63 60 62 5d 4c 4a 50 51 5c 4e 51 48 49 43 50 4e 51 4c 40 44 40 46 47 43 4c 43 46 41 3b 3d 2b 27 25 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 10 15 2f 2f 46 5a 5c 67 6a 7c 76 81 80 65 49 3c 3f 48 4b 4f 4b 54 48 51 46 4e 49 4d 55 4c 4f 4a 4a 51 51 4e 52 5a 5e 5b 58 5e 58
 56 54 54 53 56 50 54 58 56 55 56 53 51 59 52 59 5e 58 51 58 50 51 54 54 5a 50 4f 44 49 4d 4c 48 4b 48 49 52 57 5f 4f 54 50 48 41 46 41 46 3e 46 4a 49 48 4b 43 4f 4a 4b 45 43 4e 4b 53 49 4e 4f 45 48 53 4c 41 45 39 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 3e 64 67 67 6d 6a 64 65 6a 66 6a 6c 70 6d 6e 60 67 64 6a 73 79 78 76 64 66 68 5a 66 5f 64 60 5c 5f 65 63 65 68 65 52 53 4c 4e 50 4c 52 4a 4f 4e 52 54 53 57 55 57 5d 5b 59 64 5f 5c 66 62 5e 5f 55 4d 50 50 49 4b 4a 47 40 48 4d 46 46 44 3f 44 4c 3f 44 43 4d 3c 4a 4b 3c 3e 34 2c 2b 19 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 11 1a 27 31 3b 4d 52 60 6b 75 81 80 79 66 4a 46 41 44 48 48 52 48 4b 4d 50 5a 4c 51 51 4b 52 4d 4c 55 50 51 54 55 5a 5b 5b 55 5b 5d 5a 5e 55 5b 54 58 60 52 5c 53 53 59 5b 4b 54 5b 54 60 57 4e 50 51 51 53 5a 49 54 4b 4b 50 4f 52 5a 55 58 4f 54 51 4f 47 46 44 46 40 44 47 4b 51 4b 4d 50 4a 4b 47 41 4a 46 3f 4d 4b 4a 4b 49 4c 48 53 59 4c 46 3c 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 3a 5a 6b 69 68 63 5b 68 68 65 6d 73 71 76 69 6d 70 66 70 69 75 74 71 6f 66 67 61 5f 5d 5d 58 5b 51 55 54 5a 6b 68 60 5f 53 57 50 54 57 49 4a 4e 4e 51 5c 59 5c 5a 5e 5d 5f 5e 60 5a 62 57 57 5a 58 4e 53 4f 4e 50 48 4c 4b 4c 52 4b 45 46 46 42 4a 45 4d 4d 49 42 43 40 40 44 35 31 28 1f 09 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0a 19 19 2b 2f 46 4e 5c 69 68 72 7f 72 5d 4b 44 46 4b 4d 53 50 4e 44 54 48 53 45 4b 52 55 48 48 4d 48 52 53 54 55 51 52 55 53 59 56 5c 58 54 56 51 57 4f 5e 55 4b 53 52 56 4d 57 55 59 55 5a 55 5a 54 52 48 4d 53 53 53 4b 4e 54 4c 4e 59 57 5a 5d 4c 47 4d 42 49 44 46 46 4b 4f 47 4b 42 48 4d 50 4b 4a 4e 4f 56 4b 48 4e 49 4c 4d 49 4c 4e 48 3d 37 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 3b 62 6a 71 63 69 5c 68 6d 6c 64 6f 73 69 6a 6a 6f 6d 62 6e 74 75 6b 72 67 68 61 62 5e 61 57 59 5f 56 55 5c 5e 57 5f 58 56 55 52 52 4d 5b 59 50 59 5e 59 5e 63 53 5b 60 62 66 64 65 5c 53 53 57 59 4d 4e 50 4e 44 49 49 4c 46 44 51 4b 51 49 50 49 4b 4e 4b 47 47 44 44 42 3f 36 2b 18 18 14 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 13 1c 22 31 32 4a 4b 54 6b 74 77 71 60 45 3f 44 47 4a 4c 45 50 3f 3c 44 46 4c 4e 41 4d 4a 47 47 48 4f 52 51 53 5e 4b 4b 50 56
 50 5b 52 52 55 59 52 58 55 54 4a 57 4f 46 54 53 52 53 54 54 59 4d 58 50 53 47 4b 4c 4a 4f 5a 54 53 52 52 5b 4e 50 47 44 4e 3b 40 45 4b 4d 49 4d 4d 44 4a 47 47 4d 4b 47 4a 3d 47 46 42 49 4a 46 47 47 4c 47 47 3d 3a 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 32 5a 67 63 67 61 58 61 66 65 6f 70 63 71 6f 65 67 61 6c 6a 68 6f 70 65 65 64 5b 64 5b 5e 5b 57 58 59 54 5d 54 59 59 5b 52 52 4a 54 54 50 53 53 5e 63 5a 5c 55 58 4c 5a 59 59 5e 5b 5a 63 51 51 57 48 4f 4d 4d 49 4d 48 53 47 48 51 4a 47 49 44 43 47 50 48 4a 42 46 45 3d 3d 33 20 22 10 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 19 1a 26 2b 31 47 4a 61 6d 71 65 4e 43 45 3b 4a 46 4a 43 49 4a 4a 4b 46 4d 52 4d 44 47 56 4c 4a 53 4a 52 54 57 56 58 5a 56 57 51 50 54 49 50 4d 51 55 52 51 52 4f 53 44 51 52 47 52 50 51 5c 4e 55 4e 54 4e 50 4b 56 57 57 53 58 54 57 4a 45 49 47 43 49 50 46 42 45 42 46 4b 45 48 49 48 44 44 43 48 4f 4e 48 41 47 3e 4b 48 4b 4b 3c 42 40 34 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 35 59 68 60 5a 67 5f 6b 6b 65 6d 6c 6d 6d 66 69 6b 69 6d 68 64 67 63 6a 5d 62 64 64 5a 62 53 5b 55 51 4c 59 51 59 58 5d 58 58 56 4e 51 4d 4d 50 56 55 59 59 56 53 5a 59 56 5e 5c 5a 62 59 54 52 50 4c 51 4e 49 43 4b 41 45 53 46 4b 4b 42 52 49 43 44 47 49 44 44 3d 3e 42 38 34 1c 17 12 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 10 17 1c 25 31 3a 43 5a 64 63 68 4f 46 42 46 43 4d 4a 4e 47 4d 4d 4e 4c 47 47 52 52 47 4d 42 49 51 51 53 58 5c 50 54 52 54 57 5d 59 53 50 4d 58 54 4f 5c 57 51 4d 51 4b 46 4b 53 4f 57 53 58 5e 56 5c 4a 4b 4d 57 50 59 5f 59 60 53 59 50 4e 44 4d 44 4e 46 4b 4a 44 48 4b 3f 4e 4d 41 43 47 47 47 44 47 4d 4b 45 49 47 44 44 44 44 47 42 45 37 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0f 28 5a 6a 63 5d 64 5e 6a 6f 74 66 70 75 72 6c 6f 76 6d 6e 72 6a 66 6b 66 63 66 61 59 66 63 59 5c 5e 5d 51 55 57 56 55 55 54 55 56 56 56 5f 58 52 5f 55 5a 5a 56 51 4c 55 55 57 61 5e 5d 5f 55 54 54 50 51 4f 4f 4d 50 51 58 58 49 4c 41 51 4e 4a 4e 52 43 4c 4e 49 4c 3b 40 35 27 1e 10 0b 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 11 14 26 25 2e 43 50 54 5b 4e 4a 43 3f 47 41 42 4b 49 40 4e 49 4d 49 4b 4d 4b 49 4b 49 48 4d 44 47 4c 51 5c 4d 4e 4b 54
 58 5f 53 50 55 4c 51 54 51 52 49 52 54 4c 4d 4e 44 51 4a 55 4c 57 56 52 4f 46 4c 52 44 4a 53 5d 58 5a 52 4b 50 50 3f 4c 46 4a 4c 47 48 45 41 37 4c 41 45 4d 46 46 47 4a 49 48 39 3b 3e 3d 41 45 49 41 40 3a 3e 43 32 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 25 63 62 70 6b 66 68 6e 6a 64 71 6c 6f 71 6e 67 6d 60 6a 6c 6c 6c 68 62 5d 65 5a 61 5d 60 61 59 58 56 57 50 57 55 5d 5c 56 52 55 4f 57 55 51 52 57 58 54 54 52 4e 51 48 55 54 5a 5b 5d 60 5a 50 45 4b 56 51 54 49 4c 47 4b 53 50 4e 4d 4c 46 4a 52 43 48 4b 4e 4b 4b 3c 3b 36 2e 17 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 11 18 22 2b 33 45 53 59 4f 44 45 3c 47 45 44 48 3e 49 44 48 4e 47 50 4d 4e 4a 55 48 4c 4c 4a 43 50 4a 53 52 55 5d 52 4d 55 4a 54 52 52 4f 50 52 54 4d 49 49 49 4d 4e 4e 49 4f 4d 51 4d 51 4b 50 46 4a 49 4b 4a 48 4b 58 5f 5a 5f 54 4d 48 50 48 4b 4b 37 40 42 3c 46 40 3b 3f 4a 44 47 42 45 3f 4b 47 40 3f 42 48 3f 3e 41 45 3c 3a 33 34 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2d 57 6f 6f 66 66 62 61 6a 70 6c 69 6b 69 72 6a 6d 6b 6c 6a 6a 67 6b 61 62 60 59 5a 66 5a 5a 5c 59 5d 59 56 61 5b 58 56 5a 58 56 51 5b 4f 4e 51 59 53 56 51 54 55 52 56 55 54 52 54 5f 56 57 57 59 45 45 46 4f 47 48 52 4c 4a 4d 4b 4a 51 49 4f 4a 49 50 42 49 45 43 40 37 31 1d 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 1a 25 30 38 48 50 52 49 3a 43 3e 45 3e 4b 44 4e 3f 47 43 45 4b 45 47 4f 49 46 47 4a 4e 4f 59 52 4d 50 47 53 5c 50 54 5a 55 50 4a 49 46 4c 45 55 49 4b 52 4a 51 46 48 4d 53 4f 4f 50 4e 52 4c 4a 52 4b 51 4f 41 4e 52 52 5b 5b 4f 51 51 49 49 3d 40 40 44 3a 41 43 45 46 44 3a 44 4c 4f 43 4a 4b 45 48 47 46 41 45 36 3f 40 3a 36 43 2d 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 29 5e 6d 6a 70 64 61 6a 6e 73 72 73 67 66 6c 71 71 6e 71 6d 67 6c 62 63 5b 64 62 5f 56 5f 5a 57 64 54 56 59 54 54 56 5b 5a 4e 53 50 57 50 52 59 4f 5d 58 5a 52 50 49 50 51 56 5c 53 55 55 53 52 54 4a 4b 54 53 55 48 4e 4d 49 51 58 4e 54 47 4e 47 4d 4b 4f 4a 46 42 39 3c 2f 1f 0c 10 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 12 1d 28 30 48 50 50 49 3f 3f 41 48 3f 4a 45 4c 49 40 40 4b 44 4d 4d 51 51 4b 4b 4d 51 51 53 4a 4a 4a 4b 50 51 54
 4f 57 51 4d 52 50 4e 4e 52 45 4c 46 4d 52 45 45 52 49 49 46 4e 50 4a 53 53 4b 44 43 4b 48 42 4f 52 55 53 58 46 50 4f 45 4a 3c 41 40 47 39 3c 3f 43 47 3f 49 41 42 47 3d 49 46 3d 3c 3e 4d 41 3e 40 47 3c 3e 35 38 31 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 22 5c 64 6f 72 6e 62 73 76 66 76 6e 78 6e 6c 6e 66 6a 64 5f 62 5c 5d 5b 5b 5e 53 5c 56 60 5c 5d 59 52 56 5a 55 5c 57 58 56 55 57 56 52 53 4e 4d 55 59 52 54 4d 4d 54 52 56 50 53 50 51 5e 53 58 53 55 4b 50 4d 44 45 49 4d 46 4c 51 4b 4c 47 4c 4a 4a 4c 4c 47 43 3a 42 31 2a 18 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 0d 1f 22 2d 3d 4f 49 49 3d 43 39 3d 47 49 48 50 4c 46 4a 4b 4a 4a 48 4f 4e 4f 49 53 4d 48 50 47 4d 51 52 57 54 46 4e 51 4d 44 4c 4c 4a 44 48 49 4f 42 44 46 40 4b 49 49 44 44 4a 49 55 45 4e 48 4b 46 4a 49 47 51 4e 4c 56 50 59 52 50 44 49 3c 44 43 35 3a 3b 41 3f 43 38 34 3f 3d 41 43 40 44 3e 42 36 42 45 45 3f 39 37 37 35 38 29 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 21 58 68 69 6f 69 6a 73 6b 6f 69 72 68 6d 6a 6f 6b 66 6a 6f 66 68 62 67 5c 5c 58 55 5b 5a 54 58 5f 5f 5b 5b 59 54 50 5d 55 5e 55 52 57 59 53 4d 55 55 50 49 46 49 50 52 51 57 4f 51 4d 55 55 59 4b 46 4c 4a 46 4c 48 51 55 54 56 4e 50 49 4d 50 53 4b 4d 4e 47 46 41 34 31 1c 10 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 15 26 26 35 4d 52 4a 3a 41 45 3e 3c 43 4c 4b 45 45 42 47 4d 4a 4a 51 4d 4a 46 42 51 4c 4d 4f 48 49 51 53 50 4e 54 51 4c 4d 4c 50 47 51 47 4a 45 46 4a 47 41 42 4a 45 4a 44 44 4f 48 52 4c 4c 4a 41 41 4f 43 4a 49 41 47 57 59 56 53 3b 42 45 45 44 3b 42 36 3f 3e 36 3e 46 3b 3d 47 3d 3f 3b 46 43 3b 3f 3b 3c 39 41 3f 42 3c 35 32 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 53 6c 68 75 71 72 70 72 75 6a 72 6d 6c 6c 65 68 67 66 69 5f 5a 63 5c 57 5f 56 5a 55 64 53 62 61 5d 61 5e 5c 5d 51 59 58 5e 58 5c 58 52 51 56 57 53 4c 50 4d 54 55 53 51 4e 4e 4d 50 58 52 59 50 50 4d 50 48 4a 4e 4e 4f 49 54 53 4a 53 4d 4f 4f 4f 51 4b 4b 47 35 3d 21 1f 12 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 10 1c 2f 38 41 46 46 41 47 42 40 49 44 4b 54 45 47 4d 48 47 4c 4f 4d 4a 43 4d 49 50 55 52 4c 53 50 4c 4b 4b 4f
 4c 50 51 4b 4d 4a 4c 4d 46 49 45 4b 4b 45 43 3d 4b 43 3f 47 41 44 3c 44 45 4a 4a 51 45 45 43 43 48 45 42 4c 4f 4b 45 43 4a 3d 40 47 43 34 3f 3f 3e 3f 3d 45 3a 41 48 42 39 44 42 45 40 43 3d 40 3f 48 41 36 3c 37 38 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 25 52 67 6e 6f 69 65 6d 74 76 72 70 66 68 68 61 6b 65 66 66 64 63 5b 57 5c 5e 4f 5b 64 59 5e 57 55 60 54 57 61 59 63 63 63 61 61 5f 5f 5c 54 4b 59 55 4c 50 4a 55 56 55 4a 58 52 4e 59 54 54 51 4f 4c 4c 50 48 4d 4d 55 4f 50 52 54 4f 4d 5a 4f 48 48 51 51 49 47 35 2f 25 19 16 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0f 20 31 41 4d 50 47 41 3b 45 3d 46 43 49 42 4e 44 4e 53 4c 4c 4c 46 43 49 44 50 4f 4d 3e 43 4d 51 4b 48 53 50 51 4a 47 48 4e 43 42 46 45 47 3e 48 40 52 45 3f 3d 4b 3e 46 43 40 4a 50 52 48 51 40 42 44 41 3e 42 45 4c 50 51 50 44 47 3e 44 3d 3a 41 40 38 37 42 41 37 3f 41 48 43 3b 3b 3e 43 3b 41 3e 3f 3e 36 3d 3e 41 34 32 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 17 54 5f 74 65 65 6a 71 79 75 74 6f 68 67 6d 60 6a 64 5c 64 62 5f 5c 5b 59 5c 61 57 5c 55 59 58 5e 60 5e 60 62 55 5c 5e 5e 60 5a 5d 57 54 58 56 52 51 4a 48 4d 50 52 4b 49 54 51 53 54 51 53 57 4f 51 4f 4f 44 46 4a 51 50 4f 48 4f 51 52 50 4a 45 49 4e 44 44 41 33 32 25 11 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 23 2c 32 55 4f 46 44 3f 40 41 49 46 46 4a 48 49 47 4a 4a 48 49 4b 4c 45 48 4a 4d 51 4b 53 53 44 4e 4a 50 59 4f 4a 48 47 4b 49 44 4b 4c 41 49 37 4f 44 43 47 40 3e 46 3d 38 47 41 46 48 4f 4a 45 47 43 44 42 45 47 48 48 49 4a 4b 4b 46 40 3e 3c 3e 3e 35 3f 36 3d 3c 3d 34 3a 37 34 41 41 3f 40 43 42 3d 3c 3f 3f 36 37 3a 32 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 20 55 6d 6c 76 6f 70 77 72 70 74 6e 6c 6a 6b 66 67 60 68 5f 59 5e 61 5f 5d 5e 5d 62 5e 64 66 5e 5f 5a 5c 5a 58 59 61 5e 61 63 66 62 65 57 5d 5f 56 51 4d 4a 45 50 50 48 56 55 51 4c 4d 56 50 55 53 53 51 4e 55 4b 4c 4d 4a 46 4c 5f 4d 4e 4e 56 52 4a 4e 49 48 3c 32 25 1b 0a 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 16 1b 2b 36 44 50 46 4b 3f 46 42 44 4d 4b 4a 4a 3d 46 4a 56 49 52 4f 4c 47 46 50 4c 4a 4b 4e 4c 4f 49 43 4d
 51 42 45 44 46 48 3d 40 47 44 49 4a 42 3f 44 3b 41 41 3c 48 3f 3d 45 38 46 44 3f 45 40 4b 4d 46 47 43 4a 49 48 50 4c 4b 48 41 3e 3f 3f 36 3e 39 3c 3e 3d 3a 3d 40 37 40 38 45 44 46 3b 42 3c 3c 45 44 40 34 3b 3b 35 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 1a 52 69 7c 6e 75 63 68 6d 6a 69 6b 70 6a 66 66 66 61 5f 63 64 5c 5f 5c 5d 63 5e 5a 56 5a 60 5d 61 60 5b 60 67 62 66 5c 63 5f 65 5d 5d 5b 4e 5a 51 59 4b 4d 50 4a 54 4c 55 58 55 50 50 50 54 59 55 51 53 55 4b 55 4e 50 45 47 54 54 58 54 52 56 49 4c 45 40 40 44 31 21 17 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 15 21 33 41 46 43 44 41 42 48 47 49 4f 4f 4f 4d 4a 48 47 42 4d 4a 47 47 40 3f 51 42 45 4a 45 45 47 4a 4a 47 4b 44 43 3c 40 3d 43 3c 3e 36 45 41 39 39 3f 39 3f 3a 41 36 39 41 49 45 42 45 44 3f 3a 44 42 41 47 3e 3c 45 43 41 42 42 3e 3e 3e 39 45 41 3c 3d 36 3b 3c 3c 37 3c 36 39 3b 42 46 42 46 3a 41 3e 43 43 3d 3d 33 3c 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 15 4a 66 6f 78 77 70 6a 71 65 6e 6e 69 66 61 63 5f 5d 65 5d 5e 58 58 61 5b 61 5f 59 59 64 58 63 5d 5a 61 5e 62 60 5e 62 65 63 61 51 50 5c 4f 50 4a 51 4e 47 55 54 48 53 4e 51 53 55 51 4e 56 58 59 56 52 47 45 50 48 4e 4d 4d 4d 4e 45 52 4d 54 54 4c 4f 46 43 42 2c 23 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 09 19 19 24 43 42 40 45 40 42 48 4d 4f 4c 43 4b 47 46 4a 47 4a 45 51 44 48 4c 4a 44 45 4f 4d 4b 4f 41 4d 4b 4a 47 45 43 40 43 3e 3f 43 3e 45 3a 3a 3c 42 3a 35 3b 3f 40 3b 3e 41 42 3d 3b 3f 3e 44 41 47 45 47 47 3c 3f 3e 44 4a 46 48 3b 40 3d 38 3f 3e 3d 34 36 3b 3d 33 44 3a 39 40 3a 3c 3a 48 3f 47 41 3c 3c 40 44 3b 43 35 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 4f 6b 6b 73 72 62 6c 6e 6b 5f 62 66 69 65 61 62 59 5e 63 5d 5e 53 64 5d 5d 5e 5f 5a 5f 62 60 61 5a 5e 61 68 64 57 6c 65 61 61 59 51 5f 53 4d 50 50 47 49 52 4a 49 50 4a 51 58 59 55 57 60 56 58 52 4a 4d 45 3f 51 54 4d 4d 50 55 52 51 50 4f 4e 4d 4f 42 45 30 2a 16 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 14 2a 33 4f 46 3f 49 49 45 44 4b 4a 4a 48 46 47 43 40 50 4b 4b 49 3e 42 49 45 50 4b 4d 4b 44 4d 51 50
 50 49 46 46 4c 44 40 45 45 45 3d 3b 40 43 40 4a 3f 3e 3a 3e 41 3c 38 3b 41 40 38 3e 3f 41 43 3c 41 3e 38 48 39 44 3d 45 47 42 40 41 40 3e 42 3a 44 3e 3b 3b 3f 3d 33 39 3f 3b 45 45 37 46 41 43 48 45 48 41 3d 3c 39 23 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 13 4d 67 73 72 71 63 69 68 65 6c 6a 62 69 6c 60 61 61 5e 5f 5a 5d 5f 67 53 69 59 67 5f 67 62 66 64 68 65 5d 64 67 63 61 61 5d 5b 5b 57 54 54 54 5a 4a 55 50 4a 53 4e 51 43 4b 5f 54 5a 56 62 60 57 4d 50 4a 4f 4b 46 4d 52 46 52 5a 49 53 56 50 51 44 49 46 42 2f 23 12 10 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 10 20 33 3e 3b 40 44 44 43 45 4c 4b 47 42 4a 4c 46 3e 40 47 4b 49 45 42 48 4a 45 47 4a 3d 43 41 41 48 46 4e 44 45 3e 3b 3b 45 47 37 44 3d 3a 44 3d 42 41 3d 44 40 33 44 3e 3d 35 39 3d 38 36 36 3a 39 43 40 43 42 3a 44 40 3e 4a 41 3f 45 48 42 42 42 42 39 44 3a 38 3d 40 3c 41 3a 40 3f 47 3b 44 48 48 3d 38 44 45 42 3d 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 4a 68 6a 73 76 65 6b 6a 6b 62 6b 6a 6d 62 5f 61 59 62 65 64 68 5a 60 5c 65 64 62 63 5e 61 62 66 64 5a 63 60 62 64 60 5e 60 69 59 59 5b 4f 51 51 49 45 4c 54 56 4f 4a 4a 4b 54 59 57 64 60 60 58 4f 4f 49 4f 4a 47 4a 4e 54 52 48 53 4f 47 53 53 46 4a 40 3a 2a 1b 11 08 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 12 21 30 37 48 42 40 3e 48 47 4d 50 44 49 41 4c 45 42 45 50 46 49 47 46 4a 46 41 43 47 46 43 46 45 49 45 4c 44 3b 40 42 47 41 39 44 31 3d 3c 3b 48 42 41 3d 3f 3c 33 38 3c 38 36 39 3b 3a 35 37 3e 45 4a 47 3e 3e 3b 3a 45 42 40 44 42 44 45 42 38 47 49 3b 42 3e 3e 35 36 3c 40 42 44 49 45 4d 3b 46 3d 45 41 41 41 45 47 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 12 44 65 69 6e 64 62 6f 6f 66 64 5f 69 64 5f 65 59 5f 5d 60 65 64 61 60 60 6e 5e 65 60 69 62 62 60 71 68 64 6b 5b 64 63 62 66 61 5e 56 58 57 50 52 4f 48 4e 47 4e 4a 4f 52 50 54 54 61 67 62 63 57 50 4f 42 4b 42 4a 4a 57 4d 4f 50 54 4b 57 56 4e 4b 39 3a 2d 24 17 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 13 28 37 47 41 46 45 44 47 4d 4b 41 47 4e 4a 46 4b 42 40 45 44 46 43 47 41 44 48 46 41 46 44 48 47
 4b 3f 42 3f 48 3d 36 41 3a 3d 42 3f 3c 45 3c 33 3e 3c 3d 3e 3d 38 3e 31 3e 3b 41 35 39 3b 37 44 3a 3b 3a 3f 3a 40 40 3b 3d 3b 42 41 44 42 48 47 49 47 46 3c 44 39 3f 41 3d 42 46 40 3f 44 44 45 3e 44 3c 47 40 50 3f 25 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 3a 64 73 6b 65 63 69 6a 63 67 64 68 66 65 63 67 66 68 65 62 68 66 60 64 65 68 6b 68 63 6a 69 68 69 6c 60 5d 67 62 66 62 5a 5a 58 55 54 55 56 55 4e 47 4c 50 4f 51 57 4d 51 5f 63 68 5f 60 62 59 4f 4e 46 4a 48 4e 5f 4e 49 4b 52 52 59 49 54 48 3f 44 34 31 19 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 1f 2f 41 42 3b 4c 47 43 4f 4b 48 45 41 4d 42 43 45 4c 46 44 42 42 47 44 40 44 3f 44 3a 3f 3e 4b 40 3f 41 3c 3f 41 39 45 3d 40 41 40 3a 2f 41 39 37 37 36 3d 3c 30 38 37 35 39 33 36 2f 3a 46 43 44 40 37 38 4c 41 43 39 3b 42 49 46 41 3c 44 4a 52 4e 48 45 40 39 3e 40 3e 3d 40 3c 3e 41 44 46 47 38 40 3f 3f 3a 42 29 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 09 44 5f 6b 6b 65 64 6d 6f 64 6a 60 61 69 62 61 66 5d 5b 69 64 65 5a 6d 5e 6a 62 64 63 62 5d 66 6b 66 65 65 64 61 5a 63 55 53 62 51 4e 56 50 50 4e 50 53 48 4e 47 4f 51 54 50 55 62 66 67 61 5d 55 50 4b 4d 49 48 4d 42 4f 49 4e 56 52 4d 4e 4a 50 40 3b 36 29 1d 0d 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 1f 2d 46 43 42 4c 3e 4a 47 47 44 41 46 41 48 4c 3b 43 41 40 48 3c 43 40 3b 41 43 3f 45 45 47 42 47 3f 38 3e 36 3a 3e 38 42 39 38 3d 35 3a 3b 3c 41 3d 3d 30 3d 30 35 3b 36 36 36 32 3d 37 3f 3d 33 43 43 40 3e 43 36 36 39 3d 41 49 38 41 43 49 45 46 45 3d 3d 3a 44 3e 34 40 41 3f 44 3f 42 42 40 4a 3d 3a 42 42 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3a 5f 67 65 65 69 6f 6b 66 5f 6b 62 64 5c 61 62 60 62 65 69 65 67 68 63 62 68 66 62 66 5d 6f 65 65 64 5f 5f 5f 5e 52 55 59 58 57 4d 4f 4d 51 4d 48 55 44 4e 54 46 50 4b 54 56 5f 61 63 61 61 51 4b 48 4c 49 4c 48 48 4b 4e 51 55 52 54 43 47 3c 3b 3b 2d 28 10 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1d 2c 41 43 44 49 45 48 42 49 47 44 47 4d 47 3d 45 45 3c 43 45 44 4c 41 44 44 44 3a 40 41 41
 3b 42 41 47 46 42 3e 3e 3d 3d 39 3d 41 35 38 39 3e 40 3a 3d 36 3a 41 34 41 36 3b 38 32 36 39 40 40 34 3a 40 40 4a 3e 3e 45 3f 3e 47 45 3b 3e 42 48 45 47 43 42 3d 48 40 3d 3e 44 43 42 3d 3f 3c 49 47 45 49 41 44 3e 2c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 3a 5f 60 68 67 6a 6d 6d 5c 69 60 6b 68 5f 65 68 63 67 69 61 6b 67 65 6a 64 67 66 67 68 61 61 62 64 62 64 62 62 5b 51 5c 50 54 5a 54 50 4d 55 4f 54 4d 50 4f 46 4d 51 49 57 57 5b 65 65 66 5b 52 52 4c 4c 4a 4a 4b 52 46 53 55 4f 56 50 47 4b 48 45 3c 2b 26 13 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 17 28 34 3e 44 49 46 4a 49 44 3f 41 49 43 3a 41 3f 42 45 40 3d 3c 3f 3f 43 40 46 3e 45 43 40 40 43 34 41 3c 3f 39 3c 3b 36 32 32 34 3e 37 3c 38 36 38 37 39 36 38 37 38 39 42 3a 2f 2d 3a 3d 33 38 3e 3a 40 3f 49 40 45 49 45 47 40 42 45 42 45 3f 3f 43 42 45 40 3d 3a 42 46 41 3b 48 40 44 42 43 3b 42 3e 3f 38 2b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 2d 5d 60 6c 6e 67 6f 6f 69 67 61 5d 5c 5b 65 5b 5f 69 66 66 62 60 6d 63 6a 67 60 66 61 5f 62 65 5e 5d 5e 5d 5f 5d 5d 53 53 56 53 4d 4d 50 4e 51 51 48 51 43 46 47 4e 48 58 51 5d 60 5e 5c 55 55 52 4b 4a 4a 4f 4e 4c 52 57 50 52 55 55 4b 44 44 3b 3e 2c 16 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 23 2d 3b 3c 3f 44 4b 4b 48 4a 40 40 4b 3e 3a 44 40 42 3a 3e 37 37 44 43 37 45 3d 3f 3e 43 40 3c 36 3b 3d 3d 2e 3d 35 4a 32 34 3c 44 38 34 32 37 34 3a 3b 32 36 35 39 3a 41 28 37 33 3d 40 34 34 36 44 38 39 3d 42 4a 48 49 4f 46 49 39 45 46 3e 40 45 3b 46 3d 3f 42 3f 40 41 41 3a 42 43 42 43 3c 3f 3b 3a 41 2b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 34 57 61 6c 67 57 6c 62 5d 64 61 5d 5e 51 58 5c 5e 64 60 65 69 65 61 5d 67 61 67 6c 66 69 64 69 60 6d 5c 61 61 5b 5c 54 53 52 51 55 52 42 44 48 43 4d 42 4e 4a 49 4d 52 52 4f 52 51 5b 54 52 50 49 4e 4b 4c 4e 46 4a 4b 49 52 52 50 55 42 46 3e 3a 33 1f 19 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 11 12 24 33 43 43 47 4b 4b 4a 45 42 4c 4a 44 3e 43 3c 44 44 3e 41 3f 3e 3e 3d 43 35 36 37 43
 3b 42 3e 3e 3c 3e 3a 47 38 36 40 3c 34 38 39 3e 3a 3c 32 43 3a 3d 36 2e 38 36 35 3a 38 37 3d 3e 3d 39 31 3c 32 3b 42 40 42 3f 48 49 43 46 42 45 41 43 47 4a 42 4d 3f 3b 3c 37 44 3e 41 36 3f 3e 3e 3d 47 41 4a 41 3a 30 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 32 61 6e 63 62 5e 66 65 5c 5b 5b 5b 5e 55 56 58 5d 62 5f 59 65 62 6d 60 65 64 62 63 69 65 64 66 64 62 5e 5d 5d 57 55 55 58 50 4f 51 54 4c 4d 51 47 47 3d 4c 46 41 44 45 52 55 53 5c 58 52 51 50 49 4a 50 50 52 49 4c 4d 51 4a 4f 51 4d 47 49 37 35 2f 17 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 1c 32 3a 3a 47 52 4c 46 47 44 41 3f 46 47 3c 44 45 3b 3b 37 42 3e 46 3b 3d 39 37 40 3b 3c 44 3f 3c 3b 33 34 41 38 3c 37 3c 37 39 3c 35 3d 36 33 35 32 39 38 38 39 33 32 3f 3c 3b 3e 37 3d 3e 3b 3f 3e 34 38 3d 45 40 43 47 3b 46 44 41 49 41 41 44 38 44 42 43 32 3c 42 3c 40 3b 3a 3d 36 41 40 3e 3c 3e 40 34 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2c 5b 5f 5f 63 5d 64 5f 58 55 5d 51 5a 57 5a 57 5a 63 5f 5d 64 64 61 60 66 67 6b 6a 65 61 66 64 5f 5a 5d 5d 5d 58 55 52 50 50 51 4f 4e 49 46 51 4d 4a 46 4b 43 44 4a 48 4a 56 50 50 4e 50 50 47 4e 50 4a 4f 4a 4f 4c 4f 50 4e 58 51 52 3f 3c 3d 34 1f 19 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0c 0e 24 38 3b 4b 46 40 47 43 3f 48 3d 44 34 36 40 38 47 3f 3d 34 39 36 36 3b 35 39 36 3e 33 43 36 3f 34 30 33 34 34 35 3b 31 36 32 2b 40 33 37 36 3c 30 37 35 39 38 36 2d 3e 32 32 36 3b 37 37 41 3d 45 33 38 40 3b 3d 39 36 38 3c 43 3e 47 3c 40 3e 3c 42 3d 38 39 38 40 3e 3a 33 39 3f 3e 40 3d 3d 3b 3b 44 27 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 52 62 58 68 54 5c 54 51 54 51 52 55 55 50 56 52 56 59 56 64 60 61 64 62 6b 60 63 63 61 60 61 58 5a 57 59 63 5a 53 57 5b 4a 4c 51 52 4a 4b 4b 46 46 44 4d 47 45 49 48 4f 4d 50 56 51 49 4b 59 4c 50 4e 4d 4c 41 4a 49 48 51 4c 41 4e 38 39 3c 2d 1d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 09 10 1e 33 37 44 4a 41 47 42 40 46 41 48 35 3e 3c 3b 41 42 37 35 42 38 34 39 36 43 3d 43
 31 38 37 3c 3e 3a 32 3b 3e 36 3e 38 37 38 3a 39 38 32 32 35 39 35 33 3f 3d 35 36 34 39 3a 3d 33 3c 3d 39 41 34 39 3e 3e 42 38 39 34 3f 3d 3c 40 46 41 42 3f 3c 49 47 3c 3c 41 3c 3b 3a 41 45 41 36 3a 3e 3e 41 3d 3e 34 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 55 61 60 5a 56 5a 5b 55 54 50 57 54 58 54 4e 5b 51 58 59 5a 5a 5f 5f 6a 60 63 5e 5b 66 60 56 5a 59 53 59 5d 57 4c 54 54 5b 55 51 4c 4a 48 52 52 48 44 3e 48 4a 4a 4a 51 4d 4a 4e 46 44 4f 4f 44 47 50 41 4e 4e 54 4f 4f 4e 51 45 4b 40 3b 39 25 19 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 14 2b 3b 3d 45 45 43 44 46 42 34 38 3e 41 3d 3d 33 3b 39 41 36 44 3a 3f 3e 3d 3d 34 3b 3c 36 3a 3f 36 32 38 33 32 34 39 38 2f 36 39 37 32 3c 30 31 37 39 38 39 38 37 36 36 32 3d 3e 46 41 3a 37 3c 3e 43 3c 3e 38 3e 3e 3c 3f 3d 3d 44 3b 41 49 41 41 44 43 3d 3b 3e 45 3b 3e 3f 39 40 38 38 3a 3d 37 37 37 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 4c 5c 5c 5a 57 55 5c 4b 4f 51 49 5a 52 4f 4d 58 55 57 56 58 5b 5f 5a 5e 5f 64 5e 59 62 5f 59 5d 55 5a 59 5f 55 58 4c 57 54 48 4b 50 4b 40 44 47 42 41 4e 4e 4d 4b 4b 52 48 47 50 47 3d 3e 4e 49 4c 45 4a 4e 41 4f 4a 49 4e 55 4c 4f 3b 3b 25 18 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 1b 2d 3e 3f 3e 42 47 47 3b 45 42 42 38 42 3e 36 37 3e 42 39 37 40 43 37 37 37 32 38 35 37 3b 32 33 3d 33 3d 39 35 35 38 36 32 38 38 38 36 33 2a 3b 3c 38 42 3f 35 36 39 3c 41 48 48 35 3a 3f 40 33 38 38 34 3c 3e 3b 3d 3d 32 41 45 42 44 44 45 44 43 49 3a 3f 36 39 3b 3c 3a 3d 39 3e 3d 3c 3f 3f 3a 34 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 52 58 59 4f 50 52 50 4e 4e 4a 52 47 51 52 50 4f 53 53 57 52 5e 56 5c 64 63 66 5d 5f 5c 50 5b 58 4f 54 55 51 4c 52 4d 4d 4c 4d 4b 48 4a 4d 48 3d 49 4b 4b 42 4a 51 46 59 50 4b 48 4c 49 47 48 44 4b 45 4a 48 44 4c 4d 4f 4a 48 45 43 42 2f 2b 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 21 35 40 3a 3f 44 3e 44 3f 40 42 3a 39 31 38 35 38 3f 41 3b 3b 3d 43 36 3c 3d
 35 3b 40 2e 38 32 38 3b 39 31 3a 3a 3b 35 32 36 33 34 36 37 30 33 38 32 3a 34 35 34 38 37 46 34 22 2f 47 43 3b 35 32 38 39 3e 3b 35 31 35 35 3b 45 3e 4a 44 3c 40 45 3f 45 3a 37 3b 3e 43 35 3a 42 3b 40 3e 39 43 33 39 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1b 4f 51 5d 58 50 4b 51 49 48 4b 45 4e 49 4f 55 51 46 58 5d 52 55 5d 5b 5d 56 5e 63 56 56 59 4f 50 58 50 5a 52 4b 45 45 4f 52 46 45 50 45 47 4b 4a 4c 4e 4b 49 48 46 4a 53 44 47 48 49 4d 44 46 44 42 42 4e 4a 4c 4c 4f 52 49 3e 47 41 36 2e 21 10 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 18 28 39 44 41 46 3d 3f 42 40 3f 41 38 3e 3b 3d 3d 3b 3c 3b 37 39 3d 37 3a 35 35 36 37 3a 38 37 37 38 35 37 3e 35 40 35 2b 35 37 2d 37 31 39 37 35 2d 3c 32 32 3e 35 3f 3b 3e 46 4c 4d 40 35 3a 39 39 3d 37 36 3b 35 35 3b 35 35 35 39 43 49 4d 4b 4d 41 41 3e 3d 33 3a 3a 3c 3c 3d 3f 42 37 3a 3e 31 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 45 55 51 50 46 4e 4d 3d 49 47 43 4c 49 52 52 49 4e 4b 4d 4a 50 57 5e 57 5b 5f 5c 52 52 5b 5e 57 4c 52 56 52 4f 4f 55 53 4c 4b 4c 44 3e 4d 4c 49 43 48 40 52 42 42 49 51 3e 46 47 47 4b 46 4b 47 41 45 42 53 41 4c 3c 4e 45 47 4d 42 34 29 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 10 1f 39 42 3f 48 45 39 40 3e 41 3e 41 3d 3c 36 3e 37 3c 2f 3a 3a 36 3b 34 36 34 31 34 32 36 3f 32 35 38 33 30 2f 37 3d 31 33 37 34 35 2e 35 38 33 37 38 3c 34 3c 38 35 49 47 49 47 47 47 33 36 39 30 3c 3e 3a 3b 32 3b 36 3a 40 3b 3a 39 43 47 44 4a 3c 3b 39 34 3b 40 31 3d 3f 3c 42 39 32 3e 34 31 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 47 49 50 55 43 49 42 45 41 46 42 4c 41 4d 47 48 4a 4d 52 4f 4f 59 4c 59 59 5a 57 54 4a 53 50 53 53 4f 55 4b 4e 4b 49 45 4c 50 40 47 3b 47 4d 4c 47 47 44 45 3f 3e 3e 48 3c 42 3f 45 3f 4d 3d 4a 3c 46 4b 44 47 4a 45 46 44 48 45 3f 28 1f 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 06 06 18 2c 34 45 43 40 3b 43 3b 41 38 3e 35 32 3a 3d 40 3a 3e 38 35 38 30 3c 3b
 31 35 41 31 3b 33 37 35 34 37 35 34 2e 3a 38 38 31 31 32 3d 2c 31 2b 31 36 3d 33 2f 3b 34 3f 47 51 4e 4a 46 38 34 33 37 31 3a 41 41 38 37 2f 35 3a 3f 3d 42 40 4a 44 46 44 3a 3b 42 3f 3b 3f 38 3a 36 32 3e 3f 35 4a 31 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 3f 50 4d 4b 41 49 45 48 43 43 3e 41 49 4a 4a 46 4b 50 51 4b 4c 4f 4b 51 53 51 4d 54 55 58 56 51 51 53 51 4b 47 49 4b 47 3e 4a 4b 48 44 49 43 44 47 4c 3f 42 4b 46 4c 41 44 47 45 48 3f 3d 47 48 45 46 4c 4b 40 4c 47 46 47 49 44 3e 2c 13 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0c 22 2d 3e 3d 41 45 3b 39 3e 3a 39 38 34 3f 38 40 33 3b 39 37 3b 34 3b 3a 38 32 3a 35 34 33 36 3e 38 34 34 3d 33 35 34 39 34 39 30 37 35 33 34 38 37 2b 36 3a 37 3b 40 44 4e 4d 54 44 36 3f 38 43 45 36 3d 3a 37 35 40 35 30 30 3e 43 47 4a 49 44 42 3a 39 3e 32 37 3d 3c 3a 40 36 40 3f 3d 3c 3b 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 41 4a 41 49 42 4a 3d 4b 40 42 41 54 44 41 49 4a 42 49 48 4a 4f 55 53 57 4d 56 59 53 57 52 51 51 51 51 4b 4a 4a 41 48 45 42 4c 44 43 45 4b 3e 47 49 42 4c 41 3f 45 42 44 3b 44 44 45 42 45 49 44 4c 4b 52 4e 44 4d 41 4a 43 47 3b 2f 21 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 16 20 27 3b 35 3f 45 3e 41 3a 41 36 3f 36 3b 36 38 36 3b 3c 38 39 33 3e 3c 2f 31 36 34 36 39 38 2e 36 3b 36 34 35 31 31 36 2e 3b 35 34 35 36 34 33 39 3c 44 31 2c 39 3e 48 47 41 3c 36 35 38 39 46 34 32 37 38 3f 3d 3d 36 3c 41 3c 3a 3b 3e 37 3a 3a 3f 44 3c 3d 34 3e 3c 3c 31 40 42 3f 45 39 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 39 43 3d 44 41 49 3d 3e 3c 3b 3f 43 42 42 3e 4b 41 45 49 4f 4d 50 4d 4c 46 52 49 54 5a 54 58 54 48 54 4c 45 4b 49 4a 49 47 46 40 48 4a 45 4b 45 3b 3d 3f 44 38 3c 39 44 3f 3e 41 3f 3e 44 40 45 44 46 45 51 47 49 4a 43 4b 43 35 30 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0e 16 2d 40 3b 44 3a 3c 3d 3c 3d 3e 3b 31 3d 37 44 33 38 39 3a 34 32 30
 33 35 39 2b 38 32 32 35 36 32 36 35 2f 33 31 34 43 35 30 39 33 33 3b 36 41 30 31 34 37 34 37 3b 48 3b 3c 3f 3f 34 38 3f 3d 34 3f 34 33 3d 33 3f 3a 36 3e 44 47 3e 40 3d 42 36 35 39 3b 3d 34 3d 3e 43 40 3b 37 31 38 33 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2c 41 41 4a 39 47 48 44 3a 3e 41 42 4b 42 47 44 42 50 44 4a 4a 49 4a 4e 4f 4e 53 4b 56 4e 47 4c 4b 51 55 4d 3e 46 52 43 45 44 3a 47 45 3b 47 3a 43 3f 40 45 3a 46 41 43 41 43 49 42 3f 41 3f 42 47 4d 3e 47 44 45 44 41 3c 3a 3d 27 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0b 1a 1d 2e 3b 49 3d 41 3c 47 35 37 3e 34 3c 3c 43 41 3f 3d 39 38 36 30 3a 3b 35 3b 36 37 35 36 31 33 38 31 32 39 34 35 32 30 39 3d 35 3e 41 3a 39 35 39 35 3c 32 39 3a 3e 39 39 3c 3b 39 39 3e 3c 35 3b 42 3d 3d 3d 45 3e 44 3d 43 3c 4d 3f 3b 38 3d 3d 40 41 3f 3c 40 39 35 3c 41 46 3c 3d 37 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 38 46 40 44 3c 3b 3b 3c 41 42 44 3e 41 4a 42 48 41 50 4d 56 44 45 4f 4e 4a 53 53 57 52 4b 53 50 4f 51 4c 52 44 4e 42 49 4c 46 49 43 4b 42 3e 40 45 3f 45 3e 3e 46 37 47 42 3e 4f 44 38 3f 40 50 50 4e 49 45 3e 49 44 44 43 35 2b 1e 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 13 2c 39 3e 3e 37 45 41 3c 3e 37 3e 3e 3f 40 3a 41 3b 39 38 3e 31 30 41 36 39 39 38 34 36 3b 35 34 3b 3b 39 32 3a 33 2e 31 34 30 38 36 3c 37 34 3d 37 36 38 34 3b 43 42 42 42 45 37 36 36 36 35 42 39 3e 3a 3e 3d 3b 42 43 43 3e 44 36 3e 3a 39 3a 3d 3e 3c 3e 40 3f 3d 3e 38 3b 3e 47 3f 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 2d 3c 40 48 3d 3e 3f 3e 44 39 40 41 3f 48 46 4b 41 4e 49 4e 4c 42 4d 4a 4a 4b 4c 55 49 58 4d 54 4f 51 50 49 49 47 3b 44 43 46 43 44 3c 36 47 41 43 46 41 3c 41 42 42 42 42 3a 38 43 41 4f 41 49 48 48 42 4f 42 3d 3e 41 47 2f 25 1a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 1f 2b 38 3f 41 37 44 37 3c 38 40 3d 39 40 39 3e 3f 3d 39 31 37
 40 39 35 36 32 3b 35 36 33 30 37 3a 2c 2f 35 3d 31 36 35 3a 30 39 36 38 3a 35 36 3b 39 34 36 39 39 3e 3b 3d 37 34 39 39 35 34 3a 3a 38 38 3a 40 41 39 40 40 3b 3c 44 39 3a 3b 40 42 3e 44 35 3e 37 40 42 3b 37 3e 36 38 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 26 3c 3e 41 3c 37 3a 3b 39 44 38 49 37 41 43 43 46 42 45 43 43 4d 47 45 4a 4f 48 45 46 48 53 47 48 47 47 41 49 3f 3f 44 3e 3e 3b 3c 3e 39 3e 3f 3e 3a 36 38 37 43 40 42 49 43 43 46 3b 3b 39 40 45 4a 45 45 45 42 3d 45 38 23 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 14 2c 35 3e 41 40 42 3a 3d 41 40 3f 40 39 37 3e 3d 39 38 39 43 37 34 36 31 30 38 34 34 35 3b 37 2e 2c 38 3a 39 39 2f 35 40 35 30 3d 36 36 3b 39 3d 37 38 35 43 3e 3e 38 35 3a 39 37 3d 3b 35 3b 37 36 40 32 41 3f 39 38 41 40 41 42 3a 34 3d 36 42 3e 41 42 3e 40 43 3e 42 3d 41 3d 36 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 23 39 40 45 39 35 39 37 3c 3e 3d 3e 3a 43 3b 43 45 45 4b 3f 45 4c 4b 51 4b 5b 44 49 4b 4d 50 4f 47 42 47 3f 40 43 45 45 44 46 36 42 3c 40 45 43 3f 46 43 48 40 3e 3e 47 47 39 41 40 3d 46 3e 45 4a 4b 44 4f 44 41 45 34 21 1f 0d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 16 2f 35 42 3b 38 43 41 3a 3a 3f 43 38 3e 3e 3b 3b 34 35 40 41 42 31 34 39 39 34 34 36 3a 32 3a 3a 39 3a 3a 3b 37 37 3b 32 38 3b 34 3b 39 36 3e 3b 43 41 40 3e 3f 40 37 38 34 38 3f 3c 33 3b 3f 3b 42 33 40 3d 3a 39 3e 31 44 39 41 39 40 3f 3f 45 3c 39 35 3b 3a 3d 3e 3f 41 3a 3e 25 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 25 37 3c 40 39 37 3e 40 37 3a 35 40 3b 42 45 43 43 42 47 4c 45 47 4f 4b 48 54 4b 4d 48 51 48 4f 40 4b 49 40 41 41 3d 46 40 46 47 42 40 3e 46 44 39 41 42 43 42 41 3f 3b 46 42 41 3f 3c 4b 47 40 49 46 3e 49 43 45 3c 37 22 0f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 16 22 37 3b 3c 3f 3b 40 33 37 38 3e 3a 38 3a 3f 3e 3a 3b 37
 31 3b 31 34 31 32 35 38 37 3e 37 35 38 36 36 34 32 31 3e 3e 34 38 3a 33 32 35 2e 38 33 3a 36 3a 3a 39 37 3b 36 3e 3a 40 38 35 3a 3b 36 3a 38 3c 3a 34 3a 36 3b 39 36 38 3c 3b 44 3c 40 44 43 39 3e 36 46 36 3a 3d 3e 33 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 27 32 30 3f 32 39 36 3e 3b 37 3d 3f 45 44 3e 46 47 44 43 44 41 48 47 45 4d 4c 40 51 48 47 40 47 43 44 45 43 3c 3e 47 3e 41 3f 43 42 3e 3e 38 4d 3d 3a 40 44 3b 3e 3f 45 48 43 40 3a 3e 3b 45 44 42 44 42 44 39 3e 36 29 15 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 19 34 34 3c 41 41 3f 43 38 3a 40 3e 3c 42 42 38 36 37 30 38 39 30 32 30 32 38 30 39 31 34 33 32 35 36 32 34 33 3c 38 3b 35 38 35 36 34 3d 38 36 39 3e 35 3e 3e 3e 41 31 3a 3c 3d 3c 3a 40 3c 34 3a 43 3d 46 37 3e 3f 3e 39 37 32 3a 46 43 43 45 3f 3e 3f 38 35 42 3d 42 45 3f 3a 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 39 41 3c 34 36 45 3c 3e 41 42 40 43 3d 40 49 41 42 45 44 42 46 3e 44 42 44 4b 3e 48 43 4d 4a 3b 3f 3d 47 3b 3b 45 40 41 3d 45 45 4a 45 3e 40 40 3d 3c 40 3d 4a 41 47 3f 39 43 3d 3b 44 41 41 4a 4d 45 46 3b 39 34 1e 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 15 25 45 44 47 45 3a 37 3e 3b 44 3a 39 45 3b 42 42 36 38 35 3c 30 3c 35 34 34 36 39 42 2f 34 33 35 3b 3d 3a 36 39 33 33 3c 35 36 39 35 41 37 37 31 37 43 39 3c 44 38 40 39 37 37 39 44 39 42 37 39 3e 39 3d 43 3a 3d 3e 45 3d 3d 3a 35 43 3b 3c 42 3c 44 3f 40 3f 3d 3d 42 3b 3b 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 20 3e 3e 39 36 3d 38 3f 3e 42 3e 39 34 45 3c 46 44 4a 48 4b 43 49 43 47 40 4c 45 44 48 44 45 3e 44 47 3c 44 43 44 4c 3f 3b 42 3d 3f 3e 3b 3f 41 3e 3b 38 41 36 3f 44 3e 3b 3a 41 3f 43 4a 44 43 41 53 4a 47 3d 34 21 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1c 21 2b 3a 3f 45 39 3e 36 3a 41 3b 3e 37 3d 35 32 39 39
 3f 34 3c 36 3a 3b 32 34 32 2d 37 3c 35 33 32 34 42 30 3f 38 3b 31 35 3c 36 3b 3c 35 34 33 35 35 3c 34 3a 3c 37 36 38 3a 3c 45 43 3d 3b 36 38 3a 38 34 3d 3b 3a 44 39 38 36 39 34 46 41 3d 37 3a 3d 41 40 40 44 3d 36 3c 2d 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 35 3e 41 42 3f 3b 42 40 3e 36 43 41 39 43 41 45 48 3f 42 3d 47 49 42 49 49 43 3e 40 44 41 47 39 34 42 43 41 3b 43 44 45 37 41 3e 3a 40 40 3c 3c 45 39 3d 3d 3d 35 43 3a 45 42 3d 45 47 3e 43 39 43 45 3f 34 2e 1f 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 16 20 3b 4e 46 43 38 3f 40 41 3a 3e 43 3d 44 41 37 37 3b 35 3d 37 33 36 37 32 31 3c 36 2e 38 3b 37 38 39 39 3d 38 32 3e 3c 3d 3c 33 3d 3f 33 39 40 39 3e 3a 3e 3e 3d 39 45 44 3a 3d 41 39 40 41 3c 43 3c 41 41 3c 40 45 3a 40 41 41 3d 45 40 40 44 3c 42 40 3f 3a 39 3f 48 3a 28 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 35 38 35 33 41 3e 39 3d 3a 3e 42 45 49 3d 45 47 41 45 43 44 4c 42 48 46 4a 44 42 44 4b 45 3f 38 43 3e 3c 46 3e 4b 45 44 45 38 3d 41 3a 3e 43 3e 3e 3f 3a 3f 47 3f 46 3d 38 4a 48 46 40 3f 41 51 46 41 39 32 23 12 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 13 29 3d 3d 3d 38 3b 3a 39 41 42 3a 3b 3b 3d 3c 3a 3c 3c 37 3b 34 3a 33 36 30 39 39 34 37 3c 33 41 34 32 36 44 31 31 44 3a 3d 47 34 43 3b 38 33 39 43 38 45 3f 38 3a 39 3f 41 3e 40 3d 38 3b 3b 45 3c 40 43 37 40 44 3e 39 3f 3e 40 47 3d 4c 44 3c 3b 39 3c 35 39 34 42 38 2b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 37 36 3a 38 3a 43 3d 3e 3b 3c 3d 3d 41 44 47 44 42 3f 45 3d 49 43 47 45 45 45 42 4b 4b 45 48 3e 3c 45 41 39 35 40 3e 3c 40 3c 37 48 41 41 41 3c 36 3f 41 30 48 3f 41 45 3b 3f 46 40 41 44 45 48 44 41 35 2a 13 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 26 28 43 42 43 3b 35 3e 38 3b 36 33 34 3a 3e 39
 3f 33 35 34 3b 3b 35 2f 35 35 36 36 35 39 3d 3b 38 37 36 39 2f 42 38 3a 36 3a 3d 38 39 37 3f 3a 32 3a 3b 3b 44 3c 3b 40 3f 41 3d 44 3c 38 42 42 41 39 3c 3f 3a 3c 3d 3e 3d 39 3d 41 3f 43 3b 3c 3b 38 39 3d 41 3b 40 37 25 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 31 36 3d 37 37 45 38 39 42 37 3e 44 3e 49 43 41 44 43 45 36 3e 44 4a 3b 49 41 3d 42 3d 3e 40 3b 3a 3b 3f 3f 3a 3e 45 3b 46 42 3f 3a 42 44 41 44 39 3a 40 3a 3b 44 44 41 3c 44 3e 3c 47 44 41 43 3e 42 2d 19 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 15 2a 32 3f 38 3c 3b 3c 3b 3e 3d 3f 3d 39 34 39 3f 3f 3a 2f 32 35 35 35 35 34 37 30 38 36 3c 3c 37 39 31 3e 34 43 38 34 33 33 31 38 36 3a 32 3c 3b 36 3d 3a 40 42 42 44 41 34 47 38 43 45 40 40 40 3d 38 3d 3e 34 3c 3b 43 3f 41 41 3c 3d 3e 39 3a 36 48 45 3e 3a 3d 36 2c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 38 37 3d 2e 34 36 3d 3e 3b 3b 47 3f 40 39 40 43 43 3b 42 41 47 3f 44 3f 43 40 45 42 45 41 44 3b 38 44 3f 40 39 42 3d 3a 3e 3e 42 3b 38 3e 3d 43 39 3b 41 3c 37 3b 40 3f 3b 44 3f 3d 43 43 41 4b 44 33 23 15 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0e 17 27 35 38 3a 3d 3a 3d 3d 42 3c 39 3d 43 3d 3b 37 40 3c 35 32 36 36 38 36 35 39 3d 32 36 3b 40 37 3a 37 3c 39 3b 3a 35 3c 35 3e 37 37 3a 3b 41 38 39 42 44 3c 41 44 47 47 40 3d 46 3a 36 41 40 43 3a 3f 3f 3c 36 3a 43 3e 41 41 3b 43 3b 37 3c 3e 3b 39 38 3d 36 38 30 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 36 31 40 32 36 32 34 3c 42 39 42 3b 3a 44 45 4c 3e 48 48 3d 3e 3c 49 49 47 44 41 42 42 44 43 3b 39 45 40 38 3e 39 41 43 40 44 3d 38 42 39 47 3e 41 36 3b 39 3d 42 44 45 4a 3e 42 40 47 45 47 3a 38 2a 1b 0a 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 07 18 2c 2e 37 38 36 3a 46 40 3a 44 3a 39 41
 42 39 3d 3f 34 36 3a 34 3b 3c 3a 37 38 34 34 3b 41 3b 36 3f 3b 3e 35 32 41 38 3b 37 32 3c 39 39 3c 3d 37 3e 3b 43 40 46 4c 3a 38 37 36 39 37 40 36 42 3d 39 44 37 40 48 3f 42 3c 3e 45 42 3d 3b 3b 41 3f 40 40 33 3f 37 26 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 29 32 38 3c 39 40 3e 36 41 3b 44 37 3d 40 42 47 41 49 3f 43 48 40 42 42 4a 48 41 48 3e 3f 3d 38 35 33 38 41 43 3b 42 3e 3b 3e 3b 41 41 3e 42 38 41 3a 38 37 3e 37 42 3c 3a 40 3a 40 40 43 3c 36 2a 18 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 15 1b 25 2b 33 3b 40 3c 37 45 33 34 40 31 3e 3a 36 37 3a 30 39 39 33 39 34 3c 31 3c 3b 3f 35 3b 40 39 38 39 3e 38 3c 36 2f 38 33 38 38 3a 3b 36 3c 3d 3e 42 44 45 46 3c 45 3e 3c 45 39 3f 35 36 35 38 3d 3e 3c 3d 41 3a 42 43 3a 3b 3e 39 40 34 3b 34 38 37 36 34 21 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 2b 2f 31 35 35 3b 3c 39 39 41 3b 41 40 49 41 3e 41 3d 42 48 49 3e 3f 43 48 42 40 40 46 3b 36 3a 36 42 3b 3b 35 3e 41 3d 3d 45 43 3e 35 3a 37 34 3e 3f 3e 3e 3d 3a 45 3a 3f 3b 3d 3d 44 3c 36 2f 25 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 14 20 26 36 36 37 3f 3c 44 40 3f 39 3b 3b 41 3e 3d 3a 3b 3a 3a 37 3b 3d 3e 33 44 39 42 3d 36 43 40 34 3e 3b 3a 41 36 39 44 2f 39 3e 38 3e 3f 3d 3a 40 3d 4e 49 45 43 41 39 32 42 40 3b 42 3e 38 41 31 3c 3f 35 3a 42 45 3e 3c 45 40 3f 3f 41 41 41 3c 36 39 3a 2a 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 31 3a 3b 2f 39 3a 39 3f 38 4a 47 44 40 37 39 44 3b 45 45 3e 41 39 3f 47 4f 4d 40 3f 3b 3b 3b 3c 39 37 36 39 3b 46 42 46 3c 39 3c 3a 3d 40 3a 39 3c 3e 35 3e 39 3b 3e 3b 3a 3e 45 3e 42 3b 2e 24 1c 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 14 1f 29 2d 42 34 36 3f 38 31 37 43
 39 41 32 37 35 3b 31 3b 3a 36 39 38 3c 40 3e 35 37 3d 36 38 3e 3b 3f 3a 39 37 33 39 39 3b 3d 3c 33 3f 3e 40 3d 47 4c 46 48 3d 44 38 3b 3e 38 37 3c 39 39 3d 3a 3c 3c 37 3e 37 40 39 36 3e 3e 40 3f 3c 35 3f 3a 35 3c 36 2b 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 27 34 40 39 3d 39 3b 43 3d 42 38 40 3d 39 40 40 47 3b 3a 3c 42 41 4a 54 41 43 3e 45 3a 38 40 34 3d 3a 34 39 44 3c 45 3c 3b 3c 47 3b 39 3b 42 3b 3e 37 3f 39 32 3c 3a 45 3e 43 38 3c 3e 32 21 1e 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 19 1a 2a 3a 34 34 3a 35 41 39 33 3e 3d 3e 3c 37 3f 33 36 3b 36 36 36 39 3d 35 32 32 31 33 3d 3b 3b 3e 2d 39 37 38 37 36 36 35 3c 39 39 40 40 3e 47 52 4a 4c 4f 50 43 3c 39 3b 3d 33 36 38 3c 3b 40 3d 37 3c 37 3d 3f 41 35 3b 3b 3c 3a 39 32 3a 30 37 3a 35 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 31 34 39 3a 41 41 3c 35 3e 47 3d 43 3c 38 42 3a 47 3b 42 3d 3d 49 48 47 49 34 39 38 34 30 3e 3e 3b 36 39 3f 3d 3c 38 3c 3d 38 3f 3c 37 3a 38 3b 39 3e 40 36 37 33 3f 41 42 42 3d 33 29 2a 16 09 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 1b 20 2d 38 35 3e 37 38 3d 3a 45 42 3d 39 39 3f 3d 3d 37 39 35 39 37 3f 38 32 3b 32 3b 3a 35 3a 3a 39 3e 44 31 3c 3c 34 3b 38 35 32 36 42 3e 43 4a 4d 50 4c 42 3e 48 3a 3d 40 41 36 37 36 3b 3b 3b 35 39 33 46 3f 40 39 36 3c 35 3b 3a 39 32 38 3c 35 2d 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 27 34 39 36 3a 39 33 38 3d 39 40 3c 3f 48 3c 3f 41 38 41 3e 3d 48 40 47 41 39 3b 41 3e 44 45 3f 35 3f 41 3c 37 3a 38 3d 3d 37 3e 3e 38 42 39 3b 38 3e 39 3b 33 36 3e 41 39 3c 36 31 2b 1c 0d 09 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 15 20 2c 30 35 35 3c 3f 35 46
 3e 47 36 36 35 44 38 41 3b 41 30 38 32 3b 3d 33 39 3a 36 44 3e 34 39 3c 3c 35 3a 3b 35 3c 38 44 45 3a 40 42 3e 54 50 53 56 50 44 4a 49 3e 32 34 3a 37 3b 39 36 37 37 2d 3f 31 37 3c 3d 43 3e 3b 33 3d 3a 3c 3b 37 37 35 35 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 25 36 41 35 40 3d 41 42 3a 40 44 3c 3d 3a 3b 41 47 42 4c 3d 46 3a 3a 35 41 32 31 39 37 3d 38 3c 3d 44 41 3d 3b 39 3f 32 37 3e 28 45 3e 35 3f 35 37 35 40 37 3c 3b 3e 38 38 3a 32 1d 1a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 16 29 30 39 38 35 35 39 42 39 35 3d 37 3e 38 35 3c 3b 3a 40 38 34 39 36 3f 3e 38 3b 40 39 3b 30 39 38 3c 3e 34 36 39 36 39 37 3a 45 45 44 45 51 51 51 46 43 41 39 36 3d 3f 3c 30 3a 32 36 36 2e 37 3e 3e 42 3b 35 39 39 3c 37 3b 3d 3d 36 37 37 2f 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 25 3b 35 36 3c 3c 32 39 39 3f 42 3d 3e 3e 43 46 44 43 37 37 3c 3c 38 3b 3a 3a 3e 30 3d 3b 40 36 38 40 37 3a 44 38 3a 40 39 3d 43 33 36 39 37 30 3a 32 39 3d 3a 36 40 3b 34 35 2f 19 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 1c 25 28 2e 37 32 3c 3c 38 3a 3f 3a 37 47 3b 40 38 3f 3b 39 33 3a 33 39 3e 41 38 36 3a 41 3e 3a 35 38 38 32 39 3b 3f 37 37 39 3a 42 40 42 4c 4a 4b 4d 3d 49 44 39 36 37 3d 35 38 3a 3c 3b 36 3b 33 39 39 39 34 3e 3b 3a 37 33 36 42 37 39 44 43 37 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 38 3d 3c 36 40 34 44 39 34 40 3b 3e 40 3e 43 3b 41 40 38 3f 35 40 34 3d 30 36 36 3d 39 40 43 40 42 3c 38 3d 3f 37 3a 31 3d 38 32 3b 37 44 40 36 42 3b 39 41 37 38 31 25 20 16 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 1b 22 32 38 34 3c 36
 38 3e 3c 38 38 41 36 3b 39 3e 38 40 3e 36 35 36 3a 38 35 3c 33 38 3e 39 40 33 37 35 39 3e 41 3f 3a 3b 3a 45 3a 3d 3c 48 45 41 43 47 46 46 35 3b 3b 3b 34 3e 3e 36 3c 3e 38 36 44 37 3f 3d 3f 35 39 3b 34 3a 34 44 3a 3e 26 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 31 44 3f 3b 3c 34 37 3c 38 3b 3f 3f 38 3d 3a 39 3b 3e 38 3a 35 3b 38 38 3e 2d 3c 41 3e 3d 3a 3d 3d 37 44 3e 38 36 34 3b 37 42 3b 3e 3c 35 3e 3f 3c 39 39 39 34 2d 30 1a 12 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 1f 21 2a 2f 31 31 3b 36 40 37 3e 39 34 41 43 3e 37 41 32 32 36 36 34 34 36 43 33 38 3c 30 38 32 37 32 35 30 34 3b 41 35 34 3d 39 37 40 40 45 3d 4a 3e 3e 43 36 42 3d 3d 30 34 39 3b 39 3b 42 3c 3c 3c 3d 3c 3a 46 3c 3d 34 3f 3d 3b 3c 3e 30 16 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 23 37 3c 39 3e 3d 3b 31 3a 37 39 3b 3b 38 35 3e 37 34 3a 3d 3a 39 39 39 37 30 39 34 34 3a 34 3e 3b 39 3c 33 34 3d 3d 3c 36 36 3a 3b 35 3a 36 40 3a 39 34 33 2d 21 22 1e 15 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 14 25 1d 32 32 39 38 3e 3d 3c 45 3a 3d 34 34 4c 42 3f 3e 3a 3a 39 38 36 3c 38 3d 2c 35 36 3b 33 3f 42 3f 30 37 37 38 35 39 42 31 3a 38 38 3d 45 40 46 3b 44 3b 44 39 39 42 3a 39 41 41 40 3e 3a 45 42 43 3d 38 3d 38 38 3f 41 3a 3b 42 38 34 23 06 05 03 00 06 05 07 07 06 05 05 03 06 08 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 1f 34 3e 37 41 3a 42 36 3a 3e 44 36 41 32 3b 3e 35 3b 34 39 31 31 3f 3c 43 34 3c 3e 33 3b 41 3a 42 34 43 3a 39 40 3f 41 2e 3c 37 3e 3f 44 3b 39 42 38 3d 31 29 1d 1e 11 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 1b 1e 2a 35
 37 35 3d 3a 3c 40 38 3f 36 36 3c 3c 35 41 3d 3a 38 38 3d 3f 37 3a 3a 3c 32 3e 35 36 34 2e 3a 36 38 38 3d 3b 3a 3c 3b 43 4c 4a 49 43 46 4c 3b 43 44 40 3a 44 3e 42 47 43 48 47 3c 45 3f 3e 41 46 42 3a 40 37 3b 3c 3a 3b 31 1f 06 05 05 03 08 0f 06 07 0b 07 07 10 11 0c 0a 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 23 35 41 3b 44 36 42 3f 3a 3b 3b 37 3b 40 3b 41 35 3a 40 36 3d 3a 38 3b 3d 31 3d 3e 36 3d 3b 3a 3c 3e 44 3f 3d 3b 36 38 35 3c 3c 40 49 3b 3b 41 31 36 3a 2a 19 1f 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 18 25 28 2b 33 30 3d 3d 36 36 33 3b 35 36 32 37 3f 3d 35 3a 3b 37 36 3b 2c 39 3c 41 3e 3c 40 36 38 38 37 37 40 3e 36 35 3a 3b 41 44 3d 3e 43 4a 4e 4e 48 41 3d 3e 46 4c 4b 50 4d 49 55 41 4c 40 40 3d 3d 3f 40 43 3e 35 38 40 33 34 1f 06 05 07 09 0b 0f 0a 15 0f 14 14 17 14 1b 10 18 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 38 38 2d 41 3e 36 34 36 3b 3e 31 2e 31 37 3b 39 33 3b 3c 3e 3b 41 35 35 38 36 39 32 3a 44 39 3b 3c 40 3d 3d 32 3c 40 41 40 3f 41 41 47 3f 37 33 32 2c 1b 13 0d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 1a 1f 28 30 2c 38 36 3e 34 3f 37 40 3d 44 38 3a 3b 37 37 39 42 30 36 36 29 3a 36 38 36 37 37 3b 3b 3e 38 3c 38 3b 3b 43 39 3e 42 3b 44 4e 4a 54 59 4e 4c 42 41 4e 52 59 57 56 59 56 55 54 3d 45 39 41 44 3d 3c 40 41 35 3d 3c 41 2a 14 0a 05 08 15 18 20 1f 1d 22 22 21 2b 2d 2b 20 1b 17 06 09 06 05 03 00 06 05 03 00 06 05 03 21 37 37 43 3e 3a 35 2f 31 3e 39 36 31 37 31 32 33 33 36 35 3e 3b 43 3c 37 3c 30 3a 3e 43 3c 3c 40 3a 38 39 3d 44 41 46 38 3c 44 3b 3d 3e 44 2f 29 2d 1e 16 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 13 1c
 21 2c 2d 33 34 35 3e 3e 3b 3e 36 3b 39 40 3e 39 42 3d 37 3a 3f 34 35 39 35 36 40 39 39 3b 36 33 39 38 3c 40 3a 3d 3b 3a 44 42 44 4b 4a 60 55 5a 5a 4c 50 5d 62 5f 5c 5f 50 53 4a 43 3e 3c 44 43 4d 45 47 40 3c 3d 3c 3e 41 31 19 10 09 0d 1d 25 31 2d 32 34 36 41 3f 3f 3c 3e 30 23 19 07 06 05 03 00 06 05 03 00 06 05 03 27 37 43 44 3e 3a 34 3c 3b 3c 35 33 36 36 37 34 3e 33 3b 35 31 2e 34 39 35 3d 3c 3f 4a 3b 3a 44 36 3e 3b 34 3e 35 39 3f 3e 3d 47 3f 41 38 37 2c 28 22 0c 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 09 14 12 20 2b 2d 39 38 36 38 3c 3b 38 39 36 42 3c 36 3d 3a 3e 3b 31 38 36 36 34 3c 33 38 3b 41 3b 37 37 3f 3b 35 38 37 3e 3f 45 3e 44 46 4d 5d 54 55 55 4d 4b 58 4f 5c 64 52 50 4c 47 45 39 45 40 40 45 41 3d 46 40 3e 44 45 44 39 1d 16 15 1b 27 36 3b 44 3b 44 45 54 57 4a 4d 3c 3b 2e 1b 15 06 05 03 00 06 05 03 00 06 05 03 1b 31 3f 38 35 3d 3e 3c 38 35 25 33 31 32 39 30 39 34 32 3d 3f 36 44 3a 3b 39 3e 47 43 42 3e 3b 38 31 36 3c 3e 3e 32 34 36 3f 40 38 35 35 25 22 18 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1c 20 23 2f 31 32 35 41 34 39 43 3d 3c 38 3b 40 3a 3f 3f 39 33 3d 3b 39 2f 34 38 38 39 37 34 38 36 36 3d 38 39 37 3a 3f 3d 42 46 4d 54 4d 53 4a 45 46 46 50 50 51 4b 4b 3d 43 46 3c 3e 43 3a 3c 3c 46 46 44 4f 4b 46 4a 44 2c 24 23 30 38 48 4a 55 55 57 5f 68 60 54 49 4b 3e 28 19 0b 07 05 03 00 06 05 03 00 06 05 03 1f 31 3f 3b 3e 35 3b 2a 2d 29 35 2f 2e 37 35 37 33 30 3b 3e 38 3b 3a 32 39 3e 39 3b 42 3c 31 37 38 3a 33 39 39 2f 3b 3e 3b 35 31 30 2e 26 1e 13 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 0e 15 18 22 2a 31 2f 37 3a 42 44 39 42 3a 37 47 3e 42 3f 39 3d 36 33 3e 3c 3e 39 38 35 39 42 41 3f 44 3c 41 3a 39 41 3a 3c 45 41 4b 48 43 49 51 4e 4e 50 4c 49 43 46 3a 41 43 41 38 41 42 44 40 45 51 4c 4e 52 58 5e 5a 4e 38 34 34 3e 46 54 5a 5f 62 67 66 68 6d 67 5d 4e 39 30 21 11 06 05 03 00 06 05 03 00 06 05 03 17 2b 37 2e 31 3d 35 34 34 39 37 30 31 33 37 32 36 39 3b 37 37 34 44 3a 34 33 33 3e 34 37 38 3a 37 33 32 40 33 3a 39 31 29 30 30 26 23 15 0a 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 14 19 27 2d 34 35 38 36 3f 3d 41 3e 40 38 39 3a 3e 38 35 44 35 3f 39 37 33 34 3d 3b 3c 41 36 38 42 36 3b 3b 3d 3f 3b 46 42 44 47 49 4f 48 4e 4e 46 50 4e 4d 3e 3f 3f 3d 44 3d 45 3e 40 47 4c 53 54 60 5b 6f 6c 66 56 4a 48 44 45 55 64 66 64 6b 63 6a 74 73 5d 57 4c 35 2a 1f 15 06 05 03 00 06 05 03 00 06 05 03 10 2d 38 2d 2f 2e 2e 35 36 2c 35 33 2e 30 38 26 30 36 36 3b 30 39 3f 3c 3d 3d 33 3c 35 38 39 36 36 36 40 37 2a 3c 34 3a 2e 23 25 22 0e 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 17 1a 1c 30 2e 3c 3a 3a 3a 3f 47 3e 3c 36 3d 41 42 3f 36 36 33 33 3a 3c 35 39 39 3d 3c 3e 3d 39 34 3f 40 3b 42 42 42 49 43 41 42 4a 45 42 42 3f 42 44 45 44 3b 3d 3b 3c 46 42 4f 4e 50 56 64 6a 68 7a 7f 77 73 57 50 52 5b 67 69 65 6b 66 6a 6a 6f 67 64 5a 52 37 2c 1a 0d 0a 05 03 00 06 05 03 00 06 05 03 10 2b 36 31 38 2d 2a 33 30 29 35 30 35 35 38 35 32 38 38 30 35 37 3f 42 3d 30 3b 2f 3b 35 32 40 36 3b 30 35 34 33 2f 2e 2d 29 1d 06 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 11 12 20 21 2c 33 38 37 3b 38 40 3e 41 3f 3e 40 43 37 3e 3b 37 3e 3a 36 3d 39 3e 40 39 40 44 3b 3e 41 3c 48 39 47 45 3e 42 3e 46 4d 49 4a 44 45 46 43 45 41 3b 40 41 3d 4b 41 49 4a 51 68 72 7b 84 92 91 98 7d 5c 63 65 69 74 6e 66 60 64 67 69 67 67 65 55 4b 3c 29 1c 0e 06 05 03 00 06 05 03 00 06 05 03 10 28 3a 2b 2c 33 34 2f 2f 32 31 36 2f 2d 36 33 3e 38 3a 39 37 42 3d 3e 3f 36 39 3b 3c 3a 3f 41 3f 3b 37 34 34 33 2a 2e 22 1f 12 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0b 11 17 29 26 2d 34 30 43 3b 39 42 38 3e 3b 46 42 3c 39 3e 3e 3e 36 3d 3a 3b 43 42 39 43 44 42 42 45 41 42 46 3a 43 48 46 44 44 44 49 49 41 49 41 40 44 48 39 3b 44 46 3d 47 57 61 69 73 86 91 95 a5 9a 8a 6a 65 65 72 6e 6a 69 67 64 62 6d 5e 5a 59 49 3a 2c 1f 0e 0a 06 05 03 00 06 05 03 00 06 05 03 10 2e 34 29 28 34 30 32 38 2e 36 29 30 31 34 39 38 3a 30 37 39 3b 3d 37 3f 3c 37 39 31 3a 38 41 38 3a 38 38 38 33 21 22 16 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 10 18 25 29 36 3d 34 39 38 43 40 41 3d 32 3e 41 46 3c 34 3f 39 3f 3e 40 41 3f 3b 47 42 3c 44 45 4c 4a 4f 4d 44 48 45 4e 45 45 46 43 43 48 43 36 3a 41 44 39 47 4d 47 56 64 72 80 88 96 a1 a8 a4 91 7c 71 6d 66 68 6b 68 5f 62 57 58 5e 4d 49 3a 35 26 13 05 02 06 05 03 00 06 05 03 00 06 05 03 08 25 2e 2b 34 30 30 23 2f 32 30 30 2e 33 31 2c 36 36 3a 37 39 40 44 3d 3f 39 36 32 3a 38 39 3a 35 39 34 32 22 18 18 11 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 06 10 15 1c 26 2e 30 35 36 3c 44 3e 3d 40 40 42 4a 42 41 3d 34 42 40 44 4a 41 45 47 4a 49 4a 55 45 4e 53 54 4e 4c 4b 4d 57 55 5a 4f 53 50 4c 4e 44 40 47 41 44 4c 49 52 58 67 74 7a 90 96 ab b0 ac 9f 89 80 74 6a 70 68 66 60 67 59 58 51 51 49 3b 31 23 17 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 1d 37 30 35 31 33 32 2d 38 31 35 30 32 35 38 39 38 34 3c 3e 39 44 40 3c 36 36 33 36 35 38 38 2e 2d 20 1b 1b 12 0f 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0d 14 1e 25 2d 2c 3c 36 3f 3e 43 45 47 49 43 4c 44 4a 4b 4b 4c 4d 4b 53 56 47 57 58 52 55 61 66 68 61 6c 5f 64 61 60 6a 66 5c 62 57 57 56 4f 4e 4e 4f 49 49 5a 53 66 73 84 8b a0 b2 af a7 a6 8f 84 78 75 69 71 66 6d 60 61 58 53 48 43 3c 29 15 10 06 00 06 05 03 00 06 05 03 00 06 05 03 06 23 2e 2e 2c 33 2d 30 34 31 35 32 35 37 3a 39 39 37 40 40 3b 39 38 36 3d 35 2f 2d 2f 2f 39 2b 24 1e 1d 1b 11 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0f 23 1f 24 34 3a 44 41 4e 4a 44 55 52 55 50 52 55 50 5a 56 60 57 5f 67 5e 60 69 69 6f 74 75 79 76 74 77 74 74 76 71 74 6e 6f 69 65 5e 65 62 59 5c 55 57 5c 63 72 7b 8c 97 a3 ab aa aa 8d 89 7a 6a 6c 64 62 62 5b 62 4e 50 47 46 31 21 19 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 03 27 35 2f 34 2d 31 39 38 32 35 31 33 35 33 38 32 33 39 36 3d 35 34 35 30 30 27 2b 2c 22 2a 25 1a 14 0c 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 0f 1d 23 2a 36 44 41 4c 4b 50 5a 60 5f 5b 5e 65 64 6a 61 65 6b 74 6c 71 76 75 7f 78 7d 7d 79 80 7c 7f 83 79 81 7d 76 79 7c 7e 76 6e 77 77 7a 6b 6a 68 68 71 74 7f 85 95 98 ab ac a1 8d 82 7b 7d 7a 6f 67 5f 5c 5c 5a 50 50 40 2d 20 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 07 24 34 28 30 35 35 2e 34 30 34 30 37 38 3f 33 39 30 30 39 39 29 31 29 32 2a 2b 28 21 22 22 1a 16 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 17 17 22 31 3a 42 4d 59 5c 69 63 6a 64 69 6f 6c 74 77 78 77 74 78 7a 7b 76 7d 7c 7e 7f 82 80 7c 79 80 82 7c 82 86 7c 81 7b 82 7e 7e 84 82 85 7b 79 7e 7c 7e 84 8c 91 a0 a4 a8 a1 95 7f 7e 77 76 6f 73 60 57 62 57 5e 4a 3a 32 1f 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 1b 34 2f 2c 2d 31 32 2e 40 3b 2a 31 3c 33 35 35 33 39 38 2f 2f 34 2f 2a 2a 20 23 28 14 14 0d 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 17 1c 31 40 46 56 5e 64 6e 63 6a 6c 69 6d 72 73 74 73 75 7c 7c 76 7f 7c 74 72 7e 78 7c 7f 80 7a 77 74 7c 7e 89 7e 79 87 7b 7b 7b 85 86 85 84 83 82 85 8c 92 8f a1 a3 a8 aa 8f 7a 73 6d 70 70 5f 5d 5f 62 58 53 4d 44 2c 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 24 37 2d 30 30 30 32 36 37 39 30 2b 33 35 34 33 2a 33 31 30 2a 2d 2d 2d 20 19 15 1a 13 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 1d 1f 34 42 49 54 64 63 62 62 61 6b 73 70 6f 6e 70 74 7a 7d 73 70 75 75 74 7d 78 77 6a 75 7a 79 7f 83 77 7f 79 7d 7f 80 78 7b 7f 81 86 86 88 86 86 95 8b 94 a7 a1 a6 a2 84 6a 62 61 66 6f 6c 66 67 5b 55 4b 42 35 2c 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 21 3b 37 35 39 34 35 2e 35 2c 35 33 32 2e 34 2a 25 28 33 34 2a 28 21 27 1e 14 12 12 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 1d 2f 39 4e 58 58 5e 61 69 6b 6b 65 66 72 6f 74 6d 76 75 74 7a 71 76 72 70 79 79 72 7b 71 74 77 75 76 7b 79 77 7f 82 86 85 83 83 79 84 83 86 89 90 91 a4 ab a2 a7 81 5b 5a 57 5e 67 66 6c 6e 5c 55 46 41 36 29 15 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 22 38 35 31 3a 39 2e 3b 30 35 32 2d 2e 32 2c 2f 30 2c 29 27 2c 28 1b 16 12 14 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0a 16 2a 34 49 5d 5a 61 5b 60 60 65 62 69 69 63 59 6f 66 6c 6a 69 6f 6f 72 6d 72 6a 6e 6e 70 78 71 74 79 6e 76 71 73 79 7d 7b 72 77 80 80 8b 84 8c 88 97 9d 93 99 75 46 42 4e 51 5b 69 66 62 65 5b 4a 44 3a 23 18 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 3d 2d 44 3c 2d 30 2d 30 39 39 2f 2c 2e 2e 2b 28 2b 2d 22 1e 22 12 13 13 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 13 1b 22 2f 3f 4d 58 59 5f 5a 60 5e 63 67 68 62 5b 60 65 66 6f 64 5f 65 60 6b 6a 68 65 6f 67 6f 72 70 67 6e 73 7a 81 74 72 78 78 78 7b 7c 7c 7a 85 89 84 8c 80 5e 40 40 49 49 56 55 67 67 6d 65 58 39 2a 1e 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1c 35 3c 36 2c 35 2a 2b 31 27 29 31 26 26 2d 24 2d 2c 20 1e 11 13 07 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0d 16 26 33 44 48 49 52 57 62 5e 5e 5f 60 60 5c 63 5e 61 58 62 61 60 64 65 5f 62 5f 64 64 68 6c 69 5f 6b 6d 77 75 6d 73 6d 75 71 75 76 78 7c 81 82 78 7c 77 5d 30 36 38 48 50 5f 62 66 6f 67 5f 43 28 19 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 28 3a 3d 3d 34 2e 2e 2e 2b 29 29 23 2d 27 29 15 22 1a 16 16 12 06 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 17 1d 2e 32 41 44 4e 53 59 5a 60 5b 52 5a 58 5d 60 5b 56 5f 5b 56 59 5d 60 60 5c 5e 62 62 69 66 66 64 6d 6a 65 73 6d 6b 73 6e 6c 70 68 77 71 78 73 7b 55 20 25 26 3c 46 56 56 57 65 61 50 48 2d 15 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 26 45 3d 3b 36 27 2a 2d 24 25 22 22 1d 21 1f 18 15 10 05 08 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0b 13 24 33 2f 3b 52 4c 51 54 5a 59 57 51 53 56 52 51 55 57 5c 4f 57 51 56 54 51 59 5d 5e 5f 63 62 60 66 67 6e 64 6f 63 63 6a 69 70 6c 66 6f 65 69 47 18 0b 21 2d 44 4e 50 5e 5e 52 4e 42 1f 14 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 27 40 35 3a 2d 1b 24 25 1a 26 1d 14 14 12 11 07 08 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 08 15 27 2d 3a 34 3c 43 53 51 4c 4b 55 56 52 52 54 4e 4a 52 4f 56 53 4f 4b 4c 53 57 58 54 5f 55 63 62 5a 60 60 69 60 63 61 67 67 60 66 64 62 5c 40 15 0a 16 1e 36 4a 46 53 54 53 4a 38 25 0e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 28 3b 34 2e 26 20 19 1f 1f 22 11 15 06 06 04 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 10 0f 21 2f 3d 37 3e 44 48 4e 4f 45 47 45 4a 4a 4b 4a 3e 42 4d 49 3f 47 49 52 51 54 58 5a 4d 5a 55 5b 5f 56 59 57 60 5e 54 5f 53 57 56 52 3c 0c 04 06 1d 2e 3a 45 45 51 47 41 2a 1d 0d 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 24 1d 18 0d 06 0c 08 14 06 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 0a 18 29 23 2e 3a 33 3a 3e 3c 44 3f 3e 41 37 37 2f 38 36 34 38 3d 43 49 4e 46 4b 42 47 4b 41 4f 52 53 4f 4a 4c 50 4a 49 4f 47 46 3d 2c 06 03 00 07 1b 20 2f 36 3a 31 28 1f 1b 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0f 0f 22 24 35 33 2e 35 38 30 2e 2d 23 25 1e 2a 2b 27 2b 39 42 3c 41 42 39 42 3c 3f 3f 45 4a 45 3f 3b 3a 3a 3b 3a 39 39 33 27 1e 05 03 00 07 0e 10 22 24 29 23 1d 15 08 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 12 1c 1d 23 21 22 20 1a 14 16 10 0e 12 1d 17 24 22 31 33 35 32 26 24 2a 29 23 2f 29 25 30 2a 2a 29 28 1e 22 23 17 11 07 05 03 00 06 10 0e 0e 16 15 16 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 05 06 05 0b 0b 06 05 03 00 06 05 09 08 15 16 1b 1c 14 19 15 0d 0d 19 17 1e 10 14 18 0f 1b 0c 10 0f 12 0e 03 00 06 05 03 00 06 05 03 07 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 08 0b 07 0b 05 02 06 09 03 05 06 0d 03 05 0b 05 04 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
