 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 05 03 02 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 07 00 06 05 03 00 06 05 05 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 05 01 09 05 05 0a 06 05 08 00 08 07 03 02 06 05 03 01 06 07 05 04 08 05 07 09 06 05 03 0b 06 05 07 06 06 05 03 02 06 05 03 09 07 05 03 06 06 05 03 06 08 05 03 00 06 05 03 06 06 05 03 00 06 05 03 09 06 05 08 08 06 05 03 00 08 05 03 06 06 05 03 00 06 0e 07 00 06 05 03 06 06 05 03 00 06 05 04 01 06 05 04 00 06 05 03 01 06 05 03 07 06 05 04 00 06 05 03 00 06 05 05 00 06 05 03 04 06 05 03 00 06 05 03 0a 06 08 07 00 06 05 03 02 06 05 0c 05 06 05 03 03 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 05 06 05 03 06 06 06 04 01 06 05 07 00 06 07 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 02 06 05 05 04 06 05 04 06 07 05 03 0d 08 05 03 00 06 05 03 0b 06 05 07 03 06 0b 03 00 06 05 03 02 06 05 03 04 06 05 03 05 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 05 06 05 03 00 06 05 09 01 06 0c 03 00 06 05 07 00 06 05 03 00 06 05 03 06 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 00 06 07 03 00 09 05 07 02 06 05 03 00 06 05 04 07 06 05 0a 01 06 05 03 00 06 05 04 04 06 05 03 01 06 05 03 05 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 04 06 05 03 03 06 05 03 07 06 0a 05 07 06 05 0b 06 06 06 03 02 06 05 03 00 0a 05 03 04 06 05 05 06 06 07 03 05 0a 05 0c 03 08 05 03 01 06 06 09 0e 08 05 09 0c 07 07 06 00 06 05 06 06 06 06 03 07 0b 05 03 01 09 05 03 03 06 0b 05 01 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 02 06 07 03 07 06 05 0b 04 06 06 03 06 09 05 03 00 06 05 03 08 06 0b 04 10 08 09 0c 03 06 05 03 06 06 09 03 06 06 05 03 04 06 05 03 00 06 05 03 00 06 0a 03 07 06 05 03 09 06 05 07 02 06 05 03 00 06 05 03 08 06 05 08 06 06 05 07 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 03 08 06 05 10 0c 09 08 0c 02 06 05 03 01 08 05 03 02 06 05 03 00 06 05 06 0a 06 05 0f 06 06 05 04 04 06 09 0e 00 06 06 08 05 06 05 05 0b 06 0d 04 0e 06 05 04 06 06 05 08 00 06 09 03 08 06 05 04 00 06 05 05 05 06 05 03 03 0a 05 03 01 06 05 03 01 06 05 03 04 06 08 03 00 06 05 05 04 06 05 05 06 06 0b 03 06 06 05 03 00 06 05 03 03 06 06 0a 0a 09 0e 09 04 06 05 03 06 06 08 05 00 06 05 03 00 06 05 07 06 06 05 03 03 06 05 03 00 06 09 04 02 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 02 06 07 06 04 06 05 03 08 06 05 03 03 06 05 04 04 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 07 05 00 06 06 04 01 12 0c 0c 04 06 05 10 03 08 05 03 07 06 05 08 05 06 05 03 07 06 05 03 05 06 05 03 00 06 05 0a 00 06 05 03 03 06 0a 05 0d 07 05 04 0a 07 05 04 01 06 05 03 07 06 05 03 09 08 05 03 04 06 05 03 13 06 05 06 07 06 05 03 00 06 05 03 00 06 06 08 02 06 05 03 0a 06 05 03 07 06 05 03 01 06 05 03 00 06 05 03 04 06 05 03 00 06 05 06 07 06 05 05 00 07 05 06 01 07 09 08 08 06 0a 03 08 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 06 06 06 06 04 06 05 03 00 06 05 05 03 06 05 03 05 06 05 06 00 09 0a 06 00 06 05 08 01 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 07 04 06 05 03 01 06 05 04 09 06 05 0e 09 06 0a 07 0f 06 05 09 01 07 05 05 02 07 05 03 09 06 05 04 00 08 05 03 03 06 05 03 02 06 05 03 01 06 05 03 07 06 07 05 09 06 0d 06 0a 06 05 04 0a 06 05 06 0b 06 05 04 05 06 06 04 09 06 08 05 05 06 0b 06 07 06 06 08 00 08 05 03 00 06 05 03 04 07 07 03 02 06 05 03 00 06 05 04 02 0b 08 03 00 06 05 03 00 06 05 03 01 09 08 0b 0f 0c 05 08 07 06 05 06 04 09 05 07 07 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 0e 06 05 03 01 06 05 03 02 06 05 03 02 06 05 03 06 06 05 03 01 0c 09 05 06 06 05 03 02 09 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 01 06 05 04 00 06 05 03 03 0d 06 09 03 06 09 06 00 06 0c 12 09 0d 0d 07 0b 0a 05 09 0a 06 05 06 08 06 05 03 0a 06 05 05 09 06 05 0b 00 07 05 05 0b 0f 06 03 06 06 05 06 0d 06 0d 09 0b 0c 0a 09 07 09 05 08 10 06 07 06 02 06 0b 0a 01 10 05 03 0a 06 0d 09 01 07 05 05 03 06 05 03 02 06 05 07 00 06 05 03 00 06 05 03 06 06 05 03 07 06 05 03 04 06 05 08 03 06 05 03 01 06 05 03 03 0a 05 0a 06 06 09 12 05 09 05 06 06 06 05 0b 02 06 0a 03 06 06 05 04 04 06 05 03 00 06 05 03 0b 06 05 03 01 06 05 03 00 06 05 03 07 06 05 03 00 06 05 03 00 06 07 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 05 03 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 04 06 05 07 05 06 05 05 03 07 05 03 04 07 06 09 0f 0d 06 0f 0c 06 08 03 01 06 05 0e 01 06 0e 03 01 06 05 03 06 06 05 03 00 06 06 08 08 07 05 08 02 06 06 04 04 06 0d 04 08 06 08 03 07 0d 0a 03 0a 06 05 03 0a 06 05 0a 0a 06 06 03 00 06 05 03 09 06 08 03 07 06 05 03 01 06 05 03 00 06 05 03 01 08 05 0e 01 06 07 03 00 06 05 03 05 06 05 03 02 06 05 03 00 09 05 03 0a 06 0a 0b 01 12 08 03 00 06 05 06 00 06 08 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 0b 04 06 05 03 01 06 05 03 01 06 05 03 01 06 05 06 02 06 05 03 01 06 05 07 04 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 05 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 08 06 05 09 01 08 05 0c 0d 06 05 03 0b 06 10 11 11 0c 12 07 12 0f 09 0a 08 06 05 08 0b 06 05 09 06 07 0c 09 03 06 05 09 0b 06 0a 0c 04 08 09 0c 0c 06 06 06 08 0d 09 0c 0b 06 10 0b 0e 14 07 08 04 06 0a 03 0d 08 05 0e 03 09 09 0b 06 06 05 03 08 06 05 03 03 08 05 05 02 06 05 03 00 06 05 03 07 06 09 04 02 0a 05 03 09 0b 05 03 0a 06 05 03 0b 0d 05 03 02 06 07 0a 0b 06 11 07 10 0f 0f 0a 03 10 08 03 04 06 06 08 04 0c 05 03 02 06 0b 03 06 07 05 03 00 07 08 03 07 08 09 03 07 06 05 03 04 06 05 04 00 08 05 03 00 06 08 03 04 06 05 0a 03 06 05 03 09 07 09 0c 04 06 05 03 08 06 07 03 08 06 08 03 08 06 05 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0b 07 0a 09 05 06 04 06 05 0d 13 13 0c 11 17 06 0d 0e 0a 06 10 0e 0a 0c 05 08 07 06 0a 07 0c 06 05 0f 05 06 05 03 09 07 08 04 08 06 08 10 0d 07 0f 08 12 0d 10 0c 17 12 06 06 09 06 05 08 06 06 0a 10 10 0e 09 10 07 06 08 05 06 07 05 03 04 0a 05 03 06 06 08 09 0b 06 07 0a 04 06 05 0c 09 07 05 03 01 09 05 03 03 06 08 03 00 06 05 03 04 07 07 0d 00 0d 05 0c 0e 11 05 0c 0d 0a 0e 0f 05 0a 0f 07 08 06 05 03 02 06 05 03 03 06 05 04 05 06 05 03 05 0b 05 04 06 06 05 09 00 06 05 03 04 06 05 03 00 06 07 03 03 06 05 0a 04 06 05 0c 05 06 07 06 02 06 05 03 07 06 05 04 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 06 05 06 09 06 05 03 00 0b 0b 09 00 0d 0d 0d 14 0b 0f 14 0a 0b 0b 0e 0d 0b 05 10 0d 08 05 0a 0e 06 06 0c 09 06 05 05 07 06 06 08 12 13 09 0a 06 06 09 06 06 06 05 03 08 08 13 0d 11 06 11 0a 0d 0f 07 0a 07 07 09 0d 06 08 0e 09 04 0e 07 07 0f 06 0b 03 07 07 05 03 00 06 06 05 09 0a 05 05 05 06 09 04 05 06 05 05 03 06 05 03 07 06 05 03 00 06 05 03 03 06 05 07 0a 06 0c 0a 0b 0f 0e 05 0b 08 0a 09 04 06 05 06 02 06 09 03 01 06 05 03 06 06 05 03 00 06 05 0e 00 06 05 03 05 06 05 03 0a 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 05 03 00 06 05 05 00 06 05 03 02 06 05 06 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 03 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 02 06 05 03 00 06 05
 03 02 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 04 07 09 06 07 06 10 0b 07 0f 0b 13 13 11 13 14 0f 0a 0d 0a 0b 0f 0d 14 08 0f 0a 05 0d 0c 08 05 07 0c 0a 05 09 00 09 05 0a 0d 0b 0b 06 0f 08 05 0c 07 0d 06 11 0e 0d 0e 13 10 0d 0a 04 0c 09 0d 06 0c 0e 0d 09 0e 06 11 0e 07 06 0f 07 0d 07 0e 03 09 09 09 0a 02 09 05 0a 00 07 05 03 03 08 0e 03 09 06 05 03 05 06 06 03 0b 06 05 03 06 07 05 03 01 06 05 0e 0a 0a 0e 05 08 08 0a 0b 07 06 07 07 11 06 05 05 07 06 05 06 00 06 05 05 02 06 05 03 09 06 05 07 0a 0a 05 06 04 06 06 03 00 09 06 04 01 06 05 04 00 06 05 08 09 06 05 06 07 08 05 03 00 06 05 08 00 06 05 03 00 06 05 03 07 06 06 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 03 02 07 05 03 05 06 05 03 00 06 05 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 07 05 03 04 06 05 03 08 06 05 04 04 06 05 05 00 07 07 06 09 0a 09 0b 07 0b 08 09 14 0e 0d 13 12 1b 13 0b 14 10 17 0e 14 10 07 10 05 08 07 0e 0c 0e 0b 0d 10 09 10 10 0b 0b 05 04 04 17 10 12 0b 09 0d 0e 0e 0e 07 16 07 12 17 07 0c 06 06 0a 14 09 05 09 12 06 10 07 10 18 09 0a 0b 0e 08 0a 0a 06 0a 03 09 12 05 09 07 08 07 05 01 06 05 05 11 0b 0c 03 00 09 05 0a 07 06 09 03 04 06 06 03 03 07 05 07 04 06 08 0f 0a 06 05 0d 0e 11 0e 08 06 0f 05 03 11 06 09 0f 02 06 05 05 08 06 05 03 00 06 05 03 01 06 07 03 04 0b 0b 06 0a 06 06 05 00 06 09 03 05 06 05 03 05 06 05 04 01 06 05 05 01 07 05 03 05 06 05 05 01 06 0e 03 05 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 03 06 05 03 00 06 08 03 03 06 05 03 02 06 05 03 02 06 05 03 00 06 05 0a 0a 06 05 03 04 0a 0b 0a 0b 06 07 08 0a 06 05 11 10 15 14 0c 0e 0f 09 0c 0e 0d 0c 05 09 06 07 0f 11 0d 0b 1b 0d 0b 08 06 0a 0f 0e 0f 0f 10 12 0d 07 06 09 07 07 11 18 0f 12 09 11 0e 0f 10 18 0c 0f 09 06 08 04 0f 06 0e 14 11 19 05 0c 0a 09 0f 10 0a 0d 0d 10 07 07 09 09 06 06 03 02 0b 05 03 05 06 08 07 01 06 10 04 05 06 05 03 00 06 0b 03 09 06 05 04 0a 06 0d 0b 05 06 14 05 0e 06 05 06 06 0d 0f 09 09 10 05 07 06 06 05 04 02 06 06 05 00 06 05 03 0d 06 05 03 0a 06 05 03 03 06 05 03 03 06 05 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 07 06 05 03 00 06 05 04 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 09 05
 03 09 06 08 03 02 06 05 05 00 06 05 03 01 06 05 06 02 06 05 03 03 0c 05 03 01 06 05 05 0a 09 07 11 0c 10 11 11 08 0c 12 14 0d 17 10 1a 16 08 11 13 14 16 09 0c 16 15 0d 11 06 06 13 0b 0a 0e 12 0e 06 0d 09 16 0e 19 12 05 09 0f 12 10 11 09 14 0c 11 11 1a 15 0e 0d 12 13 13 06 12 0e 0b 0a 0f 11 18 13 1a 03 10 12 11 19 13 0c 0d 0a 10 0c 05 16 0e 09 0c 07 00 06 09 04 07 06 05 08 10 06 05 07 05 08 05 0e 0c 06 09 08 0d 0c 06 0b 05 06 0c 10 05 0c 0a 16 0e 0d 05 0a 0e 0e 0a 0c 10 0f 05 0e 04 06 06 03 00 06 05 03 07 06 05 03 00 06 09 08 08 06 05 03 07 06 05 06 04 07 05 03 05 06 05 08 00 06 05 03 03 08 05 08 00 06 05 03 06 06 05 03 02 06 05 03 00 06 05 03 09 06 05 03 05 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 04 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 05 06 05 0b 08 06 07 06 02 06 05 06 02 07 08 03 0b 06 05 03 01 06 05 03 08 06 05 03 02 0a 07 0a 00 06 09 0a 18 06 0f 09 0e 07 1d 0a 17 12 1f 17 11 19 12 1b 15 1c 1c 13 13 11 09 18 0a 1a 0b 0f 18 11 13 19 11 13 0a 10 0f 0c 0e 12 0f 10 14 1b 13 11 11 13 10 0e 12 16 0e 15 13 12 1b 11 14 0d 17 10 10 15 11 11 18 1d 11 16 16 0f 19 16 1b 14 13 10 1f 11 11 13 15 0e 0c 0e 05 0e 07 08 05 0d 03 06 0e 0e 06 0f 08 07 0b 06 08 0a 0b 07 0b 03 06 06 0d 09 0a 11 0a 12 12 14 0b 0b 14 10 0a 06 0f 0d 08 0c 02 06 10 0a 01 06 05 03 0b 08 05 04 0a 06 05 03 06 06 0a 07 06 0b 11 0b 09 0a 09 09 03 06 05 03 00 06 05 03 03 06 05 03 03 06 05 0a 07 07 05 07 06 08 05 04 00 06 05 03 06 06 05 04 01 08 05 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 08 04 06 05 03 06 06 05 05 00 06 05 03 09 06 05 05 06 06 05 03 00 08 05 06 00 06 05 03 00 06 05 03 0b 06 0b 0b 06 13 0a 0e 19 08 05 03 04 06 05 03 01 09 05 03 00 0e 09 04 0f 0d 0b 0b 0a 0d 15 12 11 12 11 09 0e 13 17 18 1a 13 13 1c 17 16 19 0f 15 0e 11 08 18 0b 15 13 09 16 0b 19 12 13 13 0b 09 10 1b 10 17 17 19 10 18 19 13 19 14 11 1f 18 0e 10 15 0f 17 1a 08 15 19 11 1a 16 1a 14 1b 13 14 15 16 15 13 18 18 13 13 11 1b 18 15 11 13 0c 0d 0b 08 08 14 0d 12 0a 0b 06 0d 07 09 10 0d 06 09 09 0a 0b 02 08 0b 0f 07 0b 0b 03 0b 06 0c 13 13 11 13 0b 07 0a 15 15 0c 07 06 08 0a 06 0e 0c 0c 0a 05 0a 09 06 07 03 09 06 06 0a 0d 06 08 04 0f 06 0a 05 02 0a 06 04 06 07 06 03 01 06 05 0e 01 06 06 03 02 06 05 03 00 07 06 03 01 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0b 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 04 06 05 03 05 06 05 03 03 06 05 03 00 06 05 03 00 06 05 06 08 06 0b 03 03 06 05
 03 04 06 05 03 0a 0b 11 12 16 0d 0e 05 0a 06 09 04 00 06 05 07 08 07 05 03 08 0b 12 0c 0e 10 0d 12 15 19 0f 0a 0f 15 14 14 19 1e 20 1c 19 15 16 14 0e 12 18 12 1a 16 15 1c 14 18 14 10 12 15 16 16 13 0e 11 13 15 13 1e 18 1a 1c 19 1d 11 14 12 13 17 13 1d 1b 18 10 17 13 1e 17 19 10 17 1d 16 1a 1a 1e 1a 1c 12 21 1b 1a 1a 1e 16 17 1f 19 1f 0b 19 09 15 14 0c 15 12 15 16 10 0b 0b 10 15 10 0c 0e 06 07 08 0b 06 10 0a 06 13 05 0f 0c 13 13 1c 0d 13 13 13 10 12 0d 13 0c 0c 0a 05 07 07 0c 09 05 06 0b 04 00 0d 0c 08 09 06 05 03 05 09 08 0b 0d 0c 0d 03 06 0b 06 03 0c 06 06 03 00 06 05 03 08 06 05 03 06 06 05 03 00 06 06 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 02 06 05 04 00 06 05 03 02 06 05 03 02 06 06 03 05 06 06 08 00 06 05 05 05 07 0b 08 05 06 05 05 04 06 0b 05 01 06 05 03 09 06 08 0a 07 06 08 03 0b 07 0a 0a 0f 0d 0e 0a 0b 09 09 08 0a 07 08 09 06 08 08 0a 0d 10 09 0b 0f 17 10 12 10 14 14 12 18 17 0f 19 10 20 25 1e 1f 1d 1a 18 18 19 22 11 1a 1a 19 1e 15 0c 16 14 1b 21 14 1f 16 15 22 21 19 1f 1a 17 23 3d 44 22 1b 1b 16 19 10 1a 16 1a 1b 16 1c 1c 1c 27 1f 19 12 24 33 29 2b 29 28 28 2a 26 2a 26 2e 20 26 1d 1f 1c 20 22 1b 19 19 11 11 11 1a 1a 18 12 15 15 11 15 1b 12 13 0a 09 0e 0f 11 0b 13 05 0f 0d 0b 11 11 15 11 1b 16 1b 10 0b 15 19 12 14 0e 0e 0a 12 06 0e 18 12 12 0b 0b 07 07 08 09 00 0f 06 03 0b 0c 05 0d 0a 08 11 08 0a 07 05 03 03 09 05 03 01 06 05 03 00 06 0b 06 0a 06 05 04 00 06 05 03 00 06 06 06 09 07 05 03 00 06 08 05 00 06 05 03 0a 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 09 07 05 03 00 08 05 03 00 06 05 03 04 09 05 08 04 06 05 04 00 06 05 05 00 06 05 03 06 06 05 05 07 06 05 07 00 06 05 09 05 07 05 0a 06 08 0b 0f 11 14 08 05 04 0b 05 07 00 06 05 03 03 06 0a 08 0a 09 0f 13 11 15 0f 0b 0c 13 17 1e 17 17 19 15 1c 1d 1d 1e 20 21 21 21 21 1f 19 2a 1f 18 1d 19 16 1c 18 19 1f 19 1d 1f 18 28 24 25 28 2d 31 24 32 39 34 29 23 1e 22 27 21 1d 1d 25 13 1d 1d 20 2d 21 26 25 29 39 3b 42 41 34 37 33 37 36 34 33 3a 33 31 31 28 2b 2f 2d 2e 24 24 20 21 1f 16 1d 13 16 1a 13 17 0f 1d 10 14 11 17 16 0c 13 14 15 13 16 0c 11 10 1b 17 18 16 10 1f 17 18 19 14 0e 12 0e 10 0d 0b 10 0b 11 0e 0a 0c 0e 0a 06 06 08 0e 06 05 0a 09 07 0e 03 08 06 0a 0c 03 06 0a 03 09 06 05 03 01 0a 05 05 0c 06 0a 03 00 0b 0a 04 03 06 05 03 05 06 06 03 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 09 03 00 06 05 03 00 06 05 03 07 06 05 03 10 0a 05 07 00 06 05 03 03 06 0b 03 00 06 05 03 01 06 0a 07 0a 06 0c 05 08 09 09
 07 0b 0b 07 05 11 08 08 05 0e 10 0b 0a 06 06 07 09 01 0a 0c 09 0c 0a 0c 0b 0d 06 0e 0b 0d 0d 1d 19 1a 17 24 16 1d 16 23 23 21 1e 23 1a 22 1f 1e 23 1d 27 28 30 32 27 1e 1b 25 26 23 26 22 26 22 2a 36 35 30 39 38 44 47 2c 27 2e 25 30 2a 25 27 1b 22 27 24 21 2c 25 25 25 29 22 23 2d 37 47 4a 54 5a 4d 48 3f 47 42 46 40 46 43 43 42 4d 42 36 41 3b 36 2c 2a 27 2e 2c 2c 29 2d 39 2f 27 21 22 23 1d 1e 17 1b 18 11 14 0d 15 14 14 1b 19 18 1b 1b 20 17 1f 15 16 14 19 0d 08 0c 11 03 10 14 12 12 17 15 14 0b 12 06 0a 05 0c 0b 0a 05 08 0a 0c 14 10 0c 0d 0e 0e 06 05 04 02 06 05 03 06 07 05 03 05 06 0a 03 0c 06 08 0a 00 06 05 03 05 06 05 03 00 06 05 03 03 06 0a 03 03 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 05 00 06 05 09 06 0c 0b 0b 05 0b 05 03 08 06 05 03 0a 06 05 08 02 06 05 05 05 07 0d 0a 06 06 06 06 03 0a 09 05 06 08 0c 08 06 07 0f 0d 12 0b 05 03 04 0a 14 0b 07 08 06 04 0f 0d 0d 17 18 13 10 15 1a 13 19 19 16 21 22 15 1c 1c 26 27 21 2e 20 26 22 29 1b 29 2a 2c 31 2d 2f 23 32 22 24 36 30 32 23 30 30 31 3e 4d 53 5e 5e 5a 55 3a 2e 2e 30 34 2f 2d 2d 27 2d 32 27 2a 2f 2e 33 26 3d 42 44 4b 52 54 5d 6b 74 74 6a 60 69 65 66 5f 58 50 53 53 65 58 50 3c 4a 49 43 3c 39 45 40 36 40 3e 46 4b 40 3c 34 31 2b 1f 23 28 1a 1d 18 1c 22 20 19 16 1f 1b 1e 1e 22 15 14 17 1f 1b 1c 18 1a 15 0f 0f 16 10 14 12 0f 11 05 10 0d 0b 10 14 0a 06 0a 04 11 0a 0a 09 15 0c 06 0a 0c 14 05 0c 0a 0e 05 0a 07 06 09 0a 07 08 05 03 00 07 05 09 03 06 05 05 04 06 07 03 02 06 05 03 07 06 05 03 06 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 02 06 05 03 01 06 09 0a 0a 0a 05 08 05 06 05 03 07 06 0d 05 04 06 05 04 06 0a 05 03 06 06 08 03 06 06 0c 05 06 0f 05 0a 07 06 0e 08 06 0d 0d 0a 0f 06 05 09 05 10 11 09 10 08 0d 04 12 11 10 13 11 0b 14 11 15 1c 14 1f 1f 25 20 1e 1e 22 26 1b 23 28 24 27 23 22 2c 26 2e 32 36 30 3c 34 37 3e 3a 46 43 44 46 42 49 4e 5e 76 88 85 82 85 87 60 51 51 46 53 44 44 39 3c 38 3a 32 2c 38 35 39 44 53 7a 8b 83 82 78 81 8b 90 87 84 83 81 8e 8e 88 73 6a 6e 62 6b 5d 57 52 50 4f 53 48 4a 46 43 44 4f 5a 5c 5e 60 56 4c 48 3b 25 25 26 31 2e 26 2d 1d 2d 2c 29 21 2d 1b 25 1d 21 1f 19 1e 11 1b 13 1b 18 18 21 11 14 16 13 14 12 12 09 0f 0d 09 17 14 12 0b 07 0d 0b 10 0c 12 06 0f 09 09 0b 09 16 0b 0a 05 03 00 09 05 08 06 06 05 03 03 06 07 09 00 0a 05 03 00 06 05 04 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 08 05 03 09 06 05 03 08 06 09 03 0e 08 08 07 07 0c 05 03 05 06 05 03 07 10 05 03 05 06 09 0a 0a 06 0a 0e 0d 06 0b
 08 0c 0e 0b 07 0a 0d 08 03 0b 06 0e 0b 0c 0b 09 08 0c 09 15 14 14 0d 10 0f 11 11 12 1a 1e 11 1c 1f 1d 17 24 25 21 29 28 2d 2f 29 2d 27 33 36 35 3b 37 48 47 47 51 55 52 58 5d 59 5c 61 65 66 70 76 9a b5 b2 b1 a1 a1 9f a1 93 8b 97 9d 95 90 85 6b 4a 35 3b 3f 5f 69 4f 5b 90 ac b9 a7 a1 a0 95 a2 97 9c 99 91 a1 a6 b4 9b 96 85 82 77 7c 75 57 5c 5c 52 4f 58 50 50 59 53 54 54 60 72 79 78 68 53 51 42 36 41 3e 3c 35 2f 39 3d 3e 3e 41 3d 2f 35 32 1c 23 1b 1a 21 1c 19 1a 10 16 16 1c 20 14 0c 12 0c 16 11 0f 06 07 13 14 12 07 0d 0f 07 14 07 09 0c 0d 09 07 10 0f 09 08 08 05 03 00 06 05 07 00 06 05 03 00 07 05 03 05 06 05 05 00 06 07 03 00 06 05 03 00 06 05 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 04 00 06 05 03 01 07 05 07 0d 06 0b 03 0a 06 0a 09 0a 0b 05 03 0a 06 08 09 03 08 06 06 03 09 05 06 06 06 10 15 04 0d 0e 09 0e 0e 0a 15 13 0a 14 0d 12 10 0c 12 16 0c 0d 15 10 15 19 0d 16 1b 18 16 18 16 1e 20 1e 22 25 23 1e 21 2f 2b 27 21 2f 34 3e 41 43 43 49 4d 54 5a 6e 7c 84 84 85 84 82 8b 8f 8a 86 7a 80 90 9c b1 d8 d6 cd c0 b9 b5 b6 b4 b4 b8 c4 c6 cc cf cb b3 81 51 46 56 96 ad a5 a7 b3 c2 c0 b9 b8 b4 af a6 a9 a3 9a 94 a3 bb b8 ae a3 91 8d 8d 93 9b 79 72 67 66 64 61 6d 66 64 61 61 69 73 7d 85 7d 7b 79 76 69 6c 64 5d 61 5f 54 5e 5d 5e 54 50 4a 49 35 40 36 35 2e 2c 2c 2a 28 26 18 14 23 2e 25 1c 1f 0e 19 16 15 1d 19 0e 12 15 10 0e 03 08 0f 16 12 11 15 13 0d 0e 14 08 0a 0d 08 05 09 02 08 0b 09 0c 06 05 03 0a 06 05 0a 00 06 05 04 06 06 05 04 01 06 05 03 03 06 06 03 00 06 05 03 06 06 05 03 09 06 06 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 06 01 06 05 03 03 06 05 03 01 06 07 03 05 07 05 03 05 09 0c 06 0d 12 09 0d 04 06 0b 05 06 06 05 07 08 08 06 05 04 0a 0e 0a 0c 09 14 06 0c 0c 0e 11 10 0e 13 11 0f 10 12 10 0f 16 11 15 0f 0f 0f 12 14 15 21 12 18 1a 14 26 17 20 19 1f 28 25 2a 2b 32 2e 3f 41 3b 43 49 49 46 52 57 63 6b 6b 80 98 ad c2 de d4 dc db d4 e5 e0 db b8 92 8b 96 a5 b3 d3 d8 d8 d3 c8 c5 bd c2 cc cc d6 d6 df e1 d7 ce ad 8f 75 8d b1 bf c9 c6 c2 cb d1 ce c7 c4 b6 b1 ae ab ad a1 9f ae b0 ba b0 a7 aa a1 a8 a6 9a 8b 7c 80 7a 78 71 70 79 79 71 7b 7b 81 80 86 84 86 84 86 8d 92 92 88 7f 78 7b 7e 73 64 6f 5b 55 5c 4d 54 4a 44 3c 40 38 3d 3d 2c 2c 2b 22 22 29 1a 17 1a 17 23 1f 1b 0e 0f 0f 0d 0b 0e 10 0e 13 13 0e 16 0c 10 0f 07 0c 0a 04 06 06 04 03 06 05 0f 00 06 0f 03 08 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 04 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 05 04 00 06 05 03 04 06 05 03 00 06 05 08 00 06 05 03 01 06 05 05 04 06 06 07 0b 09 07 09 06 0d 05 05 06 06 07 0a 03 06 08 09 04 07 05 06 0b 06 0b 0b 05 0c 0e
 15 10 0d 1d 15 10 11 12 17 1b 0e 1d 0a 11 13 15 12 0e 1a 1c 19 13 22 23 20 1a 25 27 30 2f 35 39 42 45 4e 4f 4d 53 4a 5b 64 6c 80 84 8f 9b a6 c2 dc fb ff ff ff ff ff ff ff ff ff cb aa 8c 94 a6 c3 d0 de df d6 d3 ce c4 cd cb de df e2 e3 db d9 c7 bc b7 bf c0 bd c0 c8 d1 dc de e4 df cd c1 b8 b2 aa ae ad a6 a4 b8 c2 c0 ce c9 cd c0 c9 c0 ac 9b 97 8d 89 80 88 8a 8f 8e 8d 93 92 91 94 94 9e 9c a2 a5 a9 a9 a6 a0 8e 82 83 81 80 6f 70 72 62 67 65 65 66 5b 57 49 50 48 4b 43 40 37 32 2e 34 23 23 1b 16 24 31 1a 14 11 11 14 11 05 0f 0c 18 16 15 15 10 0f 0e 09 0d 0a 07 0e 06 0c 00 06 0c 03 00 06 05 06 02 06 08 04 02 06 05 03 03 06 05 05 00 06 05 03 01 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 03 00 06 05 04 0b 08 06 03 00 06 09 03 0d 06 08 09 0a 11 0b 0c 0a 0c 10 10 0c 06 08 08 0a 06 05 0d 09 06 05 08 0a 08 0b 0e 0f 0f 14 0e 0d 14 13 0c 18 15 0e 13 16 10 17 13 1b 14 16 12 12 17 17 1e 19 18 2a 1e 22 1f 2a 2f 29 30 3d 43 56 55 55 66 67 6d 6f 61 67 7a 8a aa b0 bf d2 e3 e8 fd ff ff ff ff ff ff ff ff ff ff ff f9 d5 c0 bb b7 bd d2 d2 e1 e4 e9 f2 e2 d4 d1 d3 d3 d4 d9 d5 cc cf cd d3 ca cd d4 d7 dd e0 e2 e7 f6 f4 e6 d5 bc b8 ae ad b6 a8 ad aa c3 d7 db e0 e2 e4 df da c9 bb ae a9 a1 97 92 98 9b 9c 99 9e a1 a8 a9 a8 a5 ab a9 ac aa ad a5 99 94 84 88 8e 8f 84 7d 75 77 76 6b 68 72 75 77 74 75 6c 6d 67 5e 54 52 4f 4b 3f 46 3f 33 3c 2f 29 28 20 22 20 18 1b 1c 10 18 14 11 0c 17 13 0a 14 0c 12 09 0c 0c 0c 05 04 06 09 05 02 06 05 03 05 07 05 05 07 06 05 03 00 06 05 03 04 06 05 03 07 06 05 04 06 06 05 03 02 06 07 03 02 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 07 03 07 0d 0c 0d 04 06 05 03 09 09 08 05 0e 0d 05 05 12 0a 0a 0c 06 0a 0a 0f 0b 0a 08 04 04 10 05 05 0f 06 0e 10 14 15 16 15 0c 13 1a 17 1a 14 1b 1b 1b 0f 23 14 1b 19 1b 1c 1b 20 19 1f 1f 29 25 30 36 3d 36 4d 49 50 62 64 69 76 84 83 7d 80 74 76 7d 92 b4 d0 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f3 ec ec ed ee ec ee e3 e9 ee ee ed eb e0 cc cb c7 cb d3 d0 d4 d3 d3 d9 e5 ed f0 f6 ea e2 ec f3 fe fc e5 d2 c9 bc b1 ad c1 be b3 cb d2 df d7 e3 e0 db d7 ca b6 a7 a1 a4 99 9d a1 99 9a a5 ab a6 a6 ad af b3 a9 b5 ae af af ab a1 98 8a 84 87 8e 95 88 8b 8b 85 7e 77 7e 7b 8a 84 8f 94 9a 92 92 8b 7b 65 55 51 5f 54 52 55 4d 45 2f 36 37 35 2f 2b 21 21 1e 15 17 1a 17 10 12 13 15 0e 17 0d 0b 06 0a 0b 05 06 08 05 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 05 08 06 05 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 09 06 05 0b 0f 06 05 03 09 06 08 09 00 06 08 04 08 07 09 06 0e 09 05 07 09 0c 0c 04 0e 06 07 0e 0f 0b 0b 10 11 06 0d 0c 0d 0a 19 1c 1b 1b 15
 1b 11 15 14 11 15 1c 19 11 1d 1c 15 1d 21 20 27 22 34 30 3c 51 46 55 53 58 5e 63 6c 7c 82 8a 96 99 95 8c 89 7d 83 90 a1 bb e0 fc ff ff ff ff ff ff ff ff ff ff ff ff e6 d8 d9 ee fd ff ff ff ff ff ff ff ff fa ff ff e8 d9 d0 cd cd cc d6 c6 dc de e8 f1 ff f6 ef ed e9 f3 ff ff f7 e1 d3 c6 b2 bc bd cb da cc d5 cf d4 c5 c3 ba c2 b5 ab 9c 8b 8a 8f 8f 95 91 96 92 9c a5 a2 ab ac aa b3 b2 b5 b0 a6 a6 a1 94 91 7f 89 90 94 9e 97 92 96 92 93 8e 81 91 92 97 a1 b6 b6 c1 c0 b6 ab 8b 7e 67 67 5c 5c 57 59 54 4a 40 47 4a 47 3e 32 22 21 17 23 1d 19 1f 18 11 14 0c 0b 09 08 0d 05 05 0c 09 07 03 05 07 05 03 00 06 05 03 02 06 05 03 00 06 05 07 00 06 05 03 05 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 11 0d 06 05 08 03 11 0c 09 0a 0b 06 03 0a 06 05 0c 0f 06 05 08 0f 0a 06 0c 0f 07 05 08 06 06 07 05 0c 06 05 03 0c 0c 0f 0f 0f 16 18 0b 1b 19 1b 17 10 19 1f 1a 15 19 1b 17 1e 29 1e 2f 23 30 35 4d 4c 51 4f 5f 5d 66 65 69 6f 6e 85 86 90 98 a4 ac a8 a7 a2 9e 9e 9e 96 a0 a6 bc be c0 c9 ca d2 d4 ca cd ca c4 c2 bd b4 c1 dc ee ff ff ff ff ff ff ff ff ff ff ff ff ff e1 d1 ce cb d5 dd db e2 ef f8 ff ff f7 f2 f2 f2 ff ff fa ef d9 c6 c3 c0 c8 cd de d1 c7 c5 bc b5 b0 a7 a3 a5 97 96 93 84 80 8b 91 98 9b 97 a3 a4 a9 b1 a4 a9 ad ae b6 b0 b3 aa 9a a3 9e 92 8e 8b 95 9a a4 a8 a2 a1 aa 99 a3 a0 a1 a7 a3 af be cf da d6 d6 c1 a3 97 7c 6f 6e 5f 63 6b 61 5b 50 58 6a 61 4b 40 2b 2d 21 26 23 1f 20 1e 11 1a 08 11 0f 0a 0b 06 03 00 07 05 08 02 08 08 05 00 06 05 03 07 06 05 03 01 06 05 03 04 06 05 03 05 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 03 00 07 06 03 00 06 05 03 05 06 05 08 07 06 05 06 14 08 14 0c 0c 07 06 07 04 09 07 07 0b 06 06 0c 14 06 07 11 09 0c 06 08 02 0d 0e 0d 10 10 05 05 07 0c 0f 18 11 16 16 1c 19 1a 19 22 21 1c 1e 1b 1e 27 1e 21 2b 33 34 3c 4e 53 65 6f 72 6c 6b 6c 66 6f 70 6e 73 78 81 85 95 9e b5 c0 b6 b8 b4 a8 ad a3 a5 ac a8 ac a4 a3 a0 a0 9b ad af b1 ad ac aa ad ba c0 d0 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ed d8 d3 d0 d4 e7 e9 f3 ff ff ff ff ff ff ff ff ff ff ff f1 d8 ca b9 c1 c4 c6 d1 c4 af b5 ab ae aa a0 a1 a5 97 9b 8f 92 91 9a 98 9c 9f 9f a3 a9 ab a8 ae b8 b8 ba b3 b7 a7 ad aa a5 a1 9d 9c 95 97 a2 a9 aa aa a7 b5 be c1 b9 b9 bb b9 c5 d1 e5 e2 d6 c3 b4 9b 89 85 80 73 74 75 73 69 6e 76 75 84 7f 6d 5c 44 38 35 36 2c 33 24 20 18 14 11 0c 16 08 09 05 07 05 06 06 0a 00 0b 09 03 00 06 05 08 07 06 05 03 00 06 05 03 05 06 0c 03 07 06 0b 03 02 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 06 03 00 06 05 07 03 06 0a 0d 0e 0b 10 15 10 08 07 07 12 06 11 12 08 06 09 03 08 06 0e 0d 07 07 0c 0a 0f 06 0d 08 0c 10 0b 07 08 16 15 15 18 15 1c 1a 1b 23 23
 24 1f 23 24 22 23 26 25 2a 39 44 59 5f 5f 7e 84 8f 9c 96 7e 75 74 7a 81 80 75 86 83 95 9d a9 b0 c7 c9 ca bf b8 c1 ae b8 ae ad ad a6 9c 9f 98 a4 aa a7 af ab aa b0 b7 bd c7 d8 ec f3 ff ff ff ff ff ff ff ff ff ff ff ff f3 e3 d2 c7 cf e0 eb fc ff ff ff ff ff ff ff ff ff ff ff f8 dc c2 b9 bd bd c4 d0 c6 b3 af a4 ac ae aa 9c a5 9e 99 9c 9e 9c a0 98 9b 9c a3 a3 a7 ad a5 a8 b5 b8 b4 b2 ab a9 ab ac ab a3 a0 a8 a1 97 9f a8 ac b5 be be ce cf c8 c8 d2 da e1 f9 f7 ea da b6 a5 95 8f 81 88 83 80 7d 7b 7a 86 9e 9f a7 99 8b 78 69 5e 45 46 41 3a 32 25 1d 1f 12 14 16 0a 10 0f 07 06 06 05 0b 09 06 05 08 03 06 07 08 00 06 05 03 00 06 06 03 04 0a 05 03 00 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 09 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 04 0b 08 09 08 10 0b 13 13 0d 0e 08 12 14 06 07 0c 0e 11 05 08 0f 0b 0c 12 0b 06 0b 09 12 07 0f 05 12 06 0f 15 08 0d 14 12 14 13 24 25 20 26 25 21 1d 20 20 29 36 40 40 45 5b 5f 74 7c 82 8b 93 9f 9f 91 93 8a 8f 93 8d 93 8f 8e 97 a0 a9 b9 c0 cd d2 d6 d7 cd c2 bb b9 c4 b3 ad b7 ae a2 a6 aa ac a0 af b4 af bf be bd c6 d0 d3 d7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ec cb c6 cf db ea f7 ff ff ff ff ff ff ff ff ff ff ff f0 da c6 b6 bc bc c2 d1 c8 b3 b7 b1 b5 a9 ad ae ad ac a5 a2 9e a3 9d 9e a5 ac a3 a1 ab a8 ab b4 b5 b3 b0 b6 af b1 aa aa b2 b8 ad aa a9 a2 a0 a5 ae ba be c6 d4 d8 d0 da ed fe ff ff ff f7 d3 b4 a5 a0 98 97 97 93 8d 8b 86 88 99 ac c0 c0 b6 aa 98 89 75 60 71 61 5a 3a 2b 21 2a 20 1e 16 16 08 05 0b 0d 08 0f 0d 02 06 05 04 06 06 08 07 07 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 07 03 00 06 08 03 09 06 05 0d 09 06 10 0e 15 13 14 0f 16 17 11 0b 0d 08 12 13 0d 10 12 0e 08 0f 0d 14 0d 09 12 0c 0c 0d 15 11 18 0c 13 11 0e 15 22 18 20 25 26 23 2b 22 27 2e 2b 28 32 3e 41 4e 5b 65 7c 82 84 8f 8d 93 99 92 91 9d a1 a1 9c a8 a3 a6 a3 a9 ad b6 b9 c7 ce d6 dc e4 e1 d6 d4 cc cc ca c2 bc c0 b5 ae b0 b7 b8 b8 bb bb bb ba c3 c2 bf c6 cd d9 ea ff ff ff ff ff ff ff ff ff ff ff f7 eb d3 c4 ca d1 e4 f3 f2 ff fd fc f3 e8 e5 dc de e4 ec db cb d0 c4 b9 b3 b5 cd c5 bb b9 bb b5 b2 b5 b8 b0 b0 b0 ad ad b2 b0 a9 af a5 a2 aa b2 b8 b0 b4 b6 b3 b7 b4 bb bb bb b7 b5 c0 b4 b0 af b2 b2 b2 a8 b7 ba c8 ce d3 df f0 ff ff ff ff ff f1 d4 c0 af a7 a3 a6 a2 a1 97 94 8d 8f a9 c0 e7 f5 ea d4 b8 a0 9e 8b 90 75 6b 57 3d 2f 2f 2e 26 1f 11 13 16 0d 09 09 05 11 08 09 08 03 07 06 05 07 01 06 08 06 07 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 05 06 05 03 03 06 05 03 00 06 05 04 00 06 05 03 08 06 0d 0c 1a 13 14 0d 10 13 14 18 11 13 11 0e 10 0c 0a 08 0c 07 12 10 05 07 0c 0a 07 0c 13 0f 0d 15 0d 16 12 13 1b 20 20 29 23 28 26 28 25
 32 2f 3f 4d 52 54 66 76 8b a0 a4 9d 8a 96 8f 9f 9c 9d a7 aa ad b3 b7 b5 c2 b7 b6 b6 c1 c2 d7 de e2 e1 e7 e4 e0 e0 d9 de d9 d3 cc d0 b7 bb b9 ba c5 bd bf c3 ba c3 bf bd bb b8 c3 c5 d3 df f6 ff ff ff fb ff f8 ff ff ff f3 df d3 cb c5 c5 d1 d9 da e4 e7 e4 d5 d9 ca cd c8 d2 d0 ca c4 c2 b8 b5 b5 c8 d3 cb c1 b9 b5 c0 bf b7 ad b8 ae af ba ad ae b5 b6 b4 b0 b0 b2 b4 b9 b2 b2 b6 b5 b9 bb b9 b9 ba b7 bd b5 ba bb b9 b6 b3 b1 b4 b6 b6 ba bd c5 d4 f0 ff ff ff ff ff ed ca bc ae b6 aa ad a7 a5 9b 9a 98 a1 b5 d1 ea ff ff f0 cb a9 b1 a7 ac 98 84 6b 5b 41 4a 45 40 32 24 16 17 12 0f 19 1f 0e 03 0c 05 0a 06 06 05 03 02 06 05 04 00 06 05 03 00 06 05 03 02 09 05 03 01 06 05 03 00 06 05 03 00 06 05 03 06 06 06 03 05 06 05 05 03 06 05 08 00 06 05 04 01 06 06 05 10 0b 08 10 0d 14 16 1e 1f 14 1b 10 17 14 10 0b 0d 0c 0a 07 11 08 12 11 0b 0d 05 12 0b 0a 10 16 11 0e 16 0f 12 14 20 18 1f 26 27 2a 32 36 3b 40 4d 60 5f 62 63 79 8f ae bc b1 a6 92 8c 9b 9f a9 ae b6 bc c1 c2 c7 c6 cd c7 cd cb d4 e0 e5 e8 ed ef ea e8 e6 e9 e6 e2 e4 e0 d5 c9 b2 ab c4 c2 c2 c9 c1 be bf bd bc b3 c0 c0 c0 c5 c4 d0 d4 d7 d6 de e0 db e6 e0 f4 eb db cc cc c0 c7 c9 ca cc d5 d9 d8 d9 cd cf cc cd cb c9 c6 c6 c2 bd bc b6 b6 c4 cd c8 bf c0 c4 c3 c3 bc bb b8 b6 b3 b8 b1 ba b4 a7 b0 aa b5 b1 b0 bb bc b9 bb c1 be b6 bc b7 ba c3 b7 c0 b5 b7 b6 b9 b7 b1 bf b5 b9 b4 b9 c7 c0 da f2 f8 ff ff fa e0 ce bc b8 b5 b4 ad b0 a3 a2 a9 a8 aa bd ba c5 ca c7 c8 b2 ae b3 bb c4 c5 aa 85 79 68 6e 6a 66 4c 2f 1b 1a 1b 16 1b 26 1e 10 06 05 03 08 06 0a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 04 06 05 03 00 06 05 06 00 09 05 0c 09 06 07 07 02 06 09 10 15 17 1b 1a 16 1a 16 18 16 10 0f 1f 19 12 0b 12 11 06 09 17 19 12 10 0c 10 11 11 14 1a 16 13 13 20 22 27 22 20 1e 28 2d 33 4b 59 59 62 6e 68 6e 79 83 97 ac be bc b0 a5 a7 a5 b6 b6 bb c5 c8 d1 d4 d5 d8 da de df e5 e3 e4 f6 fa ff fb fc f8 ef ee f1 ed ee ed e4 e1 d3 d0 c9 cf cd ce c9 cb b8 b9 b9 bf b7 bc bb c5 bf c5 c7 bc d0 c5 c9 d2 cd d0 d9 d0 d0 cc c6 c6 c7 c9 c3 c6 d4 c5 cf cc d1 c9 c5 cb cc c6 cb ce c7 c2 b7 be bd d2 d5 c8 c5 bc cc c0 c5 ca c1 ba bd bd b8 ba b5 ba ae b7 b3 b9 ba b4 c0 c1 b1 c1 bf c3 bf c0 b8 bd bd bb bf c7 ba b7 be b6 bc c5 c5 be bd bf bb c7 c9 ce e5 f3 f1 db d2 cc c7 bb ad b2 ae bb a8 a5 aa ad ad b0 ae a7 a0 9b 94 97 99 a6 c4 e1 ea d6 bb a9 9b 9c 9b 87 61 39 2c 16 21 1b 15 1c 27 18 0d 05 03 07 06 11 05 00 06 05 0c 00 06 05 04 00 06 05 03 05 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 05 04 06 05 04 03 06 05 06 03 06 08 0a 0b 0d 06 03 06 0e 12 0d 14 1c 1d 1a 19 1c 1d 18 14 1b 17 18 12 14 0c 0c 0b 0f 10 12 19 10 0e 0b 13 11 18 08 15 25 23 17 23 1e 1b 2c 1f 2a 44 42 53 5c 5d
 70 72 75 71 7c 80 89 97 aa bc c9 bf b3 b0 b7 c4 c9 cb de e8 d7 e3 e4 e6 ef ee f0 f7 f7 fb ff ff ff ff ff fd f7 fa f5 f1 f3 e9 e8 e5 d7 d2 d1 c5 d0 cd c6 c4 c7 c1 bb b5 b4 bd bf c4 c0 c4 b9 c5 bd c4 cb c0 c8 c1 c9 d1 cd c8 ce c2 c5 bf c2 c5 d1 d4 cd c8 ca cb d1 c8 ce cd ca d0 cb c7 c7 c4 c9 d8 db d1 c6 c9 c7 c6 bf c5 be be b7 bd b6 bf bd bb c0 c3 bd b9 bd b9 bd bf b6 bd bd bc bb be b7 be be c6 c0 be c5 c3 bc c0 bf c6 c1 c9 c8 cc cf c3 d3 d2 d6 d9 de d6 cb c5 be c5 c1 c1 b8 c3 bb b2 b1 ae a4 a5 aa a2 9b 96 93 92 a1 9d a5 c4 df eb e5 e0 d0 d1 b0 8b 71 5b 40 2b 1f 1b 21 25 2a 25 17 11 05 03 0e 07 07 03 06 05 03 02 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 04 04 06 05 08 04 06 05 05 00 06 09 03 06 06 05 07 03 08 09 04 05 07 05 06 0c 12 13 1c 1d 14 20 20 1b 20 19 18 11 13 22 1a 12 18 0f 0c 12 14 1d 12 12 0c 0e 13 0e 0f 17 1d 1d 1a 1b 1f 1f 25 29 2b 3f 42 4c 61 72 70 6e 6d 7b 82 89 92 88 94 a0 ab b8 cc bd be bf bd cb d8 d9 dd ed f1 e7 f4 f7 f7 fc ff fd ff ff ff ff ff ff fe ff f9 ff f6 ed f6 e4 eb e3 df d3 cc d1 c2 c4 c5 c0 bc be bc b7 aa b9 b4 bd bb bb ba be c1 bd c6 c2 c7 c3 c6 ca b7 cb c4 c8 c5 be c5 c3 ca d0 cf cb cb cf d3 d3 d1 da d2 cf cd d0 c6 cb cd d9 d6 d0 c5 cb ca cc c9 c6 c6 c2 b5 b7 b9 b5 bb b7 bd c0 b9 bf bd b9 b7 be be b3 bb b3 b6 b5 c5 c1 c3 be c2 c4 bc bf be c0 c2 cb cf ce c7 d0 cd ce d2 d3 cc d2 d2 ca cc c8 c8 ca c7 c5 c4 b9 be b8 af b0 ad a7 a2 a5 a5 a1 99 98 a1 a4 a5 a1 ae d1 e8 e8 ea dc a2 80 77 71 56 44 25 1c 1f 1e 28 26 20 17 14 08 06 05 05 05 06 05 03 00 06 05 03 00 06 05 03 00 06 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0a 07 05 0c 0b 07 0a 05 07 0a 0d 03 06 0c 0c 11 0e 17 19 11 16 1c 1b 1d 1e 22 1b 1a 26 18 1f 1c 1b 18 1b 21 1b 19 14 1a 13 17 12 19 11 23 18 24 1a 27 28 28 26 2e 38 4b 59 67 7f 7a 7b 7b 69 72 81 8b 95 a1 ad a8 b4 c0 b9 ca c6 c8 cf d2 cf da e0 ea eb f2 f4 fa fd fb fb ff ff ff ff ff ff ff ff fe fd fa fc f7 f5 f5 ef e8 e1 d2 d6 d2 cb cf c8 c2 c2 bc c3 bc b8 b9 b2 b8 b6 b6 bb bd c2 c8 c5 bc c1 c8 c1 c2 cc c4 c7 c7 c0 c9 cd bf c7 cd cf d0 d0 d2 d0 cc d2 d6 d0 d1 dc d1 d3 ce c6 d5 de e7 d6 c9 cc cb cd ca b1 c3 c4 c0 c0 c1 b4 c1 b8 b4 b2 b6 b5 ba b5 b7 c0 b7 c0 b8 bd b7 b8 b8 c0 c7 c2 c5 be c3 c3 bc bb c0 c9 c7 cc cd cc d8 d6 d5 d2 d0 d1 d5 d6 d2 c8 c7 c4 cb c2 c8 c8 bd bf bf bc b7 b6 b3 b2 a9 ae a8 a9 a4 a4 9a a6 a2 b0 b6 d4 c7 b6 97 86 8b 85 79 67 47 32 1d 24 24 21 1e 12 0a 11 11 07 0a 07 06 05 03 01 06 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 09 0a 10 06 05 0b 06 0a 0e 08 0a 0b 06 09 10 0d 0e 13 16 10 17 19 1b 21 25 20 21 1e 1e 24 22 23 19 21 1d 1a 1d 1c 1a 1f 18 1a 1a 17 1d 18 20 1a 22 17 22 2d 37 2f 32 39 3e 59 6b 77 88 7f 72 7a 7b
 78 83 91 a9 c0 c3 c2 b7 c1 c8 ce d7 d6 e3 d2 e0 ec ed f5 f3 fb fe fc ff ff ff ff ff ff ff fe ff ff fc ff fc fc ff ff f3 fb f1 ed e6 de d9 d4 ca cb c3 c9 b9 c8 c0 c3 bf bb b6 b7 bb b6 bd c0 b8 c1 ba c3 c3 cc c2 c3 c0 c1 c5 cb ca c9 cd ca cd cb d5 d1 d1 cb d0 d1 d5 db d3 d7 d2 d4 d9 ce d2 d6 e0 e3 d7 ce ce d1 d0 cd d5 ca c5 b8 be b5 b3 b6 be bc bc b7 b4 be b9 c0 be bb be bf b8 b7 c5 c8 bc c3 bf c2 c0 c0 bf c1 bd c8 c1 ca d4 d0 d6 d4 d1 d0 ce d5 d4 d1 dc d2 cb cd cc ca c7 c7 c7 c7 c8 be c0 bf bf be bc b8 b4 b3 a9 ad a8 aa a5 a4 9e a8 b2 b8 a1 96 84 95 8a 85 78 61 49 36 22 21 17 16 07 0f 0b 0d 07 08 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 0b 05 0a 0b 0a 0c 03 07 12 14 0d 10 17 09 0f 18 19 18 13 1f 13 14 26 23 20 1c 21 20 21 21 24 20 1f 19 0c 1b 16 1f 23 1d 1b 19 21 1b 20 1f 24 2f 32 34 35 38 4c 52 5e 5e 6a 77 6d 72 75 7a 87 98 a5 bc d6 d0 d7 c7 c7 d0 d9 d7 e0 e5 ec e9 f2 f3 ee f3 f9 ff ff ff ff ff ff ff fd fa f6 ff fb f0 f9 f4 ff fa f6 fd fd ec e9 e4 e0 db d7 d2 d2 d1 c9 c0 c3 c3 b7 b3 c0 b1 b1 ba b2 ba b5 b7 c3 bd c1 c4 c2 c2 ca c8 c9 c9 c7 c6 c9 c7 ca d0 cf d4 d4 d8 d0 d1 ce d3 da da dc d6 da d5 d2 d3 de e6 e2 e0 d3 d1 db d3 d9 d2 c8 cb c0 c1 b9 b1 b6 be be bc bc be c0 b9 bf b7 bf c2 be c3 c1 c6 c6 c4 c8 c8 cd c2 c3 c2 c2 c2 c4 bd c1 c0 d2 d7 db ce d7 ce cf c6 d9 c9 cf c9 c2 c7 bc b9 c0 c5 c6 c1 ce c0 c5 c4 c2 c5 c6 bd ba b0 b1 aa b2 aa ac 9f a4 b4 af a5 93 91 88 7d 7f 7d 6e 59 4d 3b 27 23 15 0e 06 0a 07 05 08 05 06 05 03 01 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 05 05 0d 07 08 0a 0d 06 07 0b 14 0a 08 12 0f 12 10 10 17 0d 1c 0f 1c 1f 16 1c 1a 23 20 1e 24 1a 1d 2a 1c 20 22 22 2a 23 1e 1b 21 24 1f 1b 21 14 1c 28 25 2e 29 29 2f 40 48 55 65 67 61 5c 5d 71 75 77 8a 87 9e b2 bf ce d3 dd e2 dd d2 df dd e5 e3 e9 f0 f5 f7 f2 fc fa fa ff ff ff ff ff ff f9 ff f4 f5 f9 ff f8 f7 ff fe f5 f9 ff fb fb f2 ed e2 dd da d9 d3 d1 ca c3 ca ca c3 be be b4 bf b9 bc bb b5 b3 c1 b9 be c2 c8 c4 cb cb ca cc c0 c7 c6 d2 c7 d0 cc d0 cc d0 d2 d0 d5 d1 d2 d6 da d3 d4 d2 d4 de e2 ef e6 d6 d4 d6 d9 df dc d8 d2 d9 cb c2 b6 be b9 b8 b9 bc a8 bb b5 c1 c5 bb c2 c7 c4 c8 c1 c4 cf d1 cf c8 cc c4 c4 c1 ca c4 bc cf c9 c7 d4 d5 d8 cd d5 cd c7 c6 cd c4 c4 c5 c6 c6 c4 c0 be c5 bc be bf c5 c2 ca c6 bf c5 c1 b7 c0 b7 b9 b2 b4 b1 a7 aa b7 b2 a8 9b 90 81 81 73 81 7c 70 61 52 46 29 25 1b 14 0f 0b 06 0d 0b 12 05 03 01 06 08 03 00 06 05 03 00 06 05 03 01 06 05 04 00 06 05 03 00 06 05 09 04 07 09 0c 0d 15 06 09 02 10 0d 0f 16 15 17 10 19 1e 12 14 13 18 1f 25 23 22 2b 29 24 26 20 25 20 25 24 22 27 28 21 25 23 26 22 1f 21 21 21 25 36 36 3d 35 3c 3b 51 56 69 80 74 6b 69 68 75 80 8c 97 a8
 b9 c9 d6 e4 e8 ef ef e2 db db db f2 ec ec f9 f1 f5 f7 fa fb fe ff fd ff ff fe fb f8 fd f0 f8 fb f3 fc fb ff ff fc ff fe ff f6 f3 f1 e8 e2 e1 df d9 d3 d0 ce d3 cd bb bd c1 b5 b3 b5 b6 b6 b5 ba c3 c6 c7 c8 c7 c4 ca d0 c9 d0 cb cb cc c9 d4 c9 c7 d6 d4 d5 d8 d0 da cf db de db d9 d9 d4 e0 d8 e3 f3 e7 e1 d5 e0 dd e4 e6 dd d2 d4 cc cb c7 be b3 b4 b2 b5 bc b5 c1 be c0 c1 ca c3 cc c3 c5 d5 ce d0 d4 cf d6 d7 d2 c9 c8 cb cd ca cf d0 d3 d7 df d0 d3 d5 cb ce d0 cd d0 ba c6 cb c1 c7 c6 bf c3 c1 bd c1 c8 c9 c6 d0 c3 c8 bd b7 ba c4 b5 b7 b5 af b1 b5 ac b5 a1 96 8f 82 7e 73 76 79 74 69 59 48 35 24 23 12 0a 0e 0c 08 14 05 03 00 0d 05 03 01 06 05 03 00 06 0b 03 02 06 05 03 00 06 05 03 04 06 05 08 04 0c 10 13 0a 0f 0c 0c 14 0e 11 0c 10 0d 0f 17 12 1d 11 1e 1d 1a 1b 1a 1c 23 22 25 22 20 27 21 1d 23 22 22 26 2b 29 23 2a 2c 25 28 26 28 23 27 34 3a 3b 3c 44 5d 6b 73 7b 8e 82 78 77 77 80 85 9b a2 b6 d4 eb fa ff f9 fb f9 ed e3 e2 e8 f0 e9 ea ec f3 fb f1 f6 f5 f9 fd f8 f8 fd fe fe fa f1 f4 f2 f9 f4 fb fa fb ff ff ff ff fe f5 fb ed ed f0 e7 e4 dd d7 cf d1 c5 c8 cb c4 c2 bc bb be b5 bc b6 c1 c3 ba c0 c1 c9 c8 d5 d0 ce d1 cd cd cd c9 d0 ce d9 d3 d4 d1 d1 db db d3 d7 d6 db de d9 e0 d6 e2 e4 f5 ee e1 e1 e4 e6 eb e1 df dd dc ce c9 c5 c0 be be bb bd bd bc c0 c2 c6 bd ce cd c7 d0 cf d4 d4 da e0 db e1 da d9 d7 ce d8 cf cb d0 d3 d2 d0 d4 d1 d3 d4 cd cf d1 cb d0 bd c3 b9 bd c5 c3 c3 be bb c3 bb ba ca c5 c9 c4 c4 c7 c6 bf bb c7 bd af af a6 b1 ba ad a2 99 92 86 86 77 71 7d 87 76 6a 55 3c 2e 1f 17 17 0e 10 03 07 0a 03 06 07 05 05 00 0a 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 06 07 0a 11 0d 0a 09 13 0b 11 16 18 11 14 11 15 12 14 1c 18 16 23 22 23 25 20 25 27 29 23 24 27 21 23 18 27 27 29 2f 27 23 30 32 25 30 2b 33 30 2b 2d 3a 44 55 71 85 8c 91 92 92 94 80 8f 89 8e 95 9e ae c9 e5 f6 ff ff ff ff ff f5 e8 ec f0 ed ec f2 f2 f5 f7 f1 f6 f2 f7 f9 fa f9 ff f7 ff f9 fb f1 f5 f8 f1 f9 fb ff fe fe ff ff ff ff fa f7 f4 f0 f2 e6 e6 dd e0 d2 d5 d0 d1 c2 c3 c3 c4 c6 bd b7 c6 c5 bc ba cb c8 cd d1 ce cf ca cd cc d0 cb d1 cd ce cd d3 dc c9 d2 d6 d1 d4 d1 db d3 de d3 dd e3 d6 f3 f7 ef ea e2 e4 f6 e4 ea e9 e4 e0 d9 d2 c8 cb c6 bb c1 c1 bf c2 c1 c6 c5 c8 cf d0 d3 da da d8 d8 d8 dc d8 db de de dc d6 d5 da dc d5 d4 d4 da da d4 d2 da c4 d0 ce cd ce cd c2 c6 c7 c9 bf c4 c2 b6 c0 c1 bb c8 cd c9 c7 c9 ca ca c1 c2 ba b5 b9 ab af ae bc b7 a5 a2 95 8e 88 7f 73 79 7b 87 88 78 5b 45 2a 27 1b 15 0c 08 06 06 03 01 08 05 06 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 08 16 10 0d 0e 0e 11 12 12 14 1a 13 1b 17 19 1c 1b 1d 21 20 22 23 2c 25 2c 26 2a 29 27 2b 20 24 19 2d 2e 2e 33 25 2d 2f 2c 34 2e 2f 31 32 31 41 43 69 7e 96 ab a5 99 9a 99 a5 a2 ae 9e af b1 af c6 db
 e3 fb ff ff ff ff ff f0 ef f9 f2 ec f2 ed f4 f4 f9 fd f3 f8 ee f3 ff ff f7 f5 f8 fa fd f9 fd f7 ff fd fc ff ff ff ff ff ff ff f9 fe f4 fe f5 f1 e6 e5 e0 dc d9 d7 d4 ce ce cb c6 c4 c4 cb bc c0 c3 cf cf d5 d8 d5 db d6 d3 d5 d5 d2 d4 cd ce d4 d5 da d5 d4 d9 da d6 de d7 df e0 da da db de e5 f0 fc f9 ef e5 eb f3 ee eb f4 ed e7 d8 d2 c9 c8 c1 c9 ba c2 c9 c4 c2 c6 d1 d0 d4 d7 cf da dc e9 dd e9 e9 e1 ea e8 e7 e5 e3 da d9 d8 e0 de d8 d8 db d6 cf d4 d7 d4 d0 d0 ce d0 cd c5 cc c9 c7 c6 bc c0 ca c5 c7 ca cd c5 d1 c6 c8 c2 c0 c2 bf bb b7 af a8 b2 b6 b3 ad a2 93 8f 88 85 77 73 77 84 95 8e 70 55 42 2e 29 14 10 10 06 0c 03 0d 06 09 03 03 06 09 03 06 06 05 03 00 06 05 03 00 06 05 08 00 06 05 0a 0b 06 0e 10 0d 10 05 11 13 11 17 18 19 1b 1a 1c 1b 29 17 25 26 20 25 25 2c 2a 26 2c 22 2c 23 27 26 25 27 23 2d 2b 2c 2e 31 31 2e 35 33 35 3a 3f 4d 66 82 ad b7 c7 c2 9c 9f 9d af b1 c0 c2 c4 c2 ca d8 e0 f6 fb ff ff ff ff fb f4 f3 e9 e7 ee ee f1 f4 f2 f4 f0 fa f4 f6 ff f5 f9 ff f7 fb fa fa f5 fb fc fa fe ff ff ff ff ff ff ff fb ff fe fb fc ed f4 eb ea e1 e2 da db d5 cc ce cf c0 c7 c4 c5 cd c7 c4 d1 cb d5 da d1 da d7 db d1 d6 d0 d2 d6 d7 d6 d0 d2 d7 d9 da d8 d7 d5 d3 df d7 dc e2 e2 e2 de f6 ff fa ef eb f4 f4 f4 fa fb fa e7 dd d6 d3 cb cc c7 c4 c3 ca c9 d5 d5 d4 d2 da e1 d8 e3 e6 eb e9 f1 eb e8 f0 e9 ea ea ee e5 e4 e6 e8 e0 de d7 e8 db d5 d7 d2 d4 d9 d1 d5 ce cf cb c7 c9 ce c6 c6 c7 ca cc c2 c3 c7 ca c9 c4 cd c3 c0 b9 b9 b9 b3 ad ad a8 b6 b3 b6 a8 9e 8e 86 7d 7c 77 71 7e 9a 9f 92 75 53 34 26 24 1a 13 0f 0e 08 09 06 09 05 03 06 05 07 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 09 0d 13 18 0c 17 10 10 13 19 15 1b 20 1b 20 1d 12 1d 22 23 23 26 2e 28 21 26 2c 23 2d 29 27 2b 27 23 27 23 1f 2b 22 2b 26 35 34 36 36 3c 4a 45 50 69 7f a4 c4 d5 da c3 a9 9d b1 c0 c6 ce d2 e4 e7 ef fa f9 ff ff ff ff fc fe f6 ee e8 fb ec ed f2 ea ec f8 f7 f3 fb f4 f4 f9 fd f6 fa f5 ef f7 fd fb fb ff fc fe ff ff ff ff ff ff ff ff ff ff fe fc fa f2 ef ef e0 e7 db dd d8 cc c1 cf c8 cc ca c6 cb c3 ce cc d6 d7 d9 d6 e2 dc e0 de d8 de d4 d8 d1 d4 d8 dd d6 d2 d6 da d3 dd dd d8 e1 dc e1 e0 e5 f2 fb ff f0 f7 f2 f6 fc fd ff ff f6 ed db d6 d2 c9 bf cf ca c9 cc ce cf dc dd df e3 e3 e7 ed ea ed ee ed f0 e4 eb f6 f2 f0 ea ea ea e2 e4 e9 e5 eb ea e1 de d8 d6 dd e0 d8 d4 d3 cd d4 c4 c3 ca cb ce c8 d2 d0 bc c6 bd ca c8 bd c0 c8 c0 ba bd b9 b9 b4 ac aa b0 b1 a9 aa 99 92 90 87 7b 77 76 7c 9c a0 a7 92 68 51 37 2b 1d 10 0c 0d 08 10 06 05 03 02 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 0f 15 0e 12 18 18 19 14 16 19 1e 1e 1d 1b 24 24 1c 19 24 28 23 2d 2c 25 26 2f 25 2f 2c 2d 27 31 2e 29 2c 24 28 2d 2e 2b 2b 33 35 44 44 4e 54 63 66 89 a6 ca dc ee e7 cc b9 af c0 cd d0 e0 ed f2 fc ff ff ff
 ff ff ff ff fc f9 f1 ea f3 ef f2 f4 f1 fc fd f9 ff f3 f4 fc f6 f8 f9 f9 f5 fb fb ff ff fc ff ff ff ff ff ff e9 ff ff ff ff ff ff ff ff ff ff ff fa f2 eb e4 e0 e0 e0 d8 d3 cf d7 ce cb d0 cc ce c9 d0 d3 da d4 db de e5 e0 de e1 d8 db dc d6 d0 d7 d5 d6 d8 d8 d9 e1 e1 d8 dd e1 dc e5 e0 ea f4 ff ff fb f1 f1 fe fb ff fb fb f3 e6 e0 d9 d6 cf ce d0 d0 ce cd d2 dd d7 dc e7 f8 f7 ef f7 ea ed f7 f5 ef f0 f8 f6 f3 f7 f3 f5 ef ef ea e9 f0 e5 e6 e6 de dd e4 de df e0 e4 df d1 d6 cc d2 d4 da d5 cf ca cd c7 c7 c7 be c1 bc c8 cb cd d6 c1 c4 bc bc af b3 b0 ab b0 ae a5 93 94 83 85 84 78 80 8f 9f ac ac 90 62 3e 32 2b 1e 13 09 0b 0d 06 0b 03 0a 06 05 03 05 06 05 03 05 06 05 03 00 06 05 03 00 06 05 13 0e 18 13 15 19 18 15 17 14 21 1c 1e 1c 23 24 1e 22 28 24 29 2c 28 2a 2a 2a 2f 2c 2d 27 2a 25 29 2b 2d 2c 34 34 2a 33 32 3e 3f 4b 54 59 6d 82 98 b2 d2 ed fc f5 e8 cd c6 c7 cc de e7 eb f3 ff ff ff ff ff ff ff ff ff ff f1 ea ee f3 fa f8 f9 f8 fa f9 fc fe f8 f8 ff f8 fe f1 f2 f5 f9 ff fc f8 ff ff fa ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f2 f7 e8 eb e0 d9 e0 db d6 d9 d4 cf d2 d3 cf d8 dd da d7 d7 da e8 e4 e4 e5 e8 e1 db db d6 cd d7 d6 cf dd db da e0 de df e1 db ed e7 ea f0 f0 ff ff f9 f2 f3 fb fa fd ff f6 e6 ea da d4 d5 d3 d1 da ce d7 d2 d7 e6 e1 f7 ec fb fe f8 f9 f3 fc f8 fc fa f5 f5 f6 f9 fe fd fa fb fa ec f1 ef e9 ed e5 e6 e3 e9 e2 e7 e4 e6 e1 e0 d2 d7 d3 d4 d5 d0 d0 d0 c5 c2 bf c0 c1 c2 c1 c3 c7 c4 ca bb c8 b7 bb b1 b5 ad ab aa b1 9e 98 99 8e 89 80 82 85 88 93 a1 b9 a4 7f 55 44 34 21 1a 05 03 0f 06 09 08 00 06 05 03 05 06 08 03 01 06 05 03 00 06 05 03 00 06 05 0e 17 19 18 16 1b 15 14 18 1f 13 1b 21 19 1b 26 29 25 28 24 2a 29 2a 28 37 2a 2a 2e 26 2c 2f 34 2d 30 26 30 28 2e 2f 31 3d 4b 51 55 5c 77 94 ae c5 e2 fc ff ff f6 eb d8 d2 d5 de e5 f6 ff ff ff ff ff ff ff ff ff ff ff fb ea e5 e7 eb ed ef f9 fc fe ff ff ff ff ff f9 f4 fa f9 f8 fd fd ff f8 fe ff ff fd ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fd f0 e9 e8 e8 e4 e1 df d4 da d9 d8 d6 da d7 d5 dd db e0 d6 dd df e9 e4 e9 de e7 e1 d5 d5 d0 d2 d5 d6 e0 e6 dd e3 e8 e5 e9 e7 eb f1 f6 f3 ff ff f8 f8 f2 fd fa fc fb f8 f3 e7 e4 e0 d4 da ce d8 d9 de de e3 e4 e8 fa f8 ff ff ff ff ff fd fb f9 f1 f7 fa ff ff ff fc ff f8 fb fe ef f5 f2 ec e8 ed e9 ea ea eb eb de e3 e3 d9 d9 de d9 da d7 cc cb c6 c8 c4 c5 c1 ba c8 c2 be be ba bd c0 b7 b6 aa a1 aa a3 b7 af ac 9d 97 8f 88 8a 89 82 85 80 8a aa ab 90 76 4e 3c 2b 27 11 13 0a 09 05 04 00 06 05 03 00 06 05 03 06 06 05 03 05 06 05 03 00 06 05 12 19 15 1a 18 1a 19 1c 16 26 1d 24 27 22 21 1c 1c 21 2e 2b 30 34 29 36 2a 35 28 32 30 2b 2d 2b 30 2b 30 35 36 3a 39 3d 4e 4a 5a 67 88 a6 c9 dd fa ff ff ff ff f3 e7 e0 e2 df ea f1 fa ff ff ff ff ff ff ff
 ff ff ff ff fc e7 d8 e1 e8 f1 f5 fc ff ff ff ff ff f6 fc fe f4 f6 f4 f7 f9 fa ff ff ff ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff fa ff f5 ed ef f0 e4 e1 e4 da e1 de d9 da d2 d7 d5 d8 d8 d9 de e2 ea e8 e7 ea eb e9 e2 d4 dc d2 d6 e4 db e1 e2 e2 e8 e5 ec f0 ee ee f1 fc ff ff ff fd f2 f1 f8 fd ff fe fb ec ed e3 e0 dd d9 df e0 de e3 e4 eb ec f1 ff ff ff ff ff ff ff ff fd ff fd fd ff ff ff ff ff ff ff f7 ff fa fc f7 f8 f2 f5 f1 f0 f0 ec ed ee e5 e6 e2 dc dd da d8 d5 cd ce cf c0 c5 c1 c6 bb c3 c4 ba bb b8 bb b3 ac ac 98 9e 9f a3 ae b3 a5 9b a3 95 95 8d 8b 87 8a 86 8b 9c ba b3 8e 6b 4a 33 1e 1a 11 13 07 05 03 06 06 0c 03 02 06 05 03 04 06 05 03 00 06 05 03 00 06 05 14 17 1a 16 19 17 11 23 1c 1f 23 25 1c 24 2a 25 23 26 34 24 32 27 26 35 2b 39 34 36 39 36 35 2b 2b 27 32 33 34 33 49 44 53 5c 63 7c a8 d4 f0 ff ff ff ff ff f9 f4 f0 f4 e6 e8 e9 ff ff ff ff ff ff ff ff ff ff ff ff ff f0 d7 d1 d5 de eb ed eb ff ff ff ff f7 fc fe fb ff fb fb fa ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f8 f8 ee f0 eb e4 e2 e3 de db dd dd dc db d4 d7 d3 d3 d8 de dc ef eb eb eb e5 e7 e0 e0 d7 df dd df e3 e3 e4 e1 e1 e9 ee f3 f3 f4 f9 fd ff ff f9 f3 f8 fa fd ff ff fa e7 ee e7 df e6 dc e4 e6 e5 e3 e6 ea f4 ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff fd f4 fc ff fe f8 f2 f5 f9 f2 f3 ee f3 f2 e8 e9 e4 df de de d7 d6 d1 c9 c2 c7 c0 c4 c7 c2 c0 b5 b8 bc be ba b0 a6 9e a7 9f 9e ae a9 a8 a1 a3 98 98 95 93 8d 89 84 82 87 a5 b5 a1 87 65 49 35 24 14 15 0d 08 09 06 0e 05 03 05 06 05 03 06 06 05 03 00 06 05 03 00 06 05 0e 0c 1e 20 1f 1f 1d 1c 22 24 22 27 1f 2c 1e 26 2a 21 2a 24 2b 2b 2c 37 30 2f 2e 2b 32 2b 30 37 25 30 32 40 3b 42 42 46 58 5f 76 8f c4 e0 f9 ff ff ff ff ff ff ff ff f8 fe f2 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff e3 cc c6 c6 dd e0 e7 f2 f6 ff ff ff ff fe ff f9 fe ff ff fa fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f0 f8 f1 eb f1 ed e9 e0 de db dc e2 d8 d9 dc d5 d5 d4 d2 da e1 e4 ee ee eb e7 df e6 dd dc e9 e5 e7 ea ed ec e8 e8 ef ed f1 e9 fc f6 ef fb f5 ec f1 ea f9 ff ff ff f9 f0 ed e4 eb e9 e1 e3 e1 e4 ed ec f4 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff fc f6 f5 ee f8 f4 f0 f0 e8 eb e5 e0 e4 db df d9 d5 d1 d2 cc c5 cc cd c3 c9 c7 ba b6 b6 c1 b1 a5 ab a4 9e 99 99 9d a6 a5 a2 9f 97 8e 8e 91 88 86 84 79 89 8e b5 b8 9e 7b 59 43 2b 23 18 10 13 0e 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 1b 19 1c 21 20 22 1b 26 22 23 24 25 2f 1f 2a 2d 2f 20 36 24 2f 2f 2e 35 33 28 38 37 32 34 38 36 34 31 39 39 3d 44 4d 52 65 72 86 b3 d8 e6 e9 eb f6 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff
 ff ff ff e6 d4 cc c4 ce d5 e1 e7 eb f9 f9 ff ff ff fe ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f0 f1 f2 f2 e8 ea e5 df e3 e0 e3 da e1 dc d7 d2 d8 de e2 ee e9 ed f2 f2 eb eb ed ea e4 e2 ee f2 f6 fc f6 f6 f2 f5 f5 f3 fa f6 f8 f1 ef f2 eb f7 f1 ff ff ff fe fb e5 ef e8 e6 f0 eb ed ed f0 f0 f2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fa f4 fb fe f6 f5 e7 ec e4 e8 e3 e6 e6 e4 dd d4 d5 c9 c5 cd d0 d2 d2 c8 bd ba c1 ba b1 b7 af a9 a8 9f 9d 9a 97 a1 a2 95 93 96 86 8a 8c 88 85 88 88 96 a8 be ab 8e 6a 54 46 24 21 1f 16 05 09 06 05 03 06 06 09 04 04 06 05 03 00 06 05 03 00 06 05 16 0f 14 1f 17 21 24 1e 2a 2a 1e 23 24 25 29 26 26 2f 34 26 29 35 26 32 32 37 30 35 38 2a 37 37 38 34 3b 3e 42 43 54 67 7c 86 a3 cc da d5 d1 de e6 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ee d4 c6 c8 cb ca ce d0 da e4 e6 f1 ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 f1 e8 eb e8 eb ef e4 e0 e6 da dd d7 d9 d9 d4 df e2 e8 f6 f8 f5 f7 f2 f0 f3 f2 f6 f8 ff ff ff ff ff ff ff ff ff ff fb fa f8 f5 f1 f5 f4 fb ff ff ff ff ff ff fa ee f2 e7 ee f5 f0 f5 ff f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fe ff fb f9 f6 f3 f2 ef e5 ea f0 e5 ee ea e1 e2 d4 d6 d0 d8 d3 ce d1 d0 d0 d2 c5 c4 c6 b6 b3 b6 a8 ad 9e 9e a4 9b 9f 94 96 9a 8f 91 8b 89 89 86 87 93 98 a4 af b8 a3 7c 63 4d 3f 2f 1b 07 03 02 06 05 07 00 06 05 07 0e 06 05 03 01 06 05 03 00 06 05 19 1f 1d 1b 1b 21 21 22 1a 21 21 26 29 28 28 2c 28 2f 2d 29 26 2d 2d 35 2a 2f 2d 2e 33 33 2f 38 3a 3b 35 3e 43 45 5b 6f 88 a0 c1 d9 cd bd c0 ce df ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 db de d6 d0 ca c2 c2 cb c3 d0 d1 ce de de e4 ef f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 ef ef e7 ea ea e3 e6 e3 d8 e1 d7 d5 d6 db de e5 ed f3 f5 f2 f8 f8 fd fd ff ff ff ab ff ff ff ff ff ff ff ff ff ff ff f2 fd f8 f0 fb ff ff ff ff ff ff ff f8 fa ec f3 f0 f9 f7 fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fd f9 f5 fa f0 ef ec ee ea ee e2 eb df e1 d7 d3 d4 d5 d6 d1 d5 d7 d4 d2 cd c9 be bc b6 b8 ab ab a0 a1 94 9f 98 9a 91 96 93 8d 85 87 8c 85 85 91 91 94 aa bd ab 92 74 54 41 36 28 18 11 02 06 05 03 00 06 05 03 08 06 08 03 00 06 05 03 00 06 05 1d 1f 1e 25 1e 29 1d 20 25 22 26 28 27 2b 2d 2c 2b 27 28 2e 2e 20 2c 36 30 31 35 34 33 32 39 36 39 42 43 41 48 52 65 7d 95 c1 d0 cd c5 b0 ba c4 c9 df e9 ff ff ff ff ff ff ff ff ff ff ff ff f0 e0 d8 d1 d2
 d1 d1 cd c5 d4 c8 c8 ca c9 d6 d9 dc ea ef f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f8 f9 f2 f0 f6 e7 e8 e1 e0 e5 e9 da e3 e7 e8 eb ef fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f4 f2 fc ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fc ff ff f6 f6 f6 f3 ee eb f2 f4 e0 e5 e3 df db df e1 d4 d8 da da d3 d0 d2 c1 c3 b4 b1 a4 a6 a4 9f 9a 94 95 94 95 98 8d 89 95 8a 90 8a 8e 90 90 a0 ac b6 b9 9c 7e 59 45 36 26 15 0e 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 24 1c 25 1f 2a 26 27 24 23 2e 28 2b 25 2c 32 31 25 29 30 28 2b 27 39 3d 35 34 2e 38 39 2c 33 34 3a 41 3e 4d 57 5d 77 92 b4 cb ce b5 a7 a3 a1 b2 b9 d1 d5 f3 f9 ff ff ff ff ff ff ff f0 e1 d9 d5 cf d5 c6 da d7 d2 cf cc d1 c7 ca c1 ce d0 d9 d6 e8 ed f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fa f4 ef f3 ef ed ea e8 ec f3 f8 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fd ff fd ed f1 f5 ec ef e8 f2 e6 e4 e5 e6 e0 e1 e7 e2 d6 de d9 d2 d1 c5 ba b8 b8 b5 b0 a7 a9 a0 9c 9b 9d 94 97 95 90 8e 93 90 99 8f 95 97 91 a0 b6 b4 a3 8a 69 50 35 26 14 11 0a 06 05 03 02 06 05 09 03 09 05 03 07 06 05 03 00 06 05 17 1d 22 17 1e 21 25 27 2b 28 29 20 2f 31 2d 37 2a 28 2d 20 2c 2d 27 34 26 33 36 32 31 33 36 3f 3a 45 47 44 58 6f 82 a2 c4 cf b5 a1 a1 a2 a1 a8 aa b8 bc c7 d8 d6 e5 e5 ec f5 e6 e8 db cc cc c7 d5 cf d2 d8 d5 d1 d9 da d6 cd cf cf cf c9 d5 dd e2 eb ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f3 fa f7 ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff ff fc f8 f6 f9 f7 f3 f7 f0 ef ef e9 f3 e9 e2 e0 e4 e3 f0 e0 db d9 cd cf c9 c4 bd bb b5 aa ae ac a9 a4 a8 99 99 9e 9a 99 92 9e 97 98 8f 98 93 99 9c a2 b2 a9 8e 78 55 41 21 20 0b 01 10 05 04 01 06 05 03 05 06 05 04 00 06 05 03 00 06 05 19 1d 24 20 23 23 1f 22 26 26 27 22 24 2b 29 2d 2e 32 2f 2a 2a 30 33 34 35 33 2f 2d 3f 39 36 38 3f 4a 47 4c 66 78 95 bb c1 ba a9 9f a7 99 a5 a5 a2 ac b7 b6 bf c7 d3 d8 d5 d7 ce d7 d1 ca bf b5 ce cc d7 dd
 e2 df db d9 e0 da d9 cd d5 d8 d5 eb e8 e2 f5 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 f7 f1 f9 f1 f0 f1 f4 f9 f2 f2 f4 ed ee e8 e2 e6 d9 df cb c7 cf ca c8 ba c1 b5 bb b4 af ab b0 a5 9e a3 9a 91 96 9a 94 9b 8e 99 92 9d 9d 98 af b3 a7 95 7b 5b 44 29 21 14 07 15 07 06 00 06 09 03 00 06 05 03 06 06 05 03 00 06 05 1e 1f 1b 29 20 25 27 24 22 2e 2a 2e 32 31 34 27 2f 2a 35 2e 2d 33 2d 33 30 33 33 3c 42 3c 3e 46 44 4f 50 51 65 7f a6 c8 bb ae a0 9a a1 9d 9f a8 a4 a7 b0 b8 bb c6 cd d1 d7 d7 d1 d5 d0 c8 cf d0 cc d0 d9 d1 db e0 da d7 e6 de dd e5 e6 d4 e6 e6 ea e7 f3 f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 f9 f0 f2 f0 f8 fa ee f6 f2 f2 ef e8 ee ef e8 e3 dc d9 cb d1 c8 cc cf ba be bd b4 b4 ad ae aa a8 a4 ad 97 9a 9a 95 93 a0 96 a2 93 90 9e a0 ae b6 99 81 69 55 3f 32 1b 0b 0d 09 11 06 09 05 06 0e 0b 05 03 00 06 05 03 00 06 05 1e 1f 1c 26 21 22 20 26 29 23 2d 30 2c 2b 34 37 2a 37 32 2c 29 33 27 2b 36 2e 34 36 3b 3a 38 45 47 48 54 64 76 8d b5 bc b0 99 9a 99 a3 a0 a4 a6 ab 9e a7 ae c1 cc cb c6 d1 d9 d6 d5 d2 cf cb d0 cc d9 da d9 e0 dc e1 e2 ea e9 e8 ec eb e5 e5 ed f2 f6 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f9 f9 f5 f8 f8 f9 f2 f8 fa f7 f3 ef eb e9 e2 e2 e2 dd df d6 d4 cb cd c4 c7 c4 ba b5 af ac ae a6 ac 9e 9d 99 9a a2 a4 9c 9a 9b 9f 92 93 a1 98 ac aa 9f 7c 5e 54 3f 35 27 1d 15 11 0b 0e 0e 05 07 03 07 0f 03 00 06 05 03 00 06 05 1b 20 2a 29 29 25 21 25 26 20 26 29 31 2a 27 31 22 2c 34 31 34 34 33 33 2d 35 34 39 3a 3b 46 45 4f 51 52 60 7b 9f c2 b4 a6 a2 9e 9f 99 a1 a6 a6 a5 ab a4 ae bf c7 ce ce c7 d3 d4 db d8 d9 d5 d4 d4 d4 df da
 e3 de e5 ed e9 ee ed f2 ea f3 f6 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fd f9 fa f8 f3 f7 fc f4 f8 f3 ef ed ef eb e6 e4 e0 d2 d7 d0 cb ce c8 be c4 c0 b3 b2 b3 a8 ac a7 a6 a4 a3 9e 9f a0 93 98 9c 9c 9a 95 a2 a3 af 9b 86 76 5d 4a 42 31 20 16 11 0c 02 0d 08 0c 10 06 06 06 00 06 05 03 00 06 05 1a 21 22 21 22 29 26 31 2f 2a 29 27 33 2d 31 2c 2a 2e 2f 33 35 35 34 3b 33 35 37 35 41 4c 4e 55 58 5c 5d 70 86 a0 b1 ac 9f 9e 97 a2 ab a6 a4 ab a6 aa a9 b0 b6 c8 cd c9 cb d8 d8 db d7 d7 d0 ce d2 d8 e0 e4 e2 e2 e7 f1 f4 f0 f5 fb fe fb f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f5 f9 f6 f9 f3 ef f1 ef f7 f0 f4 e9 e6 e3 e4 dd dc da d3 d3 d3 d3 c2 ca c1 c1 b7 b5 ad ac ab a4 9f a6 a6 a5 9f a0 97 a2 9b a1 93 9e aa 9e 9d 84 7b 71 5b 4e 40 2b 1a 17 13 14 08 15 09 09 0b 0b 08 03 06 05 03 01 06 05 21 1b 25 1f 24 27 20 26 22 2a 36 2e 32 2e 30 25 38 2a 31 31 2f 2c 29 32 33 36 30 3c 42 4b 54 5b 64 6a 73 7c 94 a0 a7 a5 a1 a1 9d a4 a6 ab aa a6 aa a9 ad ac b5 c5 c9 d4 d6 d0 d3 dd d3 d9 d9 da db d6 d8 db ed e2 ed eb f7 eb fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fd f2 fc f4 f3 f9 f9 f2 f1 f1 ea e5 e9 e8 e7 e4 de d9 d4 d2 d2 d1 ca c1 c2 b6 b5 b2 a8 a8 aa a8 a4 97 9e a3 a0 9c 9f 96 98 89 94 8d 92 8d 82 7f 79 63 54 44 35 27 1f 17 11 11 0d 17 0b 11 0c 05 0a 06 05 03 00 06 05 19 19 21 22 20 28 25 26 20 2c 2a 33 2d 25 2c 34 2a 2f 34 2e 2c 37 31 3c 32 3e 38 49 57 56 58 5d 59 64 77 87 8d 9c a3 a5 a8 ac ad ae a9 ab b2 b4 b4 ab ae b1 b2 b9 c4 cc da da e3 e0 e0 dc e4 dc d6 e0 e1 dc
 e3 e7 ee f2 ee fd f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f7 f4 f9 f4 f4 f7 fc f8 f3 ed f6 e8 ec e0 dd de da df d5 d6 d2 d5 d2 ca ba bb b8 b6 b8 b2 b0 ad aa aa a9 a4 a5 a0 a0 98 9e 94 8e 84 7d 75 7f 6d 70 75 6f 60 4d 39 2a 29 1b 15 0c 0b 09 05 06 0a 03 02 06 05 03 00 06 05 20 1d 21 24 1a 27 23 25 2d 2d 28 30 32 2d 33 2d 2b 32 38 31 35 35 31 3d 32 3e 3a 49 57 5a 64 58 61 5c 72 94 97 9c 9e 9e a3 a8 b2 b3 b1 ab af b4 bb b4 ad b0 b4 be c7 d3 d0 da dc e4 e3 e0 e4 e0 de e0 e6 e5 e7 eb f5 ec fe f8 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fe f4 f3 f7 f7 f2 f8 ec f3 ef f3 e5 eb e5 e7 e3 e2 e0 e2 d4 d2 d6 c6 cd c4 c5 b9 ab b9 b6 b9 b3 ad ac a6 a3 ab 9f 99 a1 99 8c 8d 85 78 73 6f 67 65 78 76 64 55 44 39 25 18 1d 09 07 03 06 0d 05 03 00 06 05 03 00 06 05 25 20 22 25 22 2a 24 1e 24 32 2b 31 30 2e 2f 2a 31 2c 30 2f 3f 31 34 3c 43 39 4b 58 5f 5d 63 64 5a 59 72 93 92 a0 a3 a3 a9 a8 b1 af b3 b7 b1 b3 b9 bb b5 b0 b1 b1 bc d1 d4 d7 e7 e2 e3 dd e2 e3 da dc e7 ea f1 ed f6 fc ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fe fa f8 f5 f5 fc f0 f8 f2 eb e9 e4 e3 e9 e0 e2 e2 d9 e1 d5 d2 d6 d0 ce cc bb c9 c6 b9 bb b2 b2 af af ae a6 ac 9e ab 9e 9a 95 8f 7f 75 76 71 71 64 6f 78 80 75 55 52 3f 33 24 14 0e 0d 07 05 06 05 03 00 06 05 03 00 06 05 1c 20 25 21 22 29 21 1c 21 30 26 31 32 29 31 33 2b 30 30 26 39 2f 38 40 44 4f 4d 57 60 6a 66 6b 60 6b 7c 8f 9b 96 9e 9b a3 ac b1 b7 b6 b5 b9 bd ba b2 ba bc b0 b9 c2 c5 d7 d0 e3 e1 e0 e2 de e4 e7 e3 e3 ec
 ec ef f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 fd f7 fa f6 f2 f7 ea ed ef ee e9 e7 e5 e5 e0 de dc d8 db de d1 d6 d1 cb c4 c9 c2 bb b6 b6 ae a9 ab aa a1 a6 aa a3 9f 9c 94 90 81 75 6f 6c 72 68 66 68 79 75 72 66 52 3e 2b 1a 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 20 25 2b 24 26 1f 28 23 25 2b 2d 33 2f 2d 2e 34 30 40 37 34 3b 38 45 48 56 56 5c 6a 64 6d 72 69 70 83 94 9a 9b 9f a5 9e a4 ae b6 b8 c0 bb b8 c0 be b9 bc c0 c1 c4 d0 d6 db e5 dc e4 e6 ec ea e9 e5 ee ed f2 f7 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff f9 f9 f5 f2 f7 ee f1 f0 eb e7 ed df e8 e1 e1 e3 d9 dd cd cf c9 ce c8 c8 c7 c1 ba b6 b3 b0 a8 ac a9 a1 a3 a8 a4 9f 94 90 83 7b 79 7b 6b 70 71 6b 68 75 7e 75 63 50 47 33 1e 15 0a 05 05 00 07 05 03 00 06 05 03 00 06 05 1b 1a 22 25 2b 20 21 23 29 2d 2b 34 29 2c 2a 35 2c 33 36 30 44 31 3b 48 4d 56 53 66 6d 71 76 74 6e 7d 83 9c 93 95 a3 a2 a2 a8 b0 af bf c1 bb c3 be c0 bc be be bd c7 c7 d3 db d8 df e7 ec eb f5 ea eb ee ee f9 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa fd f9 f4 f9 f5 f9 ee f1 f7 e8 e4 e8 e8 e7 dc db db d6 d7 d5 cf cc c5 c4 c1 be b9 bc ba aa b0 b0 ab ae ad 9e a3 a4 9c 8e 89 7e 79 6f 68 6e 6b 6b 5f 6a 69 73 78 65 55 47 3a 26 1c 09 08 03 07 06 05 03 00 06 05 03 00 06 05 1f 1c 25 25 1a 20 20 24 2c 26 2a 2c 30 30 35 2d 2d 39 34 33 3b 3a 3c 46 44 57 56 6c 6a 75 76 7b 7f 7e 8b 88 95 94 8d 95 a3 ac a8 b1 b8 b9 bf bf c9 c4 c7 c3 bc c4 c9 ca d7 d6 d8 e3 e9 e6 ec f3 f3 f2 f3 f5
 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fb f7 f5 f3 f5 f8 f0 f0 ed e5 e9 e2 e2 e8 e1 da d5 c9 cc cd c4 ca c3 c0 c1 b5 bb ad b0 b2 af aa 9f a9 a9 a4 99 a1 93 87 79 73 71 71 73 75 70 6e 62 55 5e 73 75 6a 56 4c 35 1f 19 09 05 06 01 06 05 03 00 06 05 03 00 06 05 1d 20 23 23 20 1f 1b 22 31 29 24 2e 31 2c 31 33 34 32 36 35 3c 3a 47 41 51 5f 5c 6b 73 74 87 85 83 84 89 89 91 92 8f 97 a1 a8 ab b2 ba bd c6 c4 ca ca c4 c7 c4 c2 c9 c5 d2 d7 d8 de e9 e5 ee f8 f3 fc ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fb f3 f6 f7 f6 f4 f5 e5 ea f0 e4 e8 e8 dc e1 d5 d8 d3 cd cc c8 c5 c4 be b9 bd b5 b0 b6 aa b2 a6 a1 af a3 a3 a0 a1 9d 89 84 79 73 74 75 6e 78 70 68 5d 57 5e 6d 73 6b 5d 46 35 22 1c 08 0c 03 09 06 05 03 04 06 05 03 00 06 05 1f 1c 22 24 1d 1e 23 1e 1f 30 2a 29 31 2f 2f 34 32 34 3b 37 34 45 3e 51 55 56 68 6c 76 77 88 84 88 88 84 8b 88 8d 90 8d 9a a1 a8 b0 bf c3 c8 c2 ca c8 c7 c5 cb cc d0 d6 d7 dc d5 db dc e1 e9 f5 f9 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe f9 f8 f7 f0 f6 ef f4 f5 f1 f8 e9 e1 e0 e4 d9 e0 d7 d3 cc d1 c6 c8 bf be ba be b3 b1 b1 a2 a7 ab a1 a7 ac a1 9c 97 8f 81 79 74 70 74 6e 6d 6c 71 6d 5d 59 60 6b 72 6c 60 52 39 2c 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1a 11 16 20 22 1a 25 1e 23 2c 2b 2b 2a 28 2a 2d 2a 2b 35 3c 3b 45 38 42 4a 6a 62 6e 7a 79 84 89 8b 8a 7d 84 85 82 8a 85 91 95 a0 b0 bb c1 c4 c8 c2 c4 cb c8 cb d1 ca d1 d5 dd de dd e0 e9 ed ef f1 f2 fe f9
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 fa f9 f7 fa f6 f1 f4 ef ec f0 e6 e5 e3 e0 e4 ce d4 cf d5 d0 c8 ca c4 ba bb be bf b9 b6 aa ae a9 a9 aa a9 a3 9b 98 98 8c 8a 7d 74 6e 67 64 6b 64 6e 6e 67 60 57 5c 62 75 6b 60 51 3e 2a 1e 0c 06 03 02 06 05 03 00 06 05 03 00 06 05 1d 15 23 1f 27 24 23 2b 2a 22 2a 28 2f 2e 2e 33 2a 32 32 33 35 3f 40 41 4d 61 64 74 73 86 86 8f 8d 8e 85 88 83 7b 80 89 8b 98 9f a6 b2 bb c4 c8 c7 ce c9 cb c2 d0 cb d2 d0 d6 db df e2 e5 e9 ee f2 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb fb f5 f6 f1 fa f5 f4 f8 f4 fb f0 f6 ef e9 e9 e3 e0 df db d9 dd ca cf ca c5 c6 be c2 c1 bc b5 b8 ba af a7 ab a4 a2 a4 a3 95 9d 92 94 80 79 6c 6f 63 68 66 66 70 74 62 57 58 51 67 78 70 61 4e 40 27 1b 0f 05 03 0a 06 05 03 00 06 05 03 00 06 05 1c 15 1f 1f 24 25 2a 27 21 2a 23 25 28 32 30 2f 31 2f 35 30 37 39 44 46 44 60 68 74 7b 7a 91 8f 8f 90 89 84 78 7e 82 7f 89 91 95 a5 ad b9 bd be c1 c6 c5 ce d2 ce d3 d4 d4 d8 e3 e3 e2 e6 ed ee ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 fc f5 f5 ee eb ed f2 f2 ef f0 f1 f1 ec e9 ea ea e6 d7 e1 d7 d4 d3 d6 d2 ca cf c0 c0 bd c1 b8 b8 b2 aa ad ab a4 a2 a0 a8 9f 9d 97 92 88 7d 78 70 70 67 62 68 6b 76 63 5d 55 55 5c 61 73 73 63 54 3f 2c 1b 0e 05 06 06 06 05 03 01 06 05 03 00 06 05 16 17 1b 1b 1d 27 1e 25 22 28 2c 2d 29 29 2b 2d 32 34 31 35 2c 34 39 3f 48 52 60 76 82 86 88 8d 8e 94 80 80 82 7e 7c 7b 87 86 8f 94 a4 af b7 b7 c3 c0 c4 ce d0 cc d4 d4 cc ce de da e1 e3 e7 f1 f9 f7 ff ff
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 f4 f1 f4 f4 ed ed f1 ed ef eb eb ee ea e9 e4 e0 e2 d9 d3 d3 d8 d7 cc ce cb c6 c9 b8 c2 b7 b8 af b2 b5 a9 ac a0 a4 a5 a8 a0 a0 97 90 85 7d 78 72 67 6e 64 63 66 66 66 5b 65 52 4e 5d 66 76 74 60 55 41 2e 1e 06 0d 06 03 06 05 03 00 06 05 03 00 06 05 14 1b 1c 1e 1a 26 2a 28 26 23 1e 26 29 2e 29 26 28 2f 31 2d 35 34 37 42 42 57 5e 6d 82 7c 92 92 86 8b 79 7a 7f 74 7a 82 83 8c 8f 96 a5 a6 ae ba bb bd c7 c6 cf d1 d1 d6 d9 d6 da da df df e6 fa ed f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f5 fa fc f7 ed f3 e4 ec ef e6 e8 e5 ec e8 ea eb ee e9 e1 e3 d6 dd d9 d9 d8 d9 d1 c8 d6 c0 c8 bb bf c0 bb be af ae ad ac a8 a4 9e a2 96 9d 9c 92 8a 85 7f 6c 66 63 60 5f 65 62 64 61 5f 56 4e 57 5a 69 78 6a 61 5a 42 35 21 0f 07 03 00 06 05 03 00 06 05 03 00 06 05 15 15 22 25 1c 1f 1a 1d 2a 2d 1e 30 24 2e 26 28 26 2d 33 2a 32 41 31 3d 40 4b 63 6e 7a 8b 90 86 84 7f 7a 80 7f 77 7e 80 80 82 8b 89 9a a5 ad b5 b5 b7 c0 c4 c5 ca ce d4 d6 cf d7 d6 db dc de ee ea ee f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f4 f6 e9 ed ee e7 f4 e5 e1 e7 e9 e2 e3 e7 e4 e0 e5 e4 e0 e9 e6 e2 e0 d9 df d4 d2 d1 c6 c8 cb c5 ca cb b9 c7 b7 b5 b7 bb b7 ad a2 a9 a4 a5 a6 9a 9c 9b 92 84 7d 79 74 67 65 65 5c 6f 68 65 62 56 5e 58 52 60 6d 77 6f 64 54 45 30 22 0b 09 08 06 06 05 03 00 06 05 03 00 06 05 16 1a 1d 13 10 1f 23 1a 24 1a 24 24 2a 2b 24 28 30 31 36 2f 2f 2f 33 3e 40 50 59 61 7c 8a 91 97 84 79 7a 78 78 79 7f 7f 7f 85 89 8e 95 9b a3 af b3 bd bc c0 c8 c5 c8 ce cf d6 da d6 d8 e1 dd e5 e3 ec f1 fe
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f7 f0 ed eb ea e9 e7 e3 e3 e8 e1 d9 e3 de e1 e3 e0 de e6 d7 e2 db e0 e4 d6 d2 cc cc ce c8 c3 c7 c5 c5 c1 c0 b9 b8 b4 b2 ac b1 a5 a9 a2 a1 9d a4 9b 95 95 89 7d 73 6b 6a 67 66 65 61 6b 6d 64 53 58 56 4c 4c 58 65 80 6c 65 56 3e 2d 19 0d 05 03 05 06 05 03 00 06 05 03 00 06 05 12 17 1d 1d 22 26 29 1a 22 2b 20 31 25 24 21 23 20 29 2d 26 29 32 34 3d 3e 4c 55 6b 79 88 95 94 7d 75 7d 7c 79 7e 7c 7f 81 80 82 85 91 94 97 a7 b0 b0 b9 bc c0 c1 cd cb ca d4 d6 d8 d9 d7 d6 de e7 de eb f4 f8 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 f3 f3 e9 eb e4 e3 e1 e4 e3 d9 dc df da db dd db d4 d5 de da de d8 d7 d9 d8 ce d5 cf c8 c6 c2 c1 c0 bd bd b5 bc ba b3 b0 ac af a6 a8 a5 9f 95 9a 9c 94 92 84 73 6f 6c 72 68 57 61 5e 64 6d 62 60 60 4b 59 55 52 5d 6a 7b 72 5f 57 44 21 20 09 07 03 02 06 05 03 00 06 05 03 00 06 05 16 19 19 1e 20 20 24 1d 26 25 28 29 27 26 25 25 30 21 28 2b 32 36 35 3b 4d 50 57 69 6f 85 9b 8f 87 79 77 7e 74 7c 7a 81 82 81 80 86 81 93 96 a3 af b5 b8 bd c1 c1 c3 ce d5 d1 d5 d7 de dc d8 dc e2 e4 f0 f7 f9 f9 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f7 ee ed e3 e4 e3 d5 da d7 d4 da dc d6 dd d0 d0 d8 dc d8 d9 dc d7 d7 d3 d2 d7 d0 d0 c4 c9 c4 cc ca bb bf b6 bb b5 b8 b4 b5 b0 ad 8f a3 9b 9a 9e 99 97 94 8c 81 77 6a 66 69 62 5f 61 68 66 6c 65 65 66 62 59 53 50 59 69 71 66 65 58 45 37 1e 07 05 04 02 06 05 03 00 06 05 03 00 06 05 13 18 19 13 24 22 24 23 25 2a 24 1d 26 1f 28 21 25 28 2d 2a 32 37 34 3b 4a 52 5b 66 74 7f 8f 99 8b 86 76 7c 78 7d 7f 79 78 80 7b 88 8b 8a 8e 98 a1 af b4 c1 c5 c1 c9 c5 ce ce cb da e0 d6 e0 e9 e4 e6 ea f2
 f4 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f2 ee ea e1 d5 da cd d5 d9 d8 cf d5 d2 d7 ce da cf d3 d0 d3 cd d5 d6 cd d4 ce c9 ce c5 be c4 bd bf bb c1 b8 b3 b2 b7 b2 b2 ac af a4 a5 9c 9f 97 98 9a 89 85 7d 73 72 68 64 65 5e 5f 65 62 65 68 71 63 5c 5d 55 5b 5d 6b 78 69 5f 57 45 2c 22 09 07 03 00 06 05 03 04 06 05 03 00 06 05 12 10 15 10 1c 20 22 2a 20 22 1d 20 23 1f 1c 25 1e 23 26 1e 25 37 33 39 40 45 57 66 77 82 9b 95 8e 78 78 75 6e 7a 7d 7b 7c 73 79 7c 88 83 89 97 93 9c ab b3 c0 bd bd c6 c6 c9 d6 d4 d8 d6 d2 de de e6 e9 ed eb ec f4 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc f6 e4 e7 df e3 da d1 ca cd cd cd cd cc d4 c8 c8 c6 d1 d2 cb ca c3 ca ce cb cb c7 c4 cb ba bd b5 bd be ba bd b5 ba b0 a6 ae a3 a4 a9 a5 a3 a1 9b 99 97 8b 7d 7e 6c 71 62 6a 63 65 5a 5e 5b 60 6d 63 69 5e 5c 5b 58 51 51 74 73 73 69 55 42 28 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 15 16 23 14 26 23 1c 23 24 24 29 27 26 27 2a 28 26 29 25 34 38 33 3c 4c 56 65 68 7a 85 8b 94 8d 8d 81 84 77 7c 7e 7f 75 79 7b 82 80 8b 84 89 89 98 a0 b5 b5 c3 c4 c7 c7 c4 cc cc da d8 d7 e3 e0 e9 e9 e7 f6 f4 f0 f7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 eb e8 e5 e1 d9 d8 d0 cd cb ca d4 cd c7 cd c2 c8 cb ce ca cf cd c9 c9 c7 c9 c1 bf bd be bd bb ba b9 ba b3 b0 b2 b2 b0 ac ad a1 a1 9f 9f a0 9e 99 95 90 88 7c 73 73 70 66 6d 64 5d 5b 60 5f 64 62 5f 64 60 5f 5e 57 5a 5e 6c 73 6e 65 4f 41 22 15 06 05 03 08 06 05 03 00 06 05 03 00 06 05 1c 1c 22 1e 21 20 1e 16 1c 1b 14 1f 1f 1f 21 1b 1f 1d 27 20 2d 37 38 44 45 50 65 6e 73 85 90 9b 94 98 81 7b 81 75 76 78 74 80 79 7e 7c 80 8d 84 84 90 9d a5 b8 bb c2 ce c5 c4 c9 cf d6 d2 dd e1 db e5 ee e8
 f3 f2 f5 f6 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc f2 e9 e4 e0 db d8 d5 cc cd c8 cb cb bf c7 c8 ba c1 c5 c5 c9 c9 c2 cb c8 c4 c6 c3 c3 c0 bb ba b3 b2 ba af ad ab ae b8 a7 a1 a2 a4 a4 a0 9a 9c 99 91 8a 8f 81 72 6f 67 65 67 62 61 64 65 64 60 69 64 64 59 62 4f 5b 4d 52 57 6b 6f 6b 5f 56 43 28 18 08 05 03 05 06 05 03 00 06 05 03 00 06 05 18 18 20 1c 19 20 19 20 15 1a 14 15 1e 1b 1f 25 25 1a 2f 25 2d 2b 33 38 44 52 63 74 79 87 93 98 9b 8c 87 79 7b 6f 78 7b 71 79 76 7a 84 7f 88 84 85 86 8d 9e a7 af be c2 c7 c7 c4 c8 c5 ce d6 d5 dc d6 e6 e2 ed ef f9 f3 f4 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ef e6 e2 dc d1 d3 ce cc c7 c7 c6 bd c4 b8 bd c0 be b8 bf bb c0 c4 c4 b9 b6 b4 c5 b8 b7 be af b1 af ad b1 b0 af ac ad 9c 9b 9d 95 a2 9b 96 a2 90 92 8d 7d 74 71 67 68 6d 61 72 63 67 65 66 6f 5b 5e 63 59 4f 4f 57 4b 55 56 61 73 74 59 52 48 2c 10 06 06 03 07 06 05 03 00 06 05 03 00 06 05 1c 21 16 1e 16 1a 1f 1e 14 1d 16 21 1f 1e 1f 27 21 1d 1d 22 21 29 35 37 4c 5b 66 6a 78 89 93 92 93 94 85 7a 70 6f 6e 73 7a 75 7b 76 81 80 83 84 85 83 88 8d 98 a0 ad c0 bb c7 cd ce d2 d2 d8 da da de e4 e5 e9 e9 ec f4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 eb f1 e6 e0 db d2 ce cd cc b9 bc c1 bb b3 be b5 af b6 c0 b5 c1 c4 bb ba b5 b9 c3 b5 b5 af ad ad ae af b0 ad a2 a6 a8 a7 a5 9a a5 95 9d 98 9a 95 8f 8e 85 83 74 71 61 61 63 6a 6a 65 64 5f 68 61 5a 5e 52 57 53 4f 51 48 50 57 61 70 68 5c 57 42 28 18 06 05 0e 06 06 05 03 00 06 05 06 00 06 05 17 13 1a 1d 1c 1a 1a 13 11 15 1c 1d 1e 1d 17 20 19 29 26 17 2a 2f 2e 39 46 5d 66 78 7c 86 93 9f 8f 8a 80 77 68 76 73 76 78 78 81 7b 79 84 82 84 82 86 8d 93 97 94 a5 b0 b5 bf c7 cd ce d0 da d7 e2 d8 e2 e7
 e8 e9 f0 f4 fd f2 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ef ec e7 de da d4 ce c7 c3 c1 ba bf be c1 b7 bc b3 b0 bb b5 bc b6 af b8 b4 c0 ba bc b7 b0 b1 ac ab a4 a9 ab 9c ae a0 a0 a0 9e 93 9a 93 9c 93 92 8b 86 74 69 67 69 68 66 65 61 6b 60 61 5f 5c 5b 59 54 58 56 55 4d 43 50 4f 51 5b 6d 70 5d 52 3a 27 1f 0e 07 08 09 0b 05 03 04 06 05 03 00 06 05 1a 1c 19 12 18 1e 1a 12 19 21 17 19 15 1b 17 14 16 1d 19 21 23 2c 25 3c 48 5b 62 70 7d 82 91 95 8a 7c 78 69 67 71 6a 72 72 71 78 7e 7a 7a 7d 7a 74 7a 85 8e 98 91 96 9b a7 b2 bb c4 c9 ca d8 d7 d3 e0 dd e3 e9 ed f5 f2 f2 f6 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec e8 eb e4 db ce d0 c9 bb b8 c0 b4 b9 b6 b0 ad b4 ab ad b1 ad b2 b2 b4 b1 b2 af ba ae b0 b0 a8 a7 a6 a8 a3 9a a3 9e a5 a2 94 9c 8b 95 97 90 9b 89 7e 76 70 6d 67 66 6b 6b 69 64 61 66 62 60 58 58 53 51 52 4d 4e 47 53 49 45 4b 4d 65 6f 60 4e 3d 2c 21 18 0d 03 09 06 0a 03 01 06 05 03 00 06 05 0f 18 1b 1b 14 1a 1e 12 13 16 17 14 1e 15 1d 1b 1b 1e 21 22 21 29 26 31 44 58 6a 73 83 8c 99 96 8e 79 76 74 6d 74 6e 74 75 78 7e 7b 7c 7f 7a 87 7c 80 85 86 8a 88 96 98 9d a8 b8 c3 c8 c9 d2 d5 da e0 e1 e2 e9 eb f0 eb fb fa f7 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ea e8 e0 d9 da ce c8 cb c0 be b8 bb ba bc aa ab b3 a8 a1 aa aa b2 af ab b0 a4 af a7 b0 ad a7 ab a5 a1 9f a0 9f 9d 97 95 97 97 95 94 94 9c 94 8e 83 79 6d 68 66 66 6c 65 6c 64 60 67 66 64 57 60 52 48 52 49 54 4c 4a 4d 54 51 4c 59 64 6f 5c 4c 44 31 2b 22 11 0e 05 06 05 03 03 06 05 03 00 06 05 17 19 14 1b 15 19 12 15 13 14 11 1c 0f 13 15 11 1e 12 20 19 18 22 30 2f 3d 57 6a 7b 84 8f 8d 8e 90 76 69 72 72 69 77 70 74 79 7d 7a 7e 7f 7b 7f 83 83 87 8a 8a 85 90 91 96 95 ab b5 bb c3 ca d3 d3 d2 e2 e6
 e7 ed ef f2 f9 f2 fb ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 ea df e0 db dd ce c8 be be b9 b6 b9 b2 b9 a6 a6 a5 9e ad a0 a3 a4 a8 aa a6 a4 af a7 ab a6 a7 a3 a7 99 a0 9e a1 99 9d 93 97 8e 93 97 95 8b 87 89 86 74 6b 67 65 6d 69 68 69 71 66 6e 60 5c 5a 56 5d 52 51 49 55 53 4e 50 4f 52 4a 5f 61 69 61 51 40 3a 2f 20 1c 06 0d 06 05 03 00 06 05 03 00 06 05 11 12 10 1b 16 1a 0a 06 18 11 16 0e 15 14 13 1b 16 18 17 21 22 19 1d 25 3d 4b 6e 70 80 8e 94 90 84 70 63 6e 6c 75 76 75 72 78 79 79 7e 7b 76 81 82 80 84 8e 8a 82 8b 8d 90 96 a2 a8 a6 ac c3 c4 d0 d6 d6 d9 e6 e4 f7 eb f5 f1 fe fb f5 fc fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ec e9 e4 dd d0 c9 cc c1 bf bc b2 b2 b6 a8 a7 a5 a7 a9 9f a2 a7 a3 a3 a3 a5 a0 a8 a3 a1 a6 a4 a6 a2 9d 9d 98 98 8e 92 93 8f 96 8d 90 8a 90 83 81 81 6e 67 6b 65 65 65 64 66 6f 6a 62 68 65 5f 56 57 54 53 4f 4e 51 4c 4b 4e 43 4c 4d 53 61 63 5e 4e 43 38 2f 25 19 12 08 06 05 03 00 06 05 03 00 06 05 0d 0f 15 0f 16 10 0c 0d 0a 1a 11 13 15 12 17 10 18 17 1b 14 24 1f 24 2a 35 45 5c 74 7b 96 9e 98 80 65 62 66 6a 6a 6a 78 6e 74 7d 7a 80 85 7e 82 77 7e 81 84 89 8a 87 87 87 89 93 95 a1 ac aa c1 c7 cd d4 d5 db e0 e8 e9 f5 ff fd ff fc ff fb f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ea e4 e2 db d4 cc c7 c9 bd b7 b3 b1 b2 ad ad a7 a0 9b 9c a2 9c 9c 9a 96 9d a5 a0 a1 a2 a2 9d 9c 96 a0 94 97 9c 98 8e 89 86 8f 92 96 8b 87 7e 7a 71 6a 68 5f 69 67 6a 64 6c 6d 6a 6d 65 65 53 59 56 52 52 4c 54 4c 52 42 4d 48 46 4e 46 54 59 5b 52 48 35 31 2a 1b 0e 0d 06 05 03 00 06 05 03 00 06 05 12 0f 1a 0b 12 0f 0a 14 0e 0d 0f 0d 0e 13 10 17 16 10 21 1a 1d 28 22 26 31 44 5e 71 7c 89 98 94 7c 69 6b 72 6a 67 75 75 77 7d 78 86 7c 80 81 82 86 84 87 84 87 8f 8c 8b 81 86 84 91 98 a0 a9 ba bf c6 cc d0
 db de e0 ed e6 f1 fd f6 f9 f5 f8 fb fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 f1 e4 da d5 d5 c5 c6 bc ba b1 b5 af af aa a5 a7 a7 a6 a4 98 9c 95 9e 9b 92 a1 9c 9f 92 99 9d 9e 9c 98 92 98 91 8a 8d 8f 92 97 8a 8d 8a 83 87 70 73 6a 65 6d 6d 66 70 69 6a 71 73 70 6d 5a 55 5b 5c 50 4e 4f 4d 46 50 4c 4a 51 4b 52 52 52 61 5f 53 4c 3d 3f 30 1e 0f 06 06 05 03 00 06 05 03 00 06 05 0c 0f 14 16 10 13 0c 05 10 14 0c 14 10 16 09 14 1a 13 25 18 1c 22 1d 1f 27 41 55 66 81 8e 8e 97 6d 67 67 65 69 70 75 72 7e 7a 7a 84 85 7d 83 88 79 84 86 8b 86 8b 86 8b 89 90 87 90 8c 8a 9c a5 aa b5 b9 c6 d1 d6 dd de e0 ea ec f7 f3 f7 fb f6 f3 fe f9 ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f1 e8 dc df db d0 cb c0 c1 b9 b4 aa aa aa a7 a7 a0 a3 a1 9f 9a 9a 94 8d 90 93 9b 90 93 90 93 91 91 95 90 8e 8d 8a 8b 8d 8c 88 8b 88 7e 81 76 76 64 61 6d 5f 65 6a 69 69 69 6b 6c 63 61 60 5c 5a 50 56 4b 4b 50 4d 48 51 49 4e 46 4a 4c 4c 4e 50 5a 4e 4c 3e 42 36 22 18 0a 06 05 03 00 06 05 03 00 06 05 06 12 0a 11 0d 06 06 05 18 0d 10 0c 10 0a 0a 10 11 17 0f 18 18 1d 23 2b 2c 36 44 64 7f 8f 93 84 69 66 5b 63 72 6f 77 73 6f 80 81 87 89 83 8e 7e 82 89 85 88 87 85 85 83 80 85 86 8f 8b 94 98 9c 99 a9 af bb c4 c5 d1 d3 d5 da db ee f4 f0 ed f6 f2 f2 fb fb ff fe ff ff ff ff ff ff ff ff fa ff ff fe ff ff fe ff fe ff ff ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 ec e9 ee fe f7 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f0 e6 e4 da d5 cc c7 c4 c0 ba ac b7 b0 a5 a7 97 a4 9c 9f 98 9d 9d 99 8e 87 99 90 8e 89 8e 90 8e 92 87 94 8e 8a 89 85 87 82 86 85 7d 79 80 75 6a 6d 66 6c 64 68 67 6d 65 6f 6a 6d 69 5f 61 58 53 52 4d 51 54 51 4d 49 4b 4b 52 4c 47 49 48 4a 4f 5b 5f 56 51 3d 3a 2c 1c 11 0a 06 05 03 00 06 05 03 00 06 05 0d 0b 10 0d 0c 0c 0e 10 0d 05 0e 13 12 13 10 11 05 0e 11 19 1e 1c 28 25 26 38 44 63 73 84 97 8b 6c 62 5b 61 66 66 7c 76 73 7d 79 84 83 8e 8a 88 87 82 7a 83 81 85 88 84 90 87 87 87 92 8a 90 96 93 9e 99 a9
 b2 b7 c0 cc d1 d7 e0 df e2 ed f1 f5 f3 ef f4 f7 f3 ee fc ff ff ff ff fa ff fd ff ff ff f6 fc ff fd fe ff fc f9 fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ea e2 cc c4 de f2 e9 dd e1 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 eb e4 d6 d4 d6 d5 cb c2 bb b6 b6 ad a8 a5 a6 a6 ac 96 a0 a0 98 99 94 99 92 91 8f 90 87 8b 88 89 8d 85 8c 83 7c 81 89 89 83 83 7a 7f 78 71 6c 68 6a 63 64 6c 63 63 66 64 6e 69 67 61 60 52 62 55 59 51 57 4d 4a 50 50 47 4d 4b 49 4e 4b 51 52 50 58 5a 66 55 4e 42 2a 25 13 06 06 05 03 00 06 05 03 00 06 05 0d 0a 06 05 0c 0a 09 09 10 0c 12 0b 0b 14 11 11 0d 0f 16 16 21 25 20 2d 26 36 42 5a 74 7d 91 90 61 61 62 65 67 67 6e 76 73 77 7c 77 7c 81 81 7f 81 84 7f 8b 7c 7c 87 83 7f 89 89 8c 95 94 95 97 96 94 98 a8 aa b4 b7 b8 c6 d0 d6 ca e9 e1 dc e7 f1 ee f2 f3 e9 ee f7 fc fd ff ff fe ff f9 f6 f9 fa fb fb fa fd fb f6 fd fc fe f8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f7 eb de ca c0 9d ae d3 e3 eb db d0 d1 e4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ed e6 d9 d6 d2 c6 c3 b6 b7 ac a8 ab a6 aa a6 9e a0 98 9f 97 8b 8c 96 93 91 8c 84 89 8c 7b 82 89 86 85 80 80 7d 82 80 84 86 77 7e 76 6e 6e 6c 66 65 66 6a 64 67 6e 71 64 69 71 65 6d 67 5a 62 5f 52 55 4a 54 4b 51 4e 4e 51 4e 4b 49 44 4f 4b 4f 54 60 5d 58 50 45 2d 28 10 02 06 05 03 00 06 05 03 00 06 05 06 02 06 09 05 0e 09 05 04 09 08 0b 0c 0c 06 11 0f 0d 19 1b 1f 25 26 22 27 32 3b 47 60 84 91 84 71 63 62 65 61 63 66 72 70 78 71 7c 7c 71 84 85 80 83 77 86 7e 80 7f 88 89 86 8a 89 84 8e 8f 95 92 94 9c 97 a3 aa a5 b4 bf bd c1 c7 cf d3 d5 dd e1 e5 e6 e4 e1 ef e6 f3 f4 f6 fe fb fd f8 f8 f6 f6 f5 fa f6 fb f8 f9 fe ee f8 fb f8 fe fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 db d5 d8 b6 a0 87 7c 91 b8 ca d3 d1 c7 c8 d8 e5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f0 e8 e6 de d7 ce cd c1 ba b9 aa a7 a8 a4 9f 9c 9a a3 92 98 94 8f 8b 8d 8c 8a 8c 82 84 82 7e 82 84 75 75 79 7e 7b 7b 80 79 75 75 70 69 5e 61 60 60 65 56 61 6b 6a 66 67 65 72 63 6b 6f 61 60 5a 5a 4b 56 4d 47 52 4a 4c 46 47 52 49 52 46 4c 4a 4e 64 5e 61 5b 49 46 33 1b 13 04 06 05 03 00 06 05 03 00 06 05 08 06 06 05 0c 00 06 06 03 04 0a 0d 07 09 0f 0b 12 11 16 1e 1d 1e 29 2a 2f 35 35 44 63 72 87 7d 65 64 62 64 68 71 6c 6d 65 78 75 83 76 79 82 75 80 7e 7d 82 83 82 83 84 80 82 8b 85 8b 92 91 8f 9b 91 9f 9b
 9e a1 a0 a5 b1 b8 b5 c4 c0 c2 cf d4 d9 dd e0 e1 da e0 e7 df ea f4 f5 f3 f2 f6 f7 f9 fb fb f6 f6 f6 fb f8 f4 f2 f3 f6 f4 f8 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff db c6 be b6 9b 7b 70 6a 75 95 aa b6 b6 b8 ba ca d7 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f0 ea e5 e1 d9 d0 ce c5 c5 b6 b7 ab a0 a2 9f 9e a0 98 9f 91 8d 98 94 8c 85 86 8a 7f 8b 86 79 7a 78 84 74 79 77 74 74 7a 7b 72 73 72 6e 64 5e 58 5f 66 5e 6c 63 6b 69 62 6a 63 71 6d 70 64 5f 5e 63 53 57 52 58 51 47 51 50 46 4a 4a 47 4e 4a 4a 50 4c 50 60 62 57 4a 4c 38 23 0c 01 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 03 0d 06 05 03 03 08 0e 11 0a 12 0c 0c 10 16 1d 22 24 20 23 35 34 36 44 52 69 7e 80 6b 63 5f 65 5f 65 75 6d 71 6f 6b 78 7d 79 7f 71 78 85 7f 84 80 7b 83 82 83 87 82 83 91 87 91 91 89 8d 92 93 93 9d 9b a1 a7 9f a5 b1 be ba c0 c9 ce cc d6 db d6 df da e9 e3 e4 ed ea f3 ee f8 f8 f2 fa f9 f9 fd f2 f4 f9 f3 f9 f5 f7 fb f7 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 d3 c2 a3 92 74 61 60 62 6c 75 8a 99 a2 a0 ab b6 cf e6 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f2 e7 db df d3 c7 cc c0 bf b5 ac a8 a6 a5 a4 9d 9c 94 99 90 8e 90 86 87 88 88 80 82 82 7c 7b 7a 79 79 71 6d 74 75 74 6f 69 70 67 69 5e 5f 5a 66 59 64 61 5d 66 69 67 63 65 64 67 69 60 64 62 5d 63 4f 53 50 4d 51 4e 4b 4f 4f 4b 4a 45 4b 4e 50 48 59 64 6b 67 62 4f 4b 37 23 0d 06 06 05 03 00 06 05 03 00 06 05 08 00 0b 05 03 08 06 06 07 01 06 05 06 07 0d 05 09 00 0a 11 1b 26 2a 2e 28 3a 39 39 50 65 81 76 63 64 64 6a 6b 6b 69 71 69 6f 74 6e 83 7e 7c 85 85 92 90 87 83 7c 84 80 7a 7b 85 8f 7e 8a 86 86 7c 83 93 90 8e 96 99 96 98 9d a2 9e ad ae af b6 bf c8 ce cd d4 d6 de dd de e4 de e8 f0 f4 f6 f7 ee ea f2 f5 fa f4 f2 fa f1 ec f6 f5 f2 f8 f6 f8 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d4 b3 a5 89 66 59 55 50 5d 63 68 6e 7c 85 8b 94 a7 c1 d3 dc e9 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e9 e8 d6 d8 cd c4 c0 c2 b0 ae ab a3 9b 91 98 92 8f 97 89 8e 8a 8d 80 84 87 7b 7b 7c 75 79 73 70 72 6f 6d 6c 72 67 65 6d 66 69 6a 5e 5e 5f 5a 61 57 5f 5f 68 62 64 5e 62 65 63 65 69 66 5b 5e 60 59 5b 5b 55 4e 50 4a 4f 54 4d 4a 49 4e 47 49 4e 4c 4e 56 6d 68 60 51 4c 30 1e 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 01 06 09 03 0d 06 0b 08 03 0b 0a 12 0d 12 0e 23 24 31 33 30 3c 36 3a 4e 56 67 65 61 62 65 6d 71 6b 6f 70 65 70 77 80 89 87 8a 8f 8b 8b 84 83 81 7d 82 79 77 7c 7f 82 7a 7d 76 84 84 86 91 80
 88 8d 8d 88 9b 8e 9d a1 a2 b1 a2 ab c0 c0 c7 c4 cc d5 d7 da db d9 e4 df eb ed f3 fc f1 f7 f5 f0 fa f5 f8 f8 f3 f3 f5 ec fb f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe d0 a2 90 6c 58 4e 4c 55 55 58 5d 61 76 7c 7f 8a 95 b1 cd d0 d6 ee ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea e1 de d9 cb ce c4 bc b5 b0 ac ac a5 9d 97 99 96 8a 90 89 89 8d 85 85 7d 7f 84 7d 75 75 72 6f 6f 72 65 71 67 65 65 5e 62 5e 62 5d 5d 57 57 54 54 5d 59 61 5f 62 71 64 65 64 58 64 5f 65 62 5f 61 5b 5b 55 4d 54 50 4e 4e 51 4f 4c 49 48 4b 47 4b 52 50 62 6f 6f 5e 4e 4d 2f 13 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 06 05 03 06 08 09 03 00 0e 08 06 0b 0a 0d 1e 2a 30 36 31 31 38 4a 4e 50 5f 5f 64 64 6f 70 76 78 7b 77 7c 7f 7e 75 80 7a 85 85 79 7f 7b 7b 7f 78 73 7a 7e 77 80 7e 84 79 79 7e 7c 79 83 82 84 89 89 8b 8a 92 8d 95 9e 9f a9 a8 ae b3 ba bd c7 d0 da d4 d8 dc d7 e4 e6 e8 f5 f2 f4 ef f1 f4 f6 f7 f9 f5 ef f1 f4 f4 f8 f1 ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 c0 8e 71 5c 47 45 4b 49 50 52 5c 60 68 6c 79 74 93 9a b2 bf c9 d5 e6 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f1 e3 dd d3 cc ce c4 ba b5 ae aa a2 9d 9d 94 9a 92 88 8b 8c 83 84 84 75 73 80 77 74 74 6d 6d 70 6a 68 71 6d 66 67 63 60 55 5a 5b 54 5e 57 51 5a 63 56 5e 5c 64 57 60 5d 64 66 5f 60 61 6d 65 5b 5a 59 56 58 50 52 45 4b 4f 4b 4d 4f 57 4a 52 4f 4f 52 55 63 6a 75 64 54 4b 2f 18 0d 01 06 05 03 00 06 05 03 00 06 05 04 00 06 07 03 00 06 05 03 09 06 0a 0d 01 0c 05 07 06 16 0b 1d 22 2a 36 3a 34 43 40 53 60 62 68 75 6d 71 71 76 79 71 69 71 6e 6f 74 70 6f 6f 7c 73 6c 7b 79 78 7e 78 75 75 77 75 76 76 78 7b 80 7e 71 7b 83 7f 7d 82 86 85 8b 89 96 92 98 a2 a4 a5 aa b6 b6 c2 c3 c5 d1 d2 de db d4 e1 e2 e7 ed eb f1 f5 f7 f7 ee f4 f2 f4 ef ec ef f8 ed f8 fb f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 be 95 6a 4f 3f 35 44 3a 4a 4c 53 52 5b 62 6c 6f 84 8b 98 a9 bb c4 d9 e4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ef e6 de d9 ce c6 be ba b3 ab ab a5 9c 8f 96 95 8e 8d 8d 7e 84 7b 74 80 76 7b 79 75 70 6b 6a 6d 5f 6f 62 61 63 5b 5e 54 4b 51 4d 59 4f 52 57 5a 56 5a 55 56 59 5d 5d 5d 5b 60 59 58 5a 5e 62 63 58 5c 56 57 4d 51 4e 49 49 4d 4c 49 4a 50 46 4b 4a 48 56 58 64 70 75 68 50 3b 2c 13 0b 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 07 06 05 03 00 06 05 03 02 07 08 07 06 10 0e 11 26 3b 3e 44 4b 49 56 5d 62 69 6e 71 69 65 6c 6e 66 71 64 64 67 62 65 75 6d 73 73 73 71 79 75 85 7b 76 77 77 7b 75 7b 73 76 71 76 73 7e 7e 7a
 7c 81 83 84 8b 80 8e 84 8e 99 93 99 a4 a1 a3 b3 b6 b9 c9 c8 d9 d7 d6 d6 e0 e3 e6 f0 ec f4 fa fa f7 f3 f5 f7 f7 f0 f1 f3 f5 f3 f3 f8 fe fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 cd 8f 5a 44 3a 41 3b 3c 4b 51 53 55 56 5a 5b 65 6c 84 92 9f aa bc c9 dd ef fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ed e1 d7 d4 d1 c2 c1 bd ab ae a9 97 9d 98 95 84 8a 81 81 7c 7e 76 7a 7a 75 6f 6f 6e 6b 68 5e 67 68 65 5d 63 5b 60 55 4c 48 4f 4a 46 50 51 51 54 4d 5a 56 58 59 59 58 5d 5c 5c 59 5b 5d 57 62 60 5d 5c 57 4f 52 4a 4e 49 4c 51 4d 4f 4f 4e 4d 4e 4d 4f 4d 5e 62 6f 6f 5f 4d 39 23 09 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 05 00 06 05 03 00 06 07 0c 0f 0d 0a 03 0e 14 1b 23 33 40 50 56 58 55 63 61 67 67 68 5a 61 5a 64 68 68 5f 5f 57 5f 61 67 72 6d 74 7a 7a 70 70 7a 7a 76 73 75 6f 74 83 7a 73 7e 7c 7f 77 7e 7f 7f 76 7a 7f 7c 85 85 83 88 89 8f 97 93 9e 9a a7 a9 b6 b4 ba c3 c2 d1 d6 d4 dd e0 e2 eb f0 eb ef f6 f2 e9 f6 f9 f3 ee f3 f2 f5 f7 f4 fa fb ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb bd 84 50 44 38 34 3e 3b 42 4f 47 49 4f 5a 61 5f 6a 73 89 95 9f b7 b9 c2 d8 de ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ec e6 e1 e0 cc c9 c4 b9 b8 a5 a9 9e 9c 9a 91 91 8b 82 7f 7f 80 7b 75 78 7b 70 70 6f 70 63 61 6c 5f 60 5a 5a 54 59 56 4c 4d 4c 4d 53 4c 4a 51 54 4f 51 55 50 56 5a 57 59 5a 5b 5e 5b 5d 61 5f 62 64 5d 5d 57 52 50 50 50 53 46 4e 51 49 4d 4c 49 45 52 4f 4a 60 6b 67 6b 5e 49 36 1d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 06 03 08 06 05 0e 0a 0f 14 11 22 18 12 27 30 36 4b 52 4a 56 49 58 66 5c 5d 5f 5d 61 5d 63 64 5b 63 5d 69 66 70 74 70 74 78 71 6c 74 74 77 7a 77 6e 72 73 79 7d 77 7b 78 79 70 77 7b 76 72 82 79 76 7e 85 7e 84 8e 90 89 8c 96 99 9a a2 ac a5 aa ba c0 c6 cd d7 d6 d7 dd e4 ea ef f4 f2 f4 f7 f4 f8 f7 f0 f0 f4 f1 ed eb f4 fb f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff b1 73 50 41 2f 27 3b 37 41 43 42 4e 4c 55 5c 59 6c 6e 7c 82 8f 9f ac bd c3 db e8 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e8 dc d8 d6 ca c6 c4 b6 ad b0 a5 9f 97 8e 90 82 83 7f 77 7c 74 72 65 6c 75 6b 6c 6a 57 5b 5c 5c 5f 4e 4f 4d 4d 43 53 3f 45 3e 42 4d 48 48 4a 50 50 4f 4f 46 54 50 5a 55 57 58 59 5f 5e 5e 5b 5e 60 5a 59 50 53 51 52 4e 54 46 47 4d 4c 50 49 4f 4a 4b 4e 50 66 6e 78 6c 5a 42 2d 13 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 08 12 14 13 1b 14 16 1b 16 0e 0d 14 14 1f 31 3a 47 58 52 57 65 6a 61 5e 50 56 5a 63 5d 61 64 64 67 69 6d 72 74 6f 6d 66 6c 72 78 75 76 72 71 72 79 76 78 76 74 74 79 72 75 74 6c 78
 73 71 78 78 75 7b 7b 83 83 86 87 85 92 99 9a a3 a4 9b a4 b8 b4 c3 c7 c2 d6 cb dc d7 e4 ea eb ef f8 f6 f6 f7 ec ef f7 ef ec f6 f5 ff f7 fe fb f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff bd 6b 4a 38 26 26 33 37 3f 48 4f 41 4e 4a 4c 5f 60 5e 6a 76 77 8d 99 ae bb cb dc db eb f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 ef ed db d8 c2 c9 bc ba b3 ab ae 99 95 91 8f 8e 85 84 7b 76 70 78 6e 6e 6e 69 68 5b 60 5e 5c 5f 4d 54 4d 4f 49 4b 44 3d 45 43 3f 44 4a 46 4b 48 45 4c 45 51 4e 52 55 52 59 4d 5b 48 55 64 5d 56 62 58 4b 56 59 4a 51 51 52 4f 47 56 52 4c 4b 4d 46 4b 51 53 52 60 71 78 69 59 3c 26 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0c 14 14 10 16 18 0f 12 13 0d 07 07 0e 05 06 05 0a 17 27 3c 46 59 5a 58 68 64 6d 62 5a 52 54 61 5a 64 5c 65 6a 65 73 71 6a 6e 6c 6d 64 6e 76 72 73 74 72 75 70 73 74 71 6f 71 74 71 6d 72 74 72 74 78 79 74 7d 7e 87 7e 83 82 88 8b 8e 94 8d 94 9b ab aa ae af b5 b9 cd ca d0 da d6 de e9 e9 f2 f2 f8 ff fb fa f7 f6 f3 f5 f2 fd f8 fd fe f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb bf 6b 4b 36 24 27 2d 3a 3b 44 44 47 40 4d 55 52 5c 5e 65 6e 7a 86 8d 9b aa b4 c7 cf da e7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 e5 dc d3 ce c5 cb bb b6 b2 a5 a3 a1 9a 8d 89 85 7a 7c 77 79 73 75 74 6c 6c 66 5f 63 5f 50 58 4b 57 4a 47 4b 41 42 3c 41 43 45 45 3e 49 47 4b 52 4c 50 40 50 4f 52 49 4f 4b 4e 4b 4e 55 5c 5d 60 5b 5e 5a 5c 60 54 56 4f 55 50 4e 4d 47 4f 56 50 56 54 49 51 55 65 73 6f 63 4d 36 23 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0d 0b 07 05 06 06 05 06 03 06 05 03 00 06 05 0c 0b 21 3c 4a 58 6a 66 66 67 5f 5a 55 5d 58 5e 54 62 61 6b 60 6a 68 6c 6f 6a 68 65 65 6a 74 75 75 70 72 74 71 69 6f 6c 6d 74 6b 72 6f 68 6d 6b 6d 6c 76 70 70 7b 72 7c 81 89 85 84 88 8c 94 93 9e 9d a6 a7 a8 b2 b8 c3 bf bb cd d0 d7 d6 e5 ed f6 f8 f6 fb f8 ff eb fb f6 f3 f5 f9 f9 fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 a8 68 43 37 2b 1a 2d 2d 35 40 3f 45 40 43 4b 50 4c 56 59 71 6a 78 83 8a 96 a6 b3 c3 ce cf da f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 e9 e1 dc d3 cf be c5 b5 bb b3 9d a3 99 94 92 8a 81 7b 7b 74 72 70 64 70 68 6b 62 5e 59 53 51 52 48 45 39 3a 41 3d 3f 3a 3e 3f 3c 39 3a 3e 48 42 41 47 45 49 45 53 4c 4f 4d 4e 54 4b 55 59 54 55 57 59 54 59 54 57 52 52 51 51 54 54 50 4f 52 53 50 54 48 4e 51 57 65 6c 69 5f 43 29 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 02 06 05 03 00 06 06 03 00 06 05 0c 10 16 34 4b 5d 71 66 63 62 5b 54 4e 5b 51 5a 5c 5d 65 60 64 68 57 5d 60 60 5f 69 6e 6f 68 71 6c 64 76 66 69 63 65 6a 6b 6e 6a 6f 71 6a 66 6a
 68 76 72 71 68 72 71 6f 7a 77 79 85 87 7b 8f 94 94 a1 a5 b4 ab af b5 b5 bd c7 c2 c5 d4 d5 dc e4 e9 eb f8 f9 f5 f9 f6 f1 f6 f2 f6 fd f2 fc fd ff fd fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e7 a7 6b 42 2d 1f 1c 26 29 31 3a 3a 3e 44 3e 41 45 46 51 52 5a 5f 6b 77 7a 94 9b a7 ae ba c9 d2 e5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea e7 d4 d3 c1 cd bd bc b0 b4 af a4 a6 9a 90 92 7d 82 80 75 79 6a 73 6d 68 65 69 5a 55 4f 4d 4b 47 44 38 3c 37 3a 3a 45 37 2f 34 39 3b 3f 3a 3b 44 45 48 44 43 48 48 45 4f 51 49 4b 48 4f 50 52 50 58 50 4e 52 52 51 55 52 51 47 54 4a 53 4b 4d 51 4c 4b 4c 4b 59 55 6b 70 62 51 35 1f 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 06 0a 15 27 41 60 72 72 6a 5e 5a 5d 55 5e 57 5c 61 69 5e 60 61 59 5b 5f 5f 5e 69 62 71 67 69 67 69 6e 6b 65 68 67 5b 6d 66 61 6e 6a 66 66 6c 71 68 74 6d 6c 70 71 79 75 70 74 79 7a 7d 8d 86 8b 8c 9a a4 a5 ac ab b1 af bd bd bc c9 cc ce d6 e1 e6 ef ed ef ed f3 f4 f6 fb f5 fc ff f1 f6 f8 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e0 a1 64 3f 29 1e 25 23 2f 30 39 33 36 47 42 45 44 45 4a 4f 5a 5e 67 6d 70 7e 8c 94 97 a9 af c2 d5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 eb de d2 d7 c1 ce bf b9 b9 b0 ab a4 97 9c 90 8c 7d 7e 80 76 71 75 66 6f 70 60 5b 58 50 4e 4b 40 3e 43 3b 3a 3e 3b 35 35 35 3d 36 3e 35 39 3c 44 48 45 4a 43 43 45 49 47 48 55 46 57 4f 4d 55 4c 54 51 4c 57 53 5b 56 5b 5a 53 52 4f 51 4f 4d 54 50 50 50 54 4a 54 66 66 66 5b 45 1f 0c 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 05 09 14 22 38 58 63 72 7b 65 60 60 55 5e 57 64 63 65 64 6a 63 60 60 61 64 6d 6e 64 68 69 65 70 6e 69 65 5e 64 63 62 68 6a 5e 61 62 6b 67 6d 67 66 6a 6d 71 6c 6a 71 77 74 7b 75 77 7f 7b 84 85 87 95 9a a2 a4 a9 b5 a9 b5 b9 b8 c3 c5 c1 d2 da dd e3 ed ec e8 ee f3 f1 f3 ef f8 fb ff fa fb fe fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 dc a4 6d 41 2f 20 1c 23 2a 34 3e 35 39 33 3b 38 3d 45 44 4d 4b 54 61 5c 71 71 7c 8a 89 95 a2 b1 c7 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 dc d6 ce c8 c5 b7 b6 b6 b3 b0 a7 9c 9e 91 8a 86 91 82 82 7b 74 6a 68 5b 62 58 4e 56 3a 46 40 3b 3f 39 36 38 34 30 38 36 37 39 3d 38 37 3c 45 41 3e 42 48 3f 42 4b 42 40 44 50 4f 4b 4a 4e 53 46 50 50 4f 53 51 55 52 54 59 4f 55 4e 46 53 4f 5a 4d 4f 4d 54 4d 56 62 68 62 4b 33 19 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 06 13 14 1e 35 53 64 7a 6d 60 5c 5d 55 5b 62 64 5f 5e 69 5e 57 5f 57 5a 58 69 67 65 6d 68 69 6c 62 67 5b 5e 60 58 60 5e 64 65 61 63 6a 65 67 65
 6c 67 66 68 67 6b 70 72 6d 75 6f 7c 77 77 7b 84 7f 84 8e 93 9d 9e a9 af b8 b6 b1 b9 bf c4 ca d0 d2 d4 d1 ea e9 e3 e8 ec fa e4 fd f3 f1 f8 f4 ff fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee d2 9b 71 4a 2a 19 15 1a 23 2a 35 36 32 30 31 39 3a 37 39 3d 4c 4b 51 59 5f 62 6f 78 77 88 94 a0 b0 db ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e8 de da c6 c6 c3 be b0 a9 ae ac a3 9e 9a 9b 98 8f 86 7d 7f 78 6c 6c 63 60 53 4a 49 45 3d 3d 3e 3b 33 36 38 33 2e 35 33 30 36 30 34 41 31 32 3c 41 45 3c 35 42 3c 43 3e 47 44 4f 46 54 3e 48 48 47 4d 54 4b 54 4d 52 56 54 50 4b 52 56 47 4d 4b 54 51 53 4e 53 53 5a 59 60 55 3b 28 15 09 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 07 0d 1a 23 4c 69 7b 72 69 5d 5e 5d 6d 65 68 6b 6c 60 64 57 5f 55 5f 5c 60 66 6a 61 69 6c 6b 67 5e 59 54 5b 5b 5c 63 60 5f 5d 63 63 64 68 67 63 6b 5c 6a 6e 63 73 6e 72 6e 70 77 75 76 81 7e 79 83 83 86 8b 90 98 a6 a8 ae bb b7 bc bb b9 c4 cc d0 d8 db db dd e1 e1 ec ee ef f1 f0 f9 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ee d3 a4 79 47 2f 17 1a 22 1f 24 31 33 29 31 2f 2f 32 39 35 3a 47 43 4c 56 52 61 67 66 6f 78 87 91 a0 ce ff ff ff ff ff ff ff ff ff ff ff ff ff fe f0 e6 dd d2 c7 c0 bf be bb b2 b5 a7 ab 9e a4 9c 95 8d 8f 8a 81 7c 69 6a 6b 5a 53 51 49 47 41 33 34 33 36 3a 34 2d 33 37 34 33 38 34 33 35 37 40 3a 45 40 40 3d 41 45 3f 3c 47 47 43 43 51 49 3e 43 47 4c 51 4c 52 52 49 4d 51 4a 4d 4c 52 4e 54 53 53 4c 52 51 57 56 4e 4f 4f 4f 49 2e 1b 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 0b 06 06 1b 25 3c 64 78 6e 68 5f 58 59 67 65 6f 68 6d 6c 64 61 5d 59 55 5f 59 61 61 60 65 64 63 64 61 5d 59 52 5c 5d 60 66 62 5f 60 62 5b 60 60 64 66 6c 63 60 67 69 64 67 6f 6e 71 76 7e 77 76 7d 7f 82 83 84 86 8f 95 9c a4 ad ae aa b0 c0 c1 cb c6 cf d0 d4 d8 dd e4 e3 e5 eb ea ec f1 f1 f6 fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f6 ea d5 a9 80 49 29 15 12 14 22 25 2b 22 2b 28 29 2a 2b 2a 3c 33 40 4c 41 4a 55 4e 62 61 6c 6a 7f 84 8d b9 f8 ff ff ff ff ff ff ff ff ff ff ff fb e7 e0 de d5 c8 ca bf bf b7 b5 b1 af a5 a7 9b a3 a0 95 8b 8f 8c 82 79 6b 5d 52 52 49 49 3f 40 33 3f 36 31 36 31 31 32 29 34 37 35 35 31 31 34 37 37 41 42 34 34 3c 3c 4a 3c 46 3e 42 3f 4b 4a 4e 4b 40 44 42 49 4b 49 55 4f 53 52 50 55 4a 4c 54 50 4e 4d 52 4f 4a 4e 51 4f 4b 48 42 34 20 19 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 0e 19 15 34 4d 75 73 71 68 58 5d 5f 6e 64 6f 6f 64 5d 57 5a 60 60 61 5e 65 59 62 59 62 5b 5e 65 5d 5d 59 5a 5f 60 5d 5f 69 6b 65 64 6a 64
 62 60 61 60 63 5e 66 6b 6b 6a 6f 6c 6c 77 75 7e 81 7d 77 7f 78 7b 85 8a 97 98 9e 9e a6 af b5 b4 bb bb bf ca cc d3 c8 d2 d9 da de e4 e3 e8 e5 f0 f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe ff fb e9 e0 bf a0 58 25 10 0e 1c 1f 19 29 20 1f 1d 26 26 2b 30 2b 37 35 3d 42 41 4d 52 4d 59 5c 61 69 6c 81 a2 ef ff ff ff ff ff ff ff ff ff fb f6 ee e7 d4 d1 c9 cb cb c4 be bf af b0 b2 a3 ab a2 a4 9c 96 92 8e 82 76 6c 64 51 50 44 41 40 39 3c 34 36 31 35 35 31 30 2f 31 36 31 2c 38 36 33 3f 39 37 39 35 34 39 3a 34 3b 3c 3c 35 3e 44 3e 3e 3e 3d 40 4b 3d 45 46 52 44 55 57 4d 50 4c 4d 52 4a 49 46 4f 52 52 4d 44 4e 47 4a 3e 3b 31 1e 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 07 06 05 0a 0b 0b 0b 1f 30 4b 6a 77 71 67 56 5a 61 66 6b 66 62 64 5c 62 5e 5e 5f 5a 62 5a 63 64 6a 73 64 65 64 5d 61 5d 5d 66 61 62 63 64 66 69 6a 64 64 68 66 69 64 68 64 68 6f 67 6f 6b 70 78 7b 70 7b 7f 76 82 7a 72 74 79 7c 84 90 8a 9e 9f a4 af b1 b9 c0 c0 c3 b9 c1 c2 c6 ca d0 d4 d9 d5 da de e5 f0 ef f5 fb fe fe ff fc ff ff fe ff ff ff ff ff ff f6 ff ff f1 e5 d6 a9 64 27 1b 0d 11 16 21 24 21 24 27 22 22 24 2e 2f 30 3c 36 43 40 43 49 4d 57 51 5e 5e 66 74 8d d2 ff ff ff ff fd ff ff f9 f9 f5 ed ec d7 d6 d2 c5 c9 b8 b8 b4 b5 b6 ae b0 a8 a3 a0 9d 93 8f 7e 78 6a 62 69 5e 56 53 45 48 3d 3f 41 32 30 31 2d 2b 36 31 34 32 36 34 33 35 37 33 3b 33 31 34 36 31 3b 38 3b 41 37 3c 3d 40 45 3e 3b 3f 41 3c 45 44 4c 4e 4d 46 4c 4d 51 58 4f 52 53 55 4c 50 4f 4d 51 50 4d 50 42 49 3e 32 30 27 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 10 0e 15 1f 22 41 54 72 6d 6d 5d 5c 5f 57 58 63 5d 58 5c 5f 62 65 64 6a 66 69 60 72 67 6e 5e 60 63 65 58 5b 5f 5c 65 66 65 67 64 61 64 60 69 63 6a 66 63 65 60 67 61 70 6a 66 71 73 79 75 81 7b 7b 76 7b 72 79 76 76 71 79 85 89 92 92 9e a7 a4 a7 b2 b1 b5 ba b4 b8 c5 be c9 c5 c8 c7 d1 d7 d5 db db e5 ee f5 f5 f5 ff ff ff ff fd ff ff fc ff f5 f4 f5 ec dd dc bb 6b 29 18 14 12 1a 1a 22 1d 28 23 25 1e 1f 23 2b 2a 2e 37 35 3d 36 40 4c 4e 50 55 5a 60 5e 80 c2 ee fd ff ff f4 fc f8 f3 e6 e7 e6 d5 cf ca ca c5 b7 ba ba b7 b0 b4 aa ad a4 a1 97 97 84 7d 7d 6b 63 60 58 48 4c 47 41 42 3f 3c 35 43 3c 31 36 36 30 34 3c 2b 33 39 38 3c 3a 3b 34 2e 2e 33 38 32 33 38 39 33 36 35 3a 35 34 41 3f 47 41 4a 43 47 4c 4a 46 4b 4a 4e 51 53 50 4f 48 53 57 51 54 4f 54 4b 56 4b 4b 3d 36 32 1e 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 06 01 0c 09 16 1b 36 50 64 75 65 64 55 50 59 5b 5b 5a 5d 59 5d 63 67 68 69 66 72 63 5b 61 60 63 60 51 5d 59 57 57 57 60 61 5f 66 6e 5b 5d 61 64
 61 6a 61 64 66 6b 65 6c 6b 6d 67 78 75 6e 81 7c 79 76 73 74 73 66 73 72 77 6f 74 79 79 84 8f 90 96 99 9b a8 a1 a6 a6 a8 b6 a6 ae b4 b9 bb bb c1 c7 c1 cb ce d4 de e0 e0 e8 e1 ea eb e9 f0 f6 f0 f3 ef f4 ee e7 dd e2 c5 73 2b 11 0b 17 10 0b 18 1c 1a 14 1b 19 1c 23 1e 29 31 2b 2d 34 35 3c 44 46 4b 42 4e 4a 5e 6a ac df e8 f6 f1 e4 e8 e9 e5 e4 e0 cc d3 ce c1 be b4 bc b6 b2 b4 b0 a3 a0 9e 8f 95 85 83 76 6f 69 64 59 5a 4d 49 46 46 3b 3f 35 3e 3b 35 34 30 39 3d 33 33 2e 33 26 34 32 30 31 2d 2d 3a 2c 2c 37 2c 34 34 36 33 37 30 3e 35 35 3f 3b 39 3f 3b 3d 44 4a 46 4a 43 4b 4d 4b 51 4e 45 54 4e 55 50 4e 4a 4d 4d 4e 47 3f 3b 2f 25 23 06 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0b 0f 14 10 22 27 45 5a 6f 6e 5e 5c 52 59 5c 59 55 50 56 61 59 6a 66 6b 65 6e 6f 68 64 5e 61 62 5c 54 56 63 59 57 5e 54 5e 5f 63 64 64 69 68 69 60 64 65 5c 66 62 68 71 70 74 76 79 82 72 7d 7b 6c 72 6d 6c 73 68 72 6f 75 75 77 74 7d 7f 81 80 8a 8a 94 91 95 9d a0 9e a3 ac a3 a1 a3 a1 a7 b1 ae b4 bb be bf c3 c5 d1 d5 d9 d5 d3 d6 d4 e0 e1 e2 e4 d4 d9 d9 d6 cb 74 2a 16 0c 0f 0c 0e 15 15 1f 1d 15 0b 13 21 22 20 27 2a 35 2b 34 3c 42 41 3c 40 44 4d 4d 64 9e d7 df e1 ee dd e5 e4 d7 db d1 cd cb bf bd bb b6 b5 ab a2 a1 99 9c 8a 8c 88 84 73 76 65 65 5b 55 49 54 4a 4b 49 4a 44 45 44 39 3c 35 30 2f 33 30 35 36 32 2f 36 36 33 39 30 2a 31 2b 2c 30 31 31 38 35 30 29 32 2a 2f 3d 32 37 3c 38 46 3e 3b 3e 41 45 42 44 43 45 4f 4b 53 45 4d 53 4f 4e 50 50 49 47 45 45 4a 39 30 25 0e 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 04 12 09 14 18 21 27 38 51 62 6f 69 60 58 5b 5c 59 62 59 58 59 5f 5e 6a 6a 6f 69 6c 67 63 60 5a 56 61 5f 54 5b 4f 53 5b 5a 5b 5d 61 57 5a 5d 62 65 6d 6c 66 65 64 70 72 6e 7e 7d 7d 7b 7f 7c 76 74 79 72 76 6e 71 77 72 7a 6a 6d 73 7c 74 7c 7f 7a 85 7d 8d 8d 8e 8b 95 90 99 94 9a 9b 93 9a 9f 98 a5 a6 a0 a4 a8 ad b2 b0 b4 bc be b9 bd be be bd bf c1 c6 c3 c8 c6 b7 73 2a 17 0c 10 10 14 1e 1e 23 14 21 12 11 21 20 1a 21 20 2c 2e 2d 2f 32 42 38 3f 47 4c 52 4f 8e cf d5 d8 de d1 d7 d8 db c9 cd cb c3 b9 b5 b7 ab a4 a3 97 93 92 8b 81 81 76 69 73 6a 5e 5c 5b 58 4c 4f 4c 49 46 44 41 44 43 44 44 48 3f 36 40 38 3a 37 34 32 2b 33 34 34 35 2d 2b 31 29 2f 36 36 37 34 35 34 36 37 41 43 35 3a 31 43 43 42 46 4b 3d 4a 4b 4b 52 45 4f 4e 49 4c 4c 53 53 4d 59 50 51 56 4b 4b 45 3b 29 21 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 10 0c 13 18 13 34 3f 56 6f 65 5a 5e 56 51 55 51 5a 56 53 5b 56 58 64 61 59 64 5c 5f 59 5b 5d 59 56 57 55 52 55 4f 51 51 56 61 4f 51 4f 58
 63 67 61 62 6a 62 6d 72 70 74 6e 7d 7d 79 7b 79 6e 78 6f 75 69 72 71 6d 70 67 6f 76 6a 6e 76 7b 74 77 75 74 7f 82 75 84 7f 87 86 84 89 87 83 79 90 89 90 9a 97 98 9c a1 a2 a0 95 97 9c 9d a0 a6 a8 9f a0 9c a0 a5 a0 9f 6a 26 0e 09 13 06 0c 13 15 1e 13 17 13 16 15 1c 17 22 22 25 25 30 31 37 34 37 38 3a 35 4a 47 86 b7 d6 d6 d2 cb ce c5 bc c3 b6 b4 b1 a7 9a 9b 88 92 8f 8a 87 7f 76 6c 71 61 67 5f 5d 5b 55 4f 4c 4b 42 47 45 4a 49 3f 3d 41 39 42 41 3b 3a 3c 3d 37 34 31 2f 33 2a 34 31 32 2b 2a 32 2f 29 27 2d 3a 34 38 2f 32 2e 31 3a 39 3a 3a 3d 39 3b 47 38 41 45 4a 4b 4f 46 4a 4e 54 4a 52 4f 51 4f 51 4e 50 4a 4e 41 3e 33 15 17 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0d 0f 18 18 18 1b 26 28 47 5d 63 5a 52 50 50 55 55 54 58 4d 58 57 56 58 4e 5a 52 55 5a 55 5d 5a 5a 59 62 52 54 55 54 4c 56 50 58 56 5b 60 56 52 5d 53 60 64 68 6b 6b 70 75 6e 6e 71 74 79 79 78 70 74 71 71 68 6b 68 6f 68 70 6f 70 71 72 6f 76 79 76 80 78 73 70 7a 76 7a 7a 69 74 76 72 79 77 72 79 85 85 89 86 8a 88 94 90 8b 8c 8f 95 8c 8d 90 94 8a 88 82 8a 84 55 23 12 06 09 10 12 0e 16 1e 11 18 0e 0e 13 12 16 15 1c 24 1e 22 2d 2a 37 32 3b 3c 37 38 49 6e b3 c3 c0 c0 b3 ad af b1 a6 9f 9a 95 97 8a 87 84 7f 7c 7b 75 73 66 65 60 57 56 5f 53 52 51 4e 4e 49 45 4f 47 42 3d 41 41 3e 3a 43 37 36 39 40 39 3a 32 35 3a 34 36 35 31 2d 2a 33 29 2c 2f 35 25 27 2a 32 2b 2c 35 32 30 36 34 37 3f 3b 42 3d 3e 46 3a 44 44 48 48 47 4d 46 50 49 4e 47 4d 50 52 50 4b 4c 3e 2f 29 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 0d 0a 13 19 1b 19 25 36 55 65 60 5a 58 51 54 54 4b 55 50 55 4d 58 50 59 4b 53 4e 4f 57 54 54 5e 59 55 53 55 55 56 60 5a 56 5c 52 5f 66 55 5b 60 62 61 5c 5a 5b 64 5e 70 6a 70 78 70 7b 72 72 77 7c 77 72 70 6b 73 70 6f 7a 74 7a 77 6b 74 74 70 73 76 6b 70 71 6e 70 65 68 67 6d 66 6b 6e 6f 71 73 68 75 7d 83 76 7f 84 7f 85 86 84 80 84 76 7f 83 7a 77 85 79 70 58 1e 0c 08 13 0d 0b 07 1c 11 20 10 07 07 14 0b 12 17 12 1a 1c 22 2b 25 24 30 2b 31 33 31 42 69 a2 a7 b0 a5 98 9d 9d 9b 95 93 83 7f 7d 80 7b 77 77 72 67 6c 5f 5f 58 5f 5b 56 4b 51 4e 49 54 45 44 45 3f 3d 3e 43 41 35 3a 35 3c 34 36 3e 34 40 3b 3b 35 34 2c 32 32 35 3a 2e 2d 2c 28 29 2d 2c 2e 37 34 38 2b 30 33 32 3a 44 3a 42 38 3f 38 44 42 48 47 45 46 42 51 4d 4e 46 56 54 45 50 50 50 56 4b 45 3d 31 24 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0a 14 14 18 12 15 22 36 43 55 5a 55 5a 51 53 55 52 4f 50 55 4b 54 4f 55 52 47 49 52 4d 59 57 5c 5c 58 57 58 5a 5a 5a 52 55 54 56 5c 5c 5f
 5f 6c 6b 68 68 60 5d 5f 6b 61 69 64 70 76 70 71 7a 73 73 6f 74 75 70 78 78 71 6f 6f 76 70 6b 75 76 72 69 6c 5c 68 6b 66 6d 5f 65 64 6b 5e 5f 63 6a 6c 65 70 6a 6b 71 66 76 74 70 6c 6e 7e 74 72 72 77 70 72 68 6e 6d 67 4c 24 12 10 0a 0c 09 0f 13 14 15 10 0c 0c 0e 12 15 0b 1a 1d 13 19 27 1e 20 2a 29 2b 30 2f 36 59 7d 91 96 8f 7e 8c 8b 78 86 7b 82 77 6d 6d 66 69 62 5b 5d 54 55 54 53 54 49 50 4a 54 4d 4e 47 3e 41 43 3f 42 3e 3c 3a 3a 3a 39 35 35 31 30 36 3b 33 35 30 30 36 32 36 33 33 2f 2d 37 2b 2f 30 35 2c 31 32 28 28 2e 32 2d 33 3c 36 3a 36 3d 3a 3e 43 43 44 45 41 50 4a 50 4b 4f 53 54 49 4c 55 51 4e 46 48 30 22 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 11 0c 15 16 1a 1b 25 29 36 51 50 50 52 53 4a 53 4d 53 46 4a 51 54 51 58 54 4d 50 50 50 4f 4f 55 55 56 52 5d 55 50 5b 50 56 59 57 5d 59 4f 5a 65 67 60 62 5c 5a 5a 5e 62 67 5a 62 64 62 6e 6d 6f 6e 6b 70 6c 79 69 74 71 75 71 73 70 6f 76 70 6a 6e 60 6a 66 66 5f 66 5b 63 62 57 5a 5d 63 60 63 59 55 62 60 66 69 69 70 6a 6b 60 6a 6e 6d 68 61 5f 5d 5b 5f 59 58 44 1f 11 05 04 0c 09 15 10 18 11 10 10 09 09 05 07 08 09 0f 0c 18 1a 21 28 26 27 2a 2f 1f 2b 48 69 71 76 74 6e 76 6e 72 68 70 67 6a 63 66 62 5c 60 64 5a 5e 56 5b 50 52 4a 46 4c 49 41 48 4b 49 44 44 40 3b 34 41 36 3f 36 32 38 39 34 30 36 35 2f 28 28 2c 33 34 31 38 31 32 2c 2f 2c 30 27 25 2d 2c 2a 2f 2c 35 39 39 3e 36 39 36 3d 41 43 3f 43 46 41 47 49 44 4e 46 49 48 4f 52 52 4d 55 45 47 44 3d 35 1c 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0b 12 15 16 11 1b 20 35 40 4f 48 49 53 52 51 4c 4f 53 4a 44 4b 51 4f 4d 4a 47 4c 52 50 4e 53 52 51 4a 48 55 53 53 52 4c 4e 53 54 52 50 5c 5e 5d 5e 5c 5e 58 63 5a 5d 57 5c 61 60 5d 5e 6b 66 6c 64 66 6e 69 72 70 72 72 68 67 75 69 6d 68 5e 5d 65 62 62 64 52 5c 61 60 61 5a 61 54 5b 5a 54 5b 63 5b 5c 67 61 68 62 6d 66 5e 5f 5b 5c 59 5f 5b 60 5a 54 59 53 41 19 15 05 0b 03 07 0f 17 10 0f 13 06 0c 0e 09 0a 09 0a 0f 10 10 0f 20 21 19 22 24 27 1e 21 39 5c 60 6d 6c 69 67 65 64 5c 66 62 62 62 58 59 5c 58 5b 51 4a 56 4d 4a 52 47 49 43 52 3f 4e 4d 45 48 45 40 40 33 38 37 3c 35 39 35 31 2f 34 36 33 2c 31 31 38 35 31 2d 2e 2e 2a 2c 32 29 32 29 2e 2c 31 2a 2e 32 2f 34 2f 3a 3a 32 3e 3b 3e 3f 42 46 42 44 4a 40 50 44 4e 51 4e 53 52 42 4f 53 4e 48 40 38 1e 12 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 16 17 15 1e 22 1e 30 37 40 50 4e 46 49 50 50 56 51 4c 52 4b 50 5a 4d 4c 50 4d 4b 4e 53 51 4f 47 4f 4a 51 58 56 50 55 50 4f 4c 4c 50
 4f 57 59 57 55 55 57 5a 53 58 57 60 61 5d 5c 55 67 60 5d 64 60 64 5c 63 64 69 68 72 67 69 65 65 64 60 59 5d 5b 56 53 55 61 55 58 63 5f 51 5a 5c 58 5b 5a 61 58 60 6a 66 61 67 64 64 5d 5f 59 5b 59 60 5a 4d 55 52 57 4f 3f 1c 0d 09 07 03 0b 13 10 11 11 07 03 0c 06 05 0a 03 06 0c 08 10 12 15 17 1f 1d 1f 1e 24 29 32 4d 5a 5e 5e 54 5a 5d 60 5b 5c 56 56 58 52 5d 59 58 59 56 55 4c 48 4b 4f 3e 48 51 44 48 40 3e 47 3b 3b 43 37 42 3f 3e 3e 3c 39 3b 39 32 28 39 35 2e 31 29 35 35 30 26 36 33 2d 35 2e 2d 2c 28 28 2c 2f 29 30 30 38 32 35 38 3b 38 36 45 39 39 3d 44 49 45 4a 41 48 4d 50 5b 59 52 52 4a 53 48 44 47 3d 36 1c 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 0e 0b 1f 1d 24 23 27 32 32 40 48 49 51 58 53 4e 49 4f 46 4d 49 4f 46 51 47 50 57 51 4e 4f 4a 46 4c 45 52 54 4d 3e 44 4e 52 4c 4a 54 52 54 4e 4d 4f 56 4e 4c 51 52 56 4c 5a 56 67 5d 59 54 65 59 60 60 5e 66 69 6c 62 69 60 62 65 61 5b 5f 5b 5c 5c 5f 5c 54 5b 58 5c 56 54 5d 5e 52 52 5d 5f 53 5b 60 6b 6a 62 5f 5c 5c 54 58 54 55 53 4b 53 52 53 4b 4d 47 3d 19 14 0b 0a 05 06 06 12 13 0b 09 0a 0f 07 05 03 0a 07 07 07 0d 0d 0c 10 10 15 19 1b 20 1b 2e 3e 58 4c 4f 50 52 5c 58 58 56 53 54 5b 50 5c 5b 4b 58 55 50 4e 4c 49 4c 50 45 49 41 44 40 45 46 41 42 42 34 3a 3a 38 39 35 38 34 34 37 38 32 36 30 2b 2d 32 32 29 29 33 33 35 32 2b 2e 2f 2a 2d 2f 30 27 29 2e 35 34 34 2f 37 39 3c 3d 38 36 3e 45 3e 43 47 45 50 55 50 55 55 4d 52 3f 47 46 44 48 32 2a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 0e 0a 19 1c 23 24 21 29 2d 3a 44 46 40 59 56 53 53 4c 49 4a 4f 4b 4a 4d 4b 4a 48 4c 4c 49 4b 4e 4f 47 49 4c 50 51 4c 52 53 45 4f 4b 4f 5a 50 4d 4d 4e 53 51 4e 55 56 4d 56 48 60 57 57 5b 56 52 5d 54 51 60 5b 60 60 68 64 61 63 60 5e 5d 5e 5d 5a 54 53 56 5b 5d 5a 55 55 54 59 59 4e 58 4e 58 55 5c 59 63 5c 54 5f 58 54 53 56 54 4e 4d 4f 4e 46 47 4b 48 42 3a 1f 0e 09 06 05 07 1a 17 14 10 07 08 0c 06 05 08 07 06 06 0a 0b 0a 05 13 0b 15 14 11 1e 24 2c 46 4a 53 4f 4e 55 50 51 58 54 53 53 56 51 5a 53 5a 50 4c 52 52 4e 4d 4d 4a 4f 48 4f 50 43 42 3e 3d 39 36 35 3d 3a 37 3d 3f 3d 40 35 3e 41 39 37 34 2e 29 34 2f 25 33 32 32 2f 32 35 2d 2e 2c 2d 2f 2f 38 2f 31 31 2e 2c 33 47 35 3a 3a 45 42 3f 45 46 4c 49 4a 4d 57 55 63 53 49 51 48 4d 4d 49 41 2d 18 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 06 07 13 16 1d 1b 24 25 31 3d 3c 45 46 49 58 51 56 4c 4f 49 49 51 4f 4c 4c 3d 46 49 56 47 52 50 4d 48 46 51 4c 4a 4b 4d 4b 4e 4a 41 4f
 51 43 49 49 4a 4f 44 48 50 4f 54 57 50 4e 54 4b 53 54 4f 5c 53 51 5b 50 60 5d 59 5e 59 63 67 61 62 5d 62 5d 55 58 57 5a 57 53 51 52 55 4d 53 50 52 54 55 52 5b 63 5c 60 53 5c 55 56 49 50 4b 4a 50 50 49 3e 45 45 44 44 2f 15 06 05 08 05 0c 0f 10 14 09 14 03 06 06 05 07 05 06 05 03 01 09 05 0b 0a 0d 09 1a 15 1a 24 38 52 43 4d 3c 42 4a 48 4a 4e 53 51 4e 53 55 53 52 56 55 4c 4e 4b 4d 51 4a 46 41 42 45 41 45 40 38 3b 43 3d 40 33 3b 39 3d 36 3a 3c 2f 39 33 3f 34 32 33 2d 36 2b 34 35 32 30 31 2f 30 31 2d 2c 31 33 2e 37 31 33 2a 2d 3b 3d 41 41 40 44 3c 3f 3e 41 4a 5b 56 55 5d 58 56 50 44 50 4b 4a 3e 43 35 1e 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 0b 19 1e 1d 1b 22 2b 30 33 3b 3e 46 49 4c 50 50 4c 4a 4f 4c 4d 50 50 4f 4c 49 48 47 42 4d 49 48 47 40 41 51 44 45 4a 46 46 45 4b 4c 48 4d 46 47 41 45 44 4a 47 49 40 51 4e 49 49 4e 4a 51 4e 53 48 4e 57 61 5e 5b 5d 59 56 52 5f 5e 5b 60 54 52 57 50 4d 4f 51 4d 4f 4f 4a 58 57 4f 4f 4b 52 56 5b 5b 5e 51 4e 4c 51 53 4d 51 45 49 47 4b 4a 42 43 3b 48 3f 32 1b 06 05 08 00 06 05 0b 0e 10 05 03 07 0b 06 07 00 06 05 04 08 06 0a 03 05 13 14 0f 18 14 1a 31 3d 48 4c 46 43 50 44 4c 4e 4a 4a 4a 4e 4c 4e 58 4f 50 4a 48 51 47 4f 4c 44 42 4a 3e 48 3d 38 3d 38 3c 3a 36 3a 3a 3c 3b 30 2e 3d 30 30 2e 39 36 2e 3b 3b 30 3a 36 34 32 32 30 2b 33 33 33 32 30 26 26 33 2c 31 32 34 35 37 31 3e 3a 44 46 44 4c 4e 59 64 5c 5d 58 4f 4e 4a 4a 4f 4a 41 39 37 25 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 19 19 23 22 22 29 37 35 43 3c 3a 4e 4a 4b 50 4b 4a 4d 53 50 4d 41 4a 48 47 49 47 49 43 53 44 48 4d 4a 46 46 50 4c 4b 51 41 4f 4d 4c 4a 4a 48 46 4a 46 48 4d 47 50 46 45 49 50 49 45 4c 50 53 4d 50 54 57 52 52 55 52 5a 5a 60 5e 60 5f 54 55 50 54 57 53 57 4b 4e 4a 49 4f 4e 4c 45 49 4e 57 52 62 53 4d 51 47 47 43 52 45 4e 46 40 40 41 47 3d 44 3c 3e 39 1e 06 05 03 05 06 09 08 0a 06 05 03 00 06 05 03 02 0a 05 07 06 06 09 09 04 0c 0b 11 04 17 18 30 36 40 46 38 45 49 46 3b 41 45 4b 4a 4b 4f 46 4e 56 4e 4e 42 52 4a 4b 4b 4b 44 46 46 41 3f 37 39 3d 42 3c 2c 42 3b 37 3b 35 32 40 34 2e 30 34 2c 2f 3a 34 32 39 32 38 3c 36 32 32 38 32 33 2f 2b 2f 28 23 35 39 34 35 38 3d 3d 3e 40 40 45 4a 55 50 61 58 5b 50 55 4d 4f 4d 50 4d 48 3d 3c 2d 1b 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 13 12 24 1b 24 26 33 2e 33 39 45 40 54 4f 49 52 51 4b 47 4e 4a 4a 48 43 46 42 3e 50 4b 4b 4a 3d 42 49 46 51 4b 4e 4c 46 4f 51 51
 52 4d 4b 4d 51 4d 47 4d 4d 4e 48 45 4d 50 4d 59 4e 4f 4b 50 52 4f 4b 50 55 56 4f 54 55 59 5e 55 58 53 50 5c 4d 56 4a 4e 51 4e 4e 4b 4b 49 4c 47 52 4d 52 54 57 54 48 49 4b 44 4e 4b 3a 49 45 44 48 44 45 40 3a 3a 3e 3f 2f 19 0b 05 07 07 07 0b 09 10 10 06 03 00 06 05 0d 02 06 05 03 01 06 06 07 03 09 05 05 0f 0d 19 28 3c 3b 43 37 3e 42 41 46 44 3f 4a 50 47 4a 4e 4c 4f 49 49 4b 52 3e 57 45 53 4b 4f 46 45 43 44 40 33 3a 3f 38 37 35 35 35 38 37 38 36 33 39 2e 37 32 2f 38 32 34 26 31 42 34 36 2e 39 39 33 2a 30 2b 32 2f 2a 30 35 2e 3b 43 34 41 45 45 50 4b 5a 5b 5f 52 52 4d 55 53 4c 4b 52 44 44 43 36 29 0e 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 15 21 1b 1e 2a 24 37 36 3a 40 44 47 43 48 4d 4b 47 47 4e 4a 45 42 49 4a 44 3d 3e 46 48 47 46 42 4b 4f 47 4a 4e 40 45 44 42 4c 49 51 49 4c 45 42 44 4b 50 40 4e 47 45 50 4b 4e 51 4b 53 4e 44 55 51 51 48 4f 54 4e 4e 50 52 51 5a 56 56 55 4d 56 50 46 52 4b 49 4f 51 48 4a 48 4c 47 56 4e 4b 4d 50 49 4b 42 47 40 47 3b 43 45 43 36 32 3e 3f 3d 3a 35 25 11 06 05 03 00 06 05 0c 10 06 05 06 00 06 05 03 09 06 05 03 04 06 05 03 02 06 05 09 02 06 12 26 2f 3b 43 36 3e 3e 41 39 44 44 4b 45 44 49 45 4c 52 4f 54 43 4d 48 52 53 50 4f 45 45 41 42 41 33 3b 36 37 3a 35 34 36 41 36 39 3d 33 33 32 2b 28 2d 35 38 30 29 28 2c 33 34 30 37 32 37 32 30 31 2b 32 2e 2b 2f 35 3b 3a 30 3e 3d 39 50 59 5a 62 58 54 4c 4a 4f 4f 44 54 48 4b 4b 40 3f 27 1b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0c 15 19 21 17 1f 29 27 38 41 46 47 42 50 4b 49 45 4c 4a 4f 50 44 48 41 4b 42 41 44 50 46 4a 48 47 4d 4c 48 49 4b 4c 47 4b 4a 4f 4b 51 49 43 46 49 4f 48 42 4c 3c 48 48 49 55 50 52 4d 51 4d 44 4a 4e 4d 4b 50 51 51 4d 51 55 5c 5e 5c 55 54 50 4d 56 4f 4b 4d 4a 4d 4d 47 3d 4b 4f 44 4f 4b 4b 43 42 45 48 48 45 49 41 47 36 40 34 3a 39 37 39 3d 42 37 2f 1e 10 05 03 00 06 08 0c 11 08 07 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 09 09 0d 20 2e 35 33 32 40 41 39 39 34 42 43 40 49 40 46 46 4d 4f 50 4a 4a 4b 5b 4a 51 49 53 46 45 3f 4e 45 40 43 31 3c 3a 39 3d 3b 3b 36 3c 3b 35 35 34 29 2c 27 2e 2a 2d 30 2c 2f 2b 32 39 33 39 32 32 34 26 31 27 30 2f 3e 35 37 3a 40 3b 4f 59 5d 61 50 50 45 46 4b 4c 4d 4d 4c 45 50 47 3d 2c 1a 09 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 06 16 1e 1e 2f 27 2a 35 3e 3e 46 47 4f 48 4d 4a 49 49 4f 4b 40 47 4f 47 45 4a 42 40 48 46 49 47 4e 47 4d 4f 50 49 50 4d 50 51
 52 48 4b 47 52 46 3e 49 43 49 4e 4d 4a 52 4b 42 50 4e 4e 4e 50 4c 51 47 53 54 5a 4e 50 51 4d 55 4e 50 50 54 4f 55 53 48 4a 47 49 48 4b 48 4b 49 4b 4a 4e 43 4d 43 47 47 44 45 45 3c 38 3c 3d 3b 32 39 31 3e 35 45 38 37 33 1f 06 05 05 00 06 06 15 16 0a 07 03 00 06 05 03 04 06 05 03 00 06 05 05 00 06 06 03 0a 06 05 20 38 30 31 32 36 38 33 39 38 41 44 45 46 4c 4c 4d 4e 48 50 4f 4c 4f 51 51 54 4f 45 4c 4a 47 49 4a 3e 39 44 3c 3e 3d 35 37 37 37 37 39 3a 37 30 27 2a 2e 2f 2e 33 29 2d 39 37 35 2c 2e 34 35 34 34 2d 31 2f 34 45 36 34 37 3d 42 4e 47 5c 5a 53 58 48 4d 43 4d 45 4e 49 47 4a 48 47 38 22 0d 06 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 14 1b 22 1d 2a 29 35 3a 3f 44 45 4c 47 41 50 4b 44 4f 4d 47 45 40 4b 41 42 45 4d 47 45 46 47 4d 4f 4b 4f 4c 50 46 49 49 54 4a 4b 4a 44 48 4b 43 50 47 4a 50 4d 48 3f 51 4a 48 46 48 4d 4f 44 4b 4b 4a 50 4b 4f 45 4f 5a 54 54 52 4a 4a 5f 56 57 4b 4b 4f 52 4e 48 42 48 48 4c 4a 46 47 45 3f 45 44 3f 3b 3c 34 35 35 3a 3d 3a 2d 35 32 32 2f 39 38 24 21 06 05 03 00 06 09 10 0d 10 09 03 05 07 05 03 02 06 05 06 00 06 05 03 00 06 05 03 06 06 0e 16 2f 2d 30 30 36 3a 32 3b 35 39 44 42 44 48 43 3f 4d 4b 4c 3e 57 48 55 4b 4b 44 40 38 3f 43 3f 42 46 47 43 3b 43 32 31 40 31 30 3b 33 33 31 31 34 26 2d 26 2c 30 32 2d 2a 31 31 34 2d 2f 31 35 35 35 31 2f 34 29 38 34 39 43 44 49 52 53 5c 52 4b 4b 49 4d 4a 4d 53 45 42 47 41 41 29 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 13 1e 1e 1a 26 2e 2f 35 34 3b 3b 4b 44 43 4d 3e 4b 46 48 42 41 45 40 46 4c 3b 45 44 44 4e 47 50 4d 4a 50 54 4e 52 53 54 4b 51 4a 42 49 42 45 47 45 4f 46 48 4b 46 4a 4b 4c 50 4d 50 41 4f 45 47 4e 4d 4b 4d 48 54 4b 53 52 48 56 57 53 51 55 47 43 47 48 4a 50 3e 42 43 44 3d 40 43 3d 3e 3b 42 3b 30 39 35 34 35 31 34 34 30 3a 2c 2b 34 37 30 2d 15 06 05 03 04 06 0a 06 07 08 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 15 26 27 2e 34 35 31 34 2f 3e 37 3d 3d 44 45 45 48 4b 4e 48 4b 4f 4f 4e 50 49 3e 41 35 45 3a 3c 3d 3b 3e 3e 3e 2f 30 35 35 37 30 32 2c 31 2d 26 34 22 2d 34 25 2e 28 2e 2a 2d 2a 2b 2e 35 2f 31 33 37 31 36 2e 2f 30 37 3c 44 48 52 45 4a 43 44 47 42 4c 47 49 4a 4b 45 45 3b 36 29 17 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 11 21 1e 27 22 2c 2e 2e 37 39 39 44 45 43 47 44 43 3b 42 40 3e 41 48 44 38 44 45 41 48 4a 48 4f 46 49 49 4a 41 4a 48 49
 43 4a 49 50 4c 49 45 46 45 46 41 46 4a 44 48 4d 53 56 51 53 4e 4f 56 45 55 49 4b 47 3f 44 43 48 49 3e 41 46 44 4a 40 43 4a 45 40 47 46 3c 3c 42 45 41 41 3b 37 34 3e 35 32 31 35 31 30 2a 29 24 32 2e 2a 2c 26 28 24 26 1f 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 1b 2f 35 38 38 36 2c 3d 38 45 45 3f 46 4a 44 4b 4e 45 50 4a 47 4c 47 4a 49 49 49 44 42 42 44 41 45 43 44 3f 34 42 37 3d 44 3e 3a 37 3c 39 41 39 3b 38 2e 32 32 25 31 29 26 2d 2e 33 2e 2e 36 33 35 31 32 30 32 25 2d 30 29 34 2e 29 31 33 38 34 2f 3b 38 34 3f 38 3e 3d 33 31 1e 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0f 1f 25 27 23 2d 2f 3b 3a 3e 3c 3f 43 4a 44 45 42 3d 38 3a 44 3e 38 41 41 43 48 44 3e 40 45 42 49 45 4b 44 49 47 44 47 4b 3e 49 46 47 43 45 44 3e 3c 3a 3d 4b 44 4c 4c 4b 4f 51 51 4f 50 4c 4d 4d 53 4a 3e 3b 46 47 3e 41 45 41 46 42 4d 46 4a 49 42 44 3d 43 45 43 45 3b 38 37 33 36 31 30 2b 31 34 2e 27 31 2a 2d 29 29 20 25 20 22 1d 25 1f 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 1a 30 39 34 3a 3b 3a 3b 3a 39 3c 3c 49 3d 43 4d 4d 49 44 41 4e 42 49 48 41 4a 44 44 48 45 3f 40 3f 3e 42 3f 3f 36 36 3d 3e 38 3a 3b 36 38 3c 32 38 29 2a 29 2d 25 32 23 2a 2d 2d 2e 2d 33 36 32 2f 2f 35 32 2c 30 34 2d 2e 30 35 30 2c 2f 2d 39 36 32 35 31 33 3c 36 34 2a 20 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 1e 15 18 27 25 2c 34 31 42 3a 3f 3b 3b 42 48 45 42 45 3a 3b 49 3e 3d 49 45 45 3f 40 3b 3b 48 4b 43 50 47 45 43 46 46 42 3e 44 47 48 39 49 40 55 3e 3e 45 4e 43 44 42 4b 49 51 53 4a 4e 4a 4d 4f 55 3c 48 42 4a 4b 40 41 42 4f 43 44 46 4a 52 47 41 47 42 47 3b 47 45 36 35 37 29 35 2d 32 32 2d 2c 2f 2d 26 2d 2a 29 29 22 24 20 1f 29 24 17 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 2e 31 27 39 31 30 3b 3d 3c 40 36 3c 43 45 4b 46 4a 4e 47 40 3e 47 41 49 4e 49 4e 4d 4f 44 52 3e 41 42 3a 39 32 35 34 38 3e 3e 2a 2b 30 27 33 26 32 2d 29 2d 30 2c 26 24 23 2e 2a 2c 30 2c 30 2b 2f 34 2b 2b 2a 26 30 30 2f 38 27 2f 2d 31 35 30 3b 3d 30 39 33 37 33 26 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 13 23 29 2a 28 33 37 40 37 39 3a 41 3c 43 46 45 44 42 3f 48 4b 45 42 49 42 46 49 43 48 48 48 48 4b 52 40 3e 3f 46
 41 47 45 44 43 46 45 51 44 43 4c 46 3e 42 45 49 48 4d 44 57 4d 52 4a 43 4d 4a 4a 4e 4a 4b 4e 4f 4c 49 3f 4b 41 4b 51 4a 4b 44 48 44 3c 44 3f 43 3c 3a 36 37 2d 3a 2f 2a 2c 27 31 29 2e 22 29 26 26 24 2c 25 30 26 21 27 23 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 24 25 2c 2d 36 37 31 35 36 3a 44 3c 3c 40 45 49 45 3e 4a 46 4e 41 44 45 43 44 4b 48 4b 4c 47 47 43 3c 3c 35 31 30 37 31 33 37 39 33 31 35 2b 2a 20 2f 28 23 22 24 2e 2f 2b 33 31 2d 2b 2e 27 29 34 34 36 2e 2e 2d 30 29 2e 31 30 2e 32 28 30 37 31 32 38 34 3a 2e 31 32 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0f 1a 1c 29 2d 2b 35 39 30 3b 3e 3b 35 40 4a 46 40 44 40 3e 3f 48 4d 44 4b 4d 42 43 40 4c 48 4f 46 4d 46 41 49 40 43 4a 45 43 42 3a 3c 4a 43 4a 43 49 42 45 49 43 4a 45 42 46 44 4b 4b 4a 4b 46 45 50 4f 4e 50 48 4e 4e 4d 53 52 48 49 4a 51 49 49 48 38 40 3d 38 3d 35 34 33 27 30 2f 33 21 2a 2f 29 2c 26 24 26 1e 29 27 23 23 24 29 2a 22 1f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 21 2e 2d 35 34 31 30 3c 33 41 40 43 42 44 4d 48 45 49 48 44 3d 44 46 49 48 44 44 4a 49 43 3f 41 3d 3c 34 30 2d 2d 2e 32 32 33 2c 29 35 2f 2c 29 2d 24 26 27 25 26 2f 27 2a 2a 2c 2e 26 2e 31 2c 32 2b 31 2d 30 30 2e 39 33 37 28 2a 33 34 2f 36 36 3a 2a 3c 3e 30 27 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 14 20 24 26 37 34 3d 35 3a 3f 39 44 3e 3a 40 3e 3c 45 3d 44 38 3c 47 43 53 4a 4a 43 47 42 41 48 42 47 43 47 3d 4b 3f 46 3e 39 3c 3e 3e 3f 46 3e 43 3e 37 4c 42 46 49 4c 42 4b 47 49 4b 4a 41 51 43 46 49 4d 46 48 54 52 5b 49 49 4f 4a 49 3e 38 35 38 3c 34 3b 2e 31 2e 2a 30 29 25 28 26 2c 2b 24 1d 22 26 26 26 25 25 23 23 2f 1f 23 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 1b 35 25 2e 2b 2b 34 33 38 3f 40 3a 43 3f 41 44 40 4d 45 46 42 40 49 3d 42 42 44 48 49 3f 40 3a 39 43 38 30 36 39 29 2f 35 35 2f 2e 2f 28 28 27 2f 28 23 24 24 29 27 29 31 2f 29 2c 3c 31 35 31 2f 2f 23 2a 2b 2a 30 2c 24 34 23 2a 36 35 34 32 31 3a 36 3b 36 24 22 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 16 21 25 25 32 3e 3b 3c 3d 42 38 3f 43 3a 43 3e 3e 45 3f 4a 38 42 42 44 4a 4b 41 41 4e 42 3e 44 42 53 4c 51
 3b 44 43 45 4b 4a 3e 44 47 41 49 43 43 45 47 46 46 3f 42 46 4a 48 45 52 53 4b 4a 47 4d 50 55 45 4b 4e 48 52 4c 4f 50 51 50 42 3f 36 3c 38 34 37 39 33 34 2f 2b 33 31 28 27 2e 28 25 24 2b 2d 2b 20 22 27 28 2b 27 2b 2e 2b 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 14 22 29 2a 30 35 35 36 36 40 40 45 41 3e 4c 41 47 46 46 41 43 42 4a 3f 42 3e 3c 4a 49 41 48 44 3a 3d 3c 34 2b 35 36 3e 39 37 34 31 2b 34 38 2e 2a 22 2a 28 25 24 2b 28 26 2d 28 2a 37 38 2e 31 36 26 34 31 35 2e 31 31 34 2b 35 2f 2f 39 34 36 38 36 3d 36 35 39 22 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0b 1e 2e 31 30 30 3e 3a 42 42 3b 3e 3c 3e 40 42 3f 32 37 3f 42 41 42 39 41 41 48 40 4d 42 49 49 4e 4c 41 45 47 41 44 4d 4d 49 4a 3f 3c 3c 44 45 3c 43 44 44 40 4b 3f 41 47 4c 4b 4d 4d 4e 4c 4d 4d 52 4b 50 49 43 46 50 54 58 4d 4a 43 43 40 3b 38 33 32 38 2d 32 38 31 2e 2e 2a 27 27 2c 32 27 28 28 24 2a 21 23 23 28 23 26 33 25 20 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 20 29 2e 30 39 2d 34 39 34 46 41 3d 3e 4c 49 4b 48 46 47 45 3e 40 41 45 3e 3c 47 49 45 4c 45 45 3e 42 34 35 2c 39 36 2d 30 37 31 25 2a 2c 27 25 31 30 2c 25 25 2c 25 27 35 34 35 39 42 3a 37 2d 30 35 24 30 2c 2d 32 39 35 3a 2c 35 2a 2e 3d 2f 30 35 37 36 27 15 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 16 23 2d 30 3d 3a 30 3a 3a 40 3a 35 3b 42 43 39 44 40 42 39 45 43 3b 3b 44 47 3e 3e 47 49 3f 43 42 3c 40 3d 40 43 40 47 54 46 4b 43 3e 3e 41 43 3e 45 44 43 45 42 3a 4a 4d 48 52 50 47 47 4e 51 50 51 4b 3a 42 4e 55 4a 4a 45 3f 46 42 3b 3a 36 27 35 37 2f 30 2e 30 2f 2b 2f 23 2a 21 25 24 27 23 26 22 28 28 26 2b 2b 2b 30 21 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 1e 20 2a 2f 30 34 36 34 41 37 42 45 41 44 48 48 4b 43 4b 40 42 4b 46 4a 41 44 43 36 47 44 3a 3e 3c 35 2d 31 2e 2e 2f 2e 2f 2e 30 30 2e 23 2e 2e 2e 24 2a 2f 23 33 31 30 35 48 4a 45 41 35 37 2f 2f 2f 28 2f 31 34 31 2f 2f 2f 36 2f 37 32 32 34 36 3d 34 2b 20 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 17 1d 2d 36 35 34 41 3a 3d 3f 35 37 3e 3b 42 3e 41 42 3d 3c 34 39 3b 3c 44 48 41 43 43 48 3e 45 45
 3c 43 48 36 41 41 4a 4c 46 3d 44 43 46 41 3d 41 40 41 44 45 3f 43 48 42 49 44 47 43 49 48 53 3a 23 31 50 54 51 4b 40 44 43 45 3e 35 2d 2e 2c 30 38 2f 36 2e 27 27 2a 25 2e 24 23 24 2a 2e 1e 23 2c 25 29 2a 26 31 27 35 2a 1f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 22 2b 2e 29 35 31 33 38 37 41 39 42 48 48 3e 50 54 46 46 49 45 45 3d 44 47 3e 3f 41 39 3a 40 36 3f 34 2c 25 26 32 36 2b 29 36 2c 2d 32 2f 30 31 30 2d 2c 27 29 31 28 2f 3e 46 4a 3c 39 33 2e 2b 35 30 31 30 35 3b 2e 28 34 31 31 33 36 32 36 34 38 3d 37 24 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 11 22 24 2e 3c 32 39 3b 3a 3e 3f 39 41 39 3b 40 40 40 43 3a 41 40 43 40 42 43 43 3e 40 44 3f 44 3e 3d 41 40 43 41 43 43 46 42 43 47 40 4a 41 38 41 44 39 45 41 46 47 43 3d 4c 42 41 4d 41 4a 43 43 48 4e 55 4d 48 49 47 44 48 3d 39 3a 31 30 30 2b 2b 2a 2a 31 35 31 2e 34 28 2c 2a 28 21 27 26 28 2a 2a 2d 2f 28 2b 32 2e 30 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 1a 26 25 30 35 29 38 39 39 41 3e 49 49 43 47 45 49 46 48 4b 4d 45 49 4a 44 3c 3a 44 49 40 32 37 39 35 33 32 38 39 32 30 32 2a 26 33 34 31 2c 31 2a 3d 2c 29 31 39 28 32 3d 3f 42 39 3c 38 2e 2f 2a 3a 28 34 24 35 30 33 3b 37 34 36 39 30 35 37 3d 34 25 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 25 2a 33 30 3b 39 3a 43 43 3a 41 3e 34 3d 3d 41 40 42 42 40 39 42 3d 40 35 41 41 3d 43 3c 3f 3d 3a 3e 3a 40 48 3d 41 43 3d 3b 38 44 49 3b 3f 44 43 42 3e 43 46 3e 44 48 4a 43 47 41 3d 4c 45 41 42 47 4f 3f 42 43 3c 46 41 3a 39 2d 33 30 33 37 30 2c 2a 30 2e 26 2e 24 25 27 22 29 2d 1f 2b 2c 2a 31 27 23 2e 28 2d 26 1f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 30 26 30 2c 35 33 3a 3a 45 3b 46 40 43 47 4b 50 4e 4b 4f 3e 4d 4c 4a 44 40 34 3a 37 3a 38 31 39 2e 33 2e 2f 2b 33 39 2c 31 27 33 37 36 33 33 31 34 2d 29 2b 34 27 2f 2e 36 32 3c 2f 37 29 33 34 2e 30 32 30 31 31 36 36 38 2f 33 34 35 37 2f 36 31 17 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 2a 22 29 2a 38 35 3a 3e 39 3f 39 38 36 3f 38 40 39 3f 36 34 3d 3f 44 3e 43 3e 3a 3d 36 44 42
 39 3e 47 38 42 3a 40 3d 3d 42 3e 3e 38 45 44 44 3c 3d 41 4c 39 3e 37 3d 44 4a 3f 3b 42 38 40 41 42 3d 42 48 3e 3e 3e 40 38 3d 41 3d 33 30 27 2e 31 34 32 33 2a 2f 25 2a 2c 24 29 2e 2b 27 2d 25 28 26 22 2f 30 26 3c 2c 2a 2b 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 1a 25 24 30 32 38 38 3b 37 3b 44 46 45 44 4b 4f 53 4d 4b 46 3f 44 49 46 3e 3f 3c 3f 3b 38 35 37 35 31 2e 2e 32 2f 26 33 35 35 33 37 34 31 32 36 2c 2d 36 32 36 2e 2f 32 32 35 2e 2c 35 37 31 2f 34 35 29 36 31 34 35 39 3a 3e 3a 31 35 30 3b 35 34 23 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 20 2a 32 39 36 35 3e 38 3d 35 3b 3e 37 35 3e 3a 3a 39 37 42 3c 42 38 40 3d 3c 41 38 42 43 40 39 41 3b 3d 3a 3e 45 40 3e 3e 45 3e 41 3f 43 3f 46 3c 43 42 3f 41 41 42 38 43 49 40 40 40 3e 40 3f 4d 42 3b 46 40 47 48 38 3b 38 32 2f 39 2c 26 24 30 33 34 30 2f 2b 2c 26 28 2c 21 27 2c 2c 29 30 26 2e 2f 2a 2c 31 27 22 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 10 26 29 34 2b 3e 36 3a 3e 51 43 3f 47 49 44 4d 4c 4f 51 51 4d 4e 41 47 45 3e 3d 37 33 34 36 38 30 30 32 29 33 2f 2f 3a 30 31 33 39 2d 34 36 30 3b 2e 2b 31 2e 30 26 2f 32 32 30 33 36 30 37 36 3b 39 30 39 2f 38 33 39 34 35 37 3b 3a 3c 3b 33 24 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 19 2d 2f 35 38 39 34 2f 39 30 39 40 39 3f 3a 41 37 40 38 3e 39 3e 3b 40 41 3d 40 38 46 43 36 39 3f 3c 40 42 43 37 40 45 40 40 41 3d 3b 42 3b 4a 44 41 46 43 40 3f 46 49 4d 3a 33 39 39 40 3f 3c 3b 3a 3b 3c 3a 47 36 31 35 34 39 35 35 2c 31 33 2b 27 26 28 23 26 29 2e 35 2c 2f 25 2f 2c 2c 22 31 2f 2d 33 2e 24 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0f 23 2a 39 2f 33 36 36 3c 42 42 43 41 4f 47 4f 52 54 50 52 49 44 3a 42 31 3c 40 39 3c 39 2d 3b 32 2b 34 31 36 36 35 33 2f 37 37 31 3a 34 2a 2e 2f 36 26 2b 28 32 2c 2b 2e 2d 2c 32 2e 34 31 31 32 3d 34 36 39 32 3d 38 32 3f 32 39 35 3a 38 29 11 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 1f 2a 33 39 36 34 3a 41 35 3d 35 38 3b 39 3b 3d 3b 32 40 37 46 38 3b 3d 3d 39 38 38
 3a 3e 42 34 3f 3b 3a 3b 40 3d 3f 40 38 3c 3d 3e 4d 40 3c 45 42 42 47 40 4b 3b 39 3c 3b 39 39 39 45 39 3c 40 40 36 3b 41 3e 33 3e 30 2e 36 2b 36 31 29 30 32 35 2b 2d 2b 30 24 24 29 2c 2f 26 2d 2b 30 2f 2b 23 1f 24 25 26 1f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 2c 26 3a 3d 3b 35 3b 3f 43 4e 46 4c 4a 4b 5d 4f 53 4d 49 45 44 40 3b 3c 34 3d 34 2d 32 34 3a 3c 37 27 30 3d 30 33 32 27 36 33 2a 36 2c 34 30 32 35 29 34 30 33 31 32 37 30 2e 2f 2f 31 36 3d 2b 36 34 35 35 34 31 34 45 3e 3b 34 3a 31 2b 1a 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0c 26 22 2d 36 3d 31 34 3b 44 35 3c 38 45 35 35 3e 34 3e 3d 45 42 42 41 3e 3c 3b 37 3f 42 3e 43 3f 3f 3e 3e 39 3b 3f 3a 3b 44 3d 40 3d 3a 42 45 3f 49 4b 42 41 3b 3e 3d 40 36 3b 37 3c 38 37 3b 3a 3a 39 3e 3b 34 37 3b 34 33 34 3d 32 36 2d 32 2a 3a 2c 2b 26 2d 2a 2e 2f 30 2e 2e 27 22 27 2b 30 25 26 25 1c 1f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 17 28 2b 2f 33 36 3d 40 43 40 46 50 4d 52 4c 5a 55 5a 44 41 47 44 3a 3f 3c 3f 3a 32 39 38 37 39 35 3e 2f 3b 30 38 3a 34 36 33 3b 32 30 32 38 30 36 2f 2d 34 28 39 32 2f 3f 31 28 2e 30 42 40 3d 37 36 2e 39 36 37 3d 37 3a 3f 39 38 3e 30 19 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 17 21 27 35 30 31 3b 3b 3b 39 32 3e 3d 3a 3c 35 3f 3e 41 41 3b 44 3e 3c 3d 43 36 37 49 3f 42 42 41 3d 3d 42 3e 3c 44 44 42 3c 43 3d 39 3c 3b 38 41 3f 45 3e 3a 45 3d 3b 3c 36 3b 41 3e 41 42 44 36 35 35 36 30 3b 32 34 2f 30 31 2d 31 34 31 2e 31 27 2f 29 26 29 29 2c 2b 2d 2d 2a 27 27 21 23 25 2f 2b 25 20 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 32 31 35 3a 3c 43 38 40 45 44 50 51 54 49 54 50 53 4c 3d 47 40 39 37 35 3f 31 3f 36 3f 38 3b 39 35 39 35 2a 34 33 36 35 36 2e 28 38 35 35 39 33 2e 33 34 35 34 33 2a 29 34 31 41 31 3a 39 38 34 3d 34 2e 31 35 45 38 3d 44 39 2f 2a 16 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 1b 1f 2d 33 2d 36 35 3a 3b 3d 32 41 35 39 37 3f 3f 3b 41 3b 42 42 40 3d 37 3d
 45 41 3c 3f 3b 44 3b 3e 39 37 40 44 38 3a 3f 47 3b 3f 3f 43 38 43 3e 40 41 3b 3c 42 3f 39 38 3a 37 3d 39 3b 38 35 3a 38 34 32 36 31 2e 2c 2c 32 31 29 2f 2c 29 2d 34 2a 28 28 2d 2f 29 30 1f 28 22 27 2a 24 1e 26 20 27 26 19 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 18 2d 33 34 3a 3f 3b 47 3c 51 3f 4d 4f 4c 4e 4c 4e 4c 47 4b 3f 39 3a 3b 35 34 30 31 3d 33 34 33 34 2f 38 2f 31 36 31 2f 30 30 32 2e 33 35 33 2f 2b 2d 2a 37 32 34 3d 35 36 3a 2e 2f 2d 34 37 3b 38 39 38 35 33 40 3f 37 3e 35 33 2f 1d 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 16 26 2b 2e 31 3b 3a 3b 3d 3a 3c 35 38 3d 3e 3e 40 3a 37 40 40 3d 3e 3e 47 3c 38 3c 39 38 3f 3c 3c 3e 44 3f 37 34 40 44 42 42 37 3e 49 3d 3a 45 3d 3b 41 3d 44 3d 3d 3a 44 3d 3c 36 35 3a 38 37 3a 39 31 35 2e 2c 34 23 31 2e 28 27 2e 2e 2e 2e 26 20 28 21 2c 29 2b 29 28 29 2b 26 29 24 27 26 24 21 1f 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1c 35 30 32 3b 3b 40 44 44 47 46 4c 45 4e 50 50 56 47 47 49 42 44 3d 4b 31 36 38 39 3d 3c 35 31 36 2e 32 35 39 39 37 3b 2a 37 33 35 3d 37 35 3b 3a 3f 35 35 35 3d 3b 2e 35 35 31 3a 33 3b 3d 40 37 44 37 36 3e 35 32 3f 3a 3b 28 25 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 1b 1f 26 32 2a 36 34 3d 35 32 3c 3c 35 36 3d 41 38 3f 3e 3c 3e 39 39 44 46 47 36 3a 3f 40 3d 3a 3c 42 39 43 42 41 42 43 43 41 3f 44 39 41 42 3b 3f 3c 3a 43 3f 46 43 40 3c 3d 3e 35 36 33 36 3c 37 2f 34 35 31 36 24 2d 2c 27 26 29 1c 2f 25 2a 22 28 26 26 2d 23 21 1c 24 20 24 26 25 27 22 2b 28 25 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 15 2a 2d 31 3d 40 3b 3f 3d 4b 46 4b 4d 4b 4d 4c 4e 50 41 3f 44 40 3a 43 3b 3c 36 3e 35 3e 2f 3a 38 30 33 30 30 3b 34 3b 3d 36 38 33 3c 3a 30 37 39 3a 39 38 38 32 3c 36 38 36 30 40 3a 35 3e 3b 32 3d 3b 3c 38 40 3a 36 3a 32 1b 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 07 11 24 2d 2f 30 38 36 37 39 37 3b 2e 32 35 3c 38 37 39 41 3f 3c 3d 38
 33 3e 35 38 36 3a 3b 3e 3f 47 3e 3c 3f 3e 3c 3c 39 37 47 44 3d 40 42 3b 36 3a 32 3b 36 3e 37 3c 39 36 37 39 35 3d 36 3e 34 31 32 33 2c 2e 2a 2c 27 22 27 21 25 24 1f 20 23 23 2a 23 27 2a 2a 1f 24 1d 2c 1b 1f 24 25 1f 1d 20 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 29 24 31 31 3b 3d 3b 43 47 4f 4d 45 4f 51 4c 46 41 3c 3e 3d 3a 3f 3e 31 42 39 36 33 38 35 34 36 35 31 32 39 33 35 35 3b 38 36 35 30 45 35 32 39 3c 34 36 35 3b 3f 38 36 30 33 2f 39 39 38 39 35 38 30 36 39 38 35 2d 29 28 0e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 15 1b 2a 2b 37 2e 34 39 3a 38 3f 33 37 3d 3b 3a 41 42 37 38 39 32 3b 3c 35 36 36 39 40 38 40 36 3b 3a 39 3d 3c 39 3b 3c 42 41 42 3d 40 3a 3d 3a 40 3c 3a 3e 3f 35 3e 3e 3e 40 2f 39 3a 3a 39 34 39 35 2a 2d 36 2e 34 25 2a 2a 27 22 21 1b 22 2f 2a 2a 2d 25 22 25 1f 1c 27 24 27 2b 26 25 1b 20 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 15 25 25 2b 3f 36 3c 42 45 44 49 43 44 4c 44 43 42 3f 3c 3e 34 3b 38 37 3d 30 3a 35 40 3b 2f 35 31 3d 30 2f 3b 35 38 35 3e 3f 42 3d 39 3a 3a 38 37 37 37 43 3b 3e 37 30 3a 35 33 3a 36 35 3e 41 3b 3c 32 37 3b 37 33 31 1d 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0e 21 2a 2f 42 3a 3e 3c 35 34 38 37 41 38 37 44 39 41 41 37 3b 37 40 35 40 39 3a 3a 3b 40 49 36 3c 39 3c 40 44 41 3c 3e 3b 39 42 3b 3b 3f 3d 43 3b 3c 35 39 43 3a 3b 44 37 3e 36 33 34 36 40 34 39 2d 2f 32 2b 2d 31 26 28 29 2e 25 25 23 1e 2b 22 23 27 21 2b 24 25 25 23 23 26 22 25 1a 1f 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 12 23 25 30 2f 37 3b 3f 3d 3b 35 47 3c 44 41 46 43 45 3d 40 3b 3f 36 3f 39 39 3e 3a 3b 35 3c 3f 34 3a 39 3b 44 39 36 3d 38 3b 38 37 3b 3d 3a 37 36 3b 31 37 3d 39 34 31 39 37 3b 42 3a 38 37 48 40 3e 38 38 31 30 29 1f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 11 1d 30 30 2c 31 31 3b 32 37 31 36 3d 37 3a 34 3b 33 32 39 39
 40 37 3f 38 3d 3d 36 3b 37 32 3f 41 3b 39 38 3a 48 36 44 3f 41 36 3a 42 3b 41 40 3a 38 38 38 37 3c 33 39 3a 35 36 35 34 34 3d 3d 34 31 2a 2a 2d 28 25 28 25 26 2e 22 21 1f 22 1b 2e 29 25 1d 23 25 26 25 25 2b 23 20 27 28 21 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 2b 33 34 31 38 38 39 31 3f 41 36 40 3c 42 42 3a 3b 35 41 42 3a 40 40 3a 35 38 3a 37 3e 35 33 42 41 3c 36 3e 3e 3f 32 3e 3b 36 3c 3d 38 3b 41 35 37 38 38 30 3e 34 3f 3b 37 3f 3e 38 39 2d 38 3c 36 35 39 37 30 20 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 18 27 29 36 3f 38 39 32 3a 3a 3d 36 3a 41 3a 41 3e 37 36 3c 35 3e 3a 36 38 3b 36 34 41 39 34 3e 3f 3d 3d 3e 40 42 3c 37 44 3e 40 41 39 42 45 37 3a 44 3c 40 3a 3d 3c 3a 35 41 40 34 34 39 32 37 34 30 35 2d 30 30 26 2c 2f 24 29 2b 2a 26 2d 27 29 2c 24 2a 25 25 21 20 26 30 26 24 1a 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 1f 25 35 35 33 36 34 39 3d 42 44 39 43 41 3b 3e 3c 3e 45 3c 43 3e 43 3b 3b 3b 42 3f 3a 37 4b 4a 3f 43 3b 47 44 41 44 36 3b 3f 38 3c 42 3d 3b 3b 36 3a 41 3b 41 37 31 43 42 3f 39 35 37 47 3b 36 35 38 34 2e 25 0c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 1a 21 2c 35 31 32 32 36 36 36 3e 3e 36 39 37 3b 3a 3a 3c 3d 37 3e 37 3e 35 3b 33 3c 3d 38 3b 41 37 46 39 38 3b 49 34 34 49 3e 43 4c 38 47 3f 3b 36 3c 45 38 45 40 36 38 36 3a 3e 38 3b 37 31 32 30 3a 2e 30 32 25 2d 2f 28 23 2a 29 2a 33 26 35 2c 25 24 22 25 1d 23 1e 2c 25 27 1b 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 24 2b 30 3b 35 38 36 38 39 38 3e 3f 44 3f 3c 39 41 38 44 3e 43 41 3f 41 3c 46 45 41 45 41 49 51 47 3b 35 40 3d 3d 3e 3b 38 46 42 40 41 3b 34 3e 3e 2d 46 3a 3f 40 35 39 40 39 38 3a 3c 3d 38 39 33 36 2a 20 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 1f 30 27 3b 36 3b 36 31 3a 35 35 33 31 31 38 3c 38
 3f 34 37 35 3e 3c 39 32 37 39 3a 3b 39 3c 41 40 3d 3b 3b 3d 32 47 3d 3f 3c 40 44 3f 3f 3b 45 3d 34 3d 3b 39 42 39 38 3d 39 3b 39 3d 35 2f 37 39 36 2b 2e 31 29 2b 2a 2a 2b 26 28 29 29 2e 26 25 24 22 23 26 2b 24 2a 25 20 20 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 28 2c 30 3f 31 33 3e 34 39 3f 3b 45 3f 3c 3e 40 42 32 3b 41 46 37 44 3e 3a 3f 3b 3c 40 3d 40 41 43 44 3e 40 45 3d 49 44 41 3c 44 47 42 44 39 3a 41 3a 39 40 41 40 38 3f 37 33 3e 3b 35 37 34 3e 32 26 1f 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 21 31 31 37 30 36 35 37 38 3a 39 3b 39 36 32 37 3e 3e 3b 2f 33 36 36 39 38 36 3a 32 3b 37 3e 3f 3b 3b 33 42 38 45 3c 37 38 39 38 3e 3b 3e 36 40 3d 39 3f 39 3f 3f 3e 3d 3c 30 41 32 3d 3e 38 36 35 32 2d 30 30 25 2b 28 30 2e 2d 2c 29 2a 2b 25 26 21 32 31 2b 25 29 24 26 1a 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 2a 23 2e 32 35 39 37 36 44 3b 3b 34 3d 3f 3f 37 40 3f 45 3d 43 3d 41 3f 44 42 45 41 47 3e 3e 49 44 45 3d 44 3f 3e 40 40 45 3b 3b 3f 3e 44 3b 3c 41 3b 36 3b 3e 3e 37 3f 37 36 3a 39 35 43 3d 35 2a 20 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 13 1f 2d 33 32 32 37 36 37 39 3e 38 35 38 3f 3b 3a 37 40 3d 36 33 36 37 38 38 37 39 41 35 3a 3e 43 39 3e 39 3e 3b 3e 3c 38 41 38 42 3b 3b 3e 3e 43 39 3b 41 41 39 3a 3c 40 40 3a 38 40 34 2f 39 38 38 30 33 34 2f 28 2b 33 2f 2f 31 28 2f 29 25 28 2a 27 26 23 29 23 26 2a 21 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 28 30 2d 2f 37 3c 36 3d 36 35 3f 42 49 3d 44 45 3c 3d 3d 48 49 47 43 42 40 43 46 45 41 3f 4a 44 3c 44 3e 44 46 42 47 41 3b 44 3b 4a 41 41 38 3c 39 3c 42 44 44 45 38 3c 38 3f 3d 41 35 3a 2c 1f 0e 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0d 20 30 2c 32 32 32 36 42 3d 36 40 36 36 3c
 41 38 3d 3f 34 38 3c 36 3d 3d 3d 39 3b 37 36 3e 42 3d 37 41 3d 40 35 33 45 3d 3f 3b 37 42 3d 3d 40 40 39 3e 38 3e 39 3d 43 33 33 35 32 34 35 3b 30 3b 35 2f 3b 2d 34 3c 32 32 2c 2f 35 30 2d 2a 2a 2f 2d 2e 2e 21 2d 28 21 21 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 25 33 34 3c 39 33 3c 37 3f 35 3a 3c 3f 44 3f 46 40 43 48 40 43 42 4b 48 41 48 41 44 42 3e 3c 3a 3d 46 4a 3f 46 42 3e 41 3e 44 42 40 44 3b 44 3c 39 38 3f 36 41 3a 34 3b 35 39 38 3f 38 36 2b 16 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 18 1f 25 29 2f 37 3d 39 34 42 31 30 3e 2f 3b 39 35 35 3b 30 3a 3a 35 3a 36 40 32 3e 3e 41 37 3e 41 3b 3a 3b 3f 3b 3d 3d 32 3b 38 3d 3f 3f 3f 3c 3f 3d 3b 3b 3a 3a 3b 34 41 3b 3a 42 37 3b 32 32 30 32 35 35 34 32 35 2e 35 35 2d 2c 30 29 32 26 2d 25 29 27 28 25 1d 25 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 2d 32 39 39 34 36 3e 37 3f 3e 49 41 3d 40 3c 42 49 49 3f 41 44 46 42 41 43 4b 42 3d 43 41 4a 43 41 3b 42 46 42 42 4a 47 44 39 3e 39 37 43 42 42 41 3e 3c 45 37 3c 36 38 38 3d 37 33 2b 20 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 15 22 23 34 33 32 3a 38 3f 3c 3d 36 3a 37 3e 3e 3c 3a 3b 3c 39 37 3c 3e 3f 35 45 3c 44 3e 36 43 3f 36 3e 3b 38 43 38 3c 44 32 3d 42 3f 44 46 40 3a 3a 33 41 3c 3b 3b 3c 35 32 41 3e 39 3f 3b 35 3c 2d 37 38 2e 32 38 3c 33 32 39 35 32 32 35 35 33 2e 25 2c 2d 27 2c 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 29 29 38 39 35 3c 36 47 45 43 3e 37 38 45 3b 46 48 3f 42 3c 40 45 48 4b 43 44 44 43 43 45 40 40 3c 3f 42 4b 46 4b 41 3f 42 40 40 45 40 3c 41 42 39 40 3e 3d 3d 37 37 3a 3e 37 3b 31 24 18 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 12 1b 26 28 3e 32 33 38 35 2f 34 40
 37 3e 2f 35 34 3a 31 3b 3c 35 3c 39 3d 42 41 35 36 3e 37 38 3f 3c 3f 3a 3a 36 35 3d 3c 3e 41 42 38 44 42 40 37 3b 3e 38 3b 32 3e 34 38 3d 38 37 3a 36 37 3b 38 38 38 34 39 30 39 31 2b 34 34 33 33 2f 2a 33 2e 28 2e 2b 29 23 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2f 33 3c 39 39 41 3b 40 37 40 3d 39 41 42 48 3d 3c 3f 44 41 47 4e 3c 46 43 4b 44 41 48 3c 46 43 39 3f 4c 40 4a 43 40 40 4b 40 3e 40 44 3f 41 39 41 3a 34 3c 38 41 3b 3e 31 31 31 24 12 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 14 17 25 35 30 30 36 32 3e 37 30 3c 3b 3c 3c 36 40 34 39 3a 36 36 36 3b 3f 37 35 33 32 33 3d 3c 3c 3e 2d 39 39 39 39 3a 39 38 41 40 3f 45 42 3a 3c 41 3a 3c 40 46 3d 39 38 3c 3c 33 36 38 3d 3b 3f 3c 34 3a 32 37 39 3b 2f 32 33 34 30 30 26 2f 23 2b 31 32 2a 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2a 36 3f 42 3b 33 3d 46 3c 42 3d 38 42 3a 4b 3d 44 40 3f 49 48 46 4b 3c 42 42 40 38 44 47 43 3f 3f 45 43 42 3e 40 43 3e 45 41 3c 3f 3e 40 3e 40 43 39 37 33 3e 3c 3e 3a 36 29 1d 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 17 1a 27 33 31 3c 33 34 3a 37 43 3f 3a 39 36 3e 3f 3c 37 39 35 3b 38 41 3a 35 3c 34 3c 3b 37 3b 39 38 3d 45 33 3d 3d 37 3e 3d 3a 3a 3b 44 3b 37 38 3c 3c 3b 35 34 44 39 3f 41 43 3a 3a 39 3c 3d 3c 35 38 32 44 3e 3c 33 30 35 2e 33 32 30 29 2e 30 2b 29 29 1e 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 29 33 3a 3c 34 39 3e 39 40 3d 41 4a 3f 42 44 3a 43 42 41 4b 43 49 47 40 44 4b 49 4e 4c 48 3f 49 48 45 3e 41 3f 44 44 3f 43 43 3e 47 3d 3f 3c 41 3b 3e 36 36 3c 3f 35 39 2f 26 1f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0d 19 25 29 30 2f 37 3b 33 44
 3d 44 35 35 34 42 39 40 3a 3e 2f 37 32 3c 3f 33 3b 3b 38 44 3e 35 38 3b 3d 35 3a 3a 34 3e 3a 44 48 3c 44 44 3b 49 3f 40 3f 3c 36 40 44 3d 33 35 3c 38 3c 3b 37 3a 38 2e 3f 30 35 38 3a 3e 38 34 2b 34 33 32 31 2d 2a 28 2f 2b 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2e 33 3e 3f 41 42 3b 42 44 3e 3e 3d 3f 42 48 43 4d 41 4b 40 40 3b 49 3b 3a 43 41 45 41 43 44 4b 46 44 41 40 47 39 3e 47 2e 4a 44 39 44 39 3a 39 43 3a 3d 3b 3c 33 32 31 26 10 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0d 20 28 33 34 31 34 37 3e 35 33 39 35 3c 37 33 3a 3a 3a 40 37 34 3a 36 40 3e 38 3b 41 39 3a 2c 37 36 3d 3c 35 37 3a 37 3c 3a 3d 45 41 3a 36 3a 3c 3f 37 3a 3e 38 36 3f 3f 3d 31 3b 33 38 35 2f 37 3e 3e 40 39 32 35 33 34 2f 32 34 33 29 29 29 29 2c 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 2f 39 3d 33 39 39 3f 42 3e 3f 41 45 45 42 43 3b 3e 42 42 3f 42 44 42 46 39 46 43 48 3d 42 47 3d 41 4b 3e 41 46 3f 45 48 38 3c 3d 3a 34 3d 36 3c 3e 39 35 3a 2f 27 25 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 1d 20 27 32 30 39 39 35 38 3d 36 36 44 39 3f 39 3f 3b 3a 34 3b 35 3b 41 41 39 37 3a 40 3c 3a 34 38 3a 32 39 3d 41 35 39 3b 3c 42 3e 3d 42 3c 39 3a 30 42 40 36 35 39 3e 36 39 3b 3d 3d 36 3c 34 39 36 37 31 3b 36 36 32 2d 2e 39 2d 2e 38 37 32 29 24 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 26 35 32 41 35 44 3a 35 44 3d 42 44 42 44 3d 45 44 3f 48 3d 47 3e 45 39 3f 3e 46 41 46 4c 49 4a 44 40 44 46 3e 41 39 43 3f 3a 41 3d 45 42 38 43 3e 3b 40 31 2c 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 11 1a 2a 36 34 3e 36
 38 3c 3a 36 37 3d 35 39 37 3d 39 41 3f 36 35 38 3d 38 37 3e 34 39 3d 38 40 33 36 36 39 3f 43 41 3b 3d 3b 46 3a 3b 39 41 3a 35 3a 3f 41 43 34 3b 3c 3b 36 40 40 37 3d 3e 38 36 45 37 3c 3c 3c 34 33 36 2c 31 2a 38 30 34 23 30 25 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 39 38 40 36 3b 3e 3b 3f 42 44 3d 41 3f 3f 42 45 41 43 40 44 3f 41 47 36 44 4c 48 47 45 47 47 3f 4b 48 42 3f 3b 43 3e 48 41 45 40 39 40 3f 3b 3a 36 32 28 1a 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 18 24 30 34 34 3d 37 3f 35 3b 36 31 3d 40 3c 36 42 33 32 38 39 35 35 39 43 33 38 3b 2e 37 32 35 2f 35 31 35 3d 42 35 35 3e 37 35 3d 3b 3c 32 41 37 39 3f 33 40 3b 3a 30 34 3a 3a 39 39 3f 38 39 39 3a 38 37 42 36 36 2c 35 34 31 33 36 2f 2b 29 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 24 34 3f 48 40 33 3e 3a 3c 3e 3f 3e 3a 44 40 3d 44 46 45 42 42 44 41 3a 43 3c 3e 44 3c 48 47 43 46 3e 40 48 47 44 3f 3e 42 42 3a 3c 37 40 38 35 2d 29 1d 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 18 15 2f 37 43 42 44 3f 3b 42 36 3a 31 32 4a 40 3f 3c 39 3b 3a 38 36 3d 38 3d 2c 35 35 39 30 3f 41 3e 30 37 35 38 33 38 40 2f 38 34 31 33 3c 37 3f 35 3d 37 40 35 36 41 38 36 3e 3e 38 37 33 3d 3b 3e 38 35 3a 32 30 36 37 31 34 3a 30 33 35 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 37 4a 48 47 39 3f 41 46 3b 45 38 40 47 3f 45 3d 43 3d 3b 49 47 4e 3e 45 49 40 48 4d 45 4f 42 4d 46 46 4b 4b 4c 38 44 3b 41 3f 42 3a 36 3a 2d 2b 1c 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 10 16 2b 3d
 46 43 48 3e 3d 3e 35 3d 34 33 3a 39 33 40 3d 3c 3a 39 3f 3e 36 3c 39 3b 34 3c 35 35 33 2d 39 35 3a 3a 3c 3a 37 3a 36 3e 44 42 42 3d 3e 42 30 3b 3b 3a 37 40 38 3a 3c 36 3a 38 30 3a 37 36 3b 40 3c 34 37 2d 33 35 33 34 2c 2d 23 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 39 4c 3f 45 40 3e 40 40 3c 42 49 44 4b 42 45 4a 43 49 48 44 49 4e 40 4d 4e 47 53 4c 50 50 55 58 56 52 50 49 4a 43 45 41 3d 40 32 30 33 22 21 20 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 20 2c 39 46 42 49 44 38 36 2f 39 33 33 2e 36 3f 3e 35 3b 3c 36 36 3c 2e 3b 3e 40 3e 3b 40 35 37 39 37 37 3f 3d 35 34 39 38 3d 3f 39 3c 3e 3e 3d 3d 39 35 34 35 3d 3d 3a 3d 36 32 3e 2b 3b 34 36 37 37 38 34 39 35 2e 30 39 28 2e 2a 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 29 45 44 39 39 3c 41 44 3b 38 3c 44 48 49 44 4d 4e 51 50 56 4c 4e 54 52 55 52 5e 67 60 62 63 66 62 64 59 5b 5d 59 4f 42 39 32 34 28 20 1b 12 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 1a 2d 3e 3f 4d 44 45 35 3d 35 3b 3a 3f 36 37 39 38 38 3a 42 30 36 39 29 3a 38 39 37 36 38 3b 3a 40 38 3d 36 39 39 3f 37 3b 41 38 41 46 38 3a 3f 36 39 32 31 38 35 3b 35 38 3a 39 3e 41 2e 3b 31 38 39 32 31 35 39 2e 35 31 38 2f 30 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 19 3e 3f 40 39 36 39 47 43 44 42 49 44 49 4f 4e 53 53 5f 5e 65 62 62 68 5c 67 6a 75 72 70 73 71 6b 6a 6d 70 67 65 50 47 42 2c 26 20 25 0d 06 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 14
 1c 2f 39 43 47 44 44 3f 38 3b 30 37 34 3d 3c 39 40 3d 38 3c 3f 34 35 39 36 38 41 3a 39 3a 36 35 39 38 39 40 38 39 37 35 40 3e 3d 3f 32 41 31 38 41 36 38 3f 40 36 35 3d 32 3b 36 32 31 31 3c 39 43 38 3a 35 30 32 32 30 33 30 2c 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 41 43 45 3e 47 49 4f 4a 4b 51 54 5a 59 67 60 68 65 64 60 66 6d 6e 75 72 72 81 79 75 80 71 77 72 67 6e 5f 5a 59 4f 3d 38 26 20 13 10 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 09 1c 2e 35 48 49 42 3f 3b 37 33 35 31 3f 38 34 3b 37 3d 3b 31 3a 36 39 35 3e 35 38 3d 44 3c 37 37 3d 39 34 35 35 3a 39 41 39 3c 39 37 3f 31 35 3b 37 35 3f 30 38 43 35 37 39 36 39 2f 3a 36 35 3a 33 31 39 33 30 36 36 31 2f 27 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 39 41 52 53 53 52 55 42 5b 5e 62 6e 69 73 72 70 7b 7d 75 7f 77 78 76 78 80 7c 7e 7b 76 71 67 66 68 65 5f 48 41 36 33 25 18 0f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 15 1a 23 34 3b 41 3e 45 33 36 3e 37 38 35 38 3e 38 3d 3e 39 33 3e 3c 3b 30 35 39 38 39 39 34 39 35 35 3e 37 35 36 38 3c 37 38 38 39 3e 33 3a 33 32 33 31 37 38 39 36 3b 30 39 3f 34 36 3a 32 30 30 36 35 30 3a 36 30 30 33 29 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 47 59 5b 63 55 5d 5e 6b 69 6d 76 76 7c 76 75 7f 80 79 7c 79 70 76 7c 75 75 7d 76 6a 6e 6b 69 5a 59 56 42 40 39 2b 1c 0e 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 07 0d 13 20 2d 36 36 3d 3d 41 41 34 3c 35 33 43 3a 3e 3e 39 3d 37 34 3f 3d 41 3a 38 36 3b 42 43 3f 43 39 3e 38 36 40 35 36 3e 36 3e 38 34 3a 40 3d 3c 3c 38 35 32 3c 2f 38 3d 3a 32 39 3b 3b 32 34 3c 33 32 33 37 3c 35 2f 2a 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 23 49 5f 75 6d 71 73 7b 7b 75 78 7a 7c 78 7f 7f 7f 79 79 74 80 77 70 6e 6d 78 6b 6d 6a 6a 61 56 4d 50 3c 39 2d 1a 0f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 11 21 2c 33 36 3c 36 3f 38 3a 37 3b 33 34 36 3b 34 34 44 36 3f 39 39 35 34 3f 3b 3c 40 38 36 3e 34 38 39 38 3b 35 40 39 3a 3b 41 43 3c 42 3e 35 3e 3c 40 34 37 38 36 40 37 3d 35 35 38 36 37 30 38 2d 3e 37 32 2a 2e 1f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 27 58 6b 75 73 78 7b 74 7a 7a 74 76 7d 6c 76 7a 78 7b 6d 76 78 74 73 75 69 71 67 66 61 58 51 48 46 34 1d 27 15 14 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 13 16 2c 2d 3c 38 36 34 38 41 39 35 31 37 3c 3d 3d 35 37 33 33 3b 3c 36 3a 38 3c 3b 3b 39 36 32 3b 3d 36 3d 3d 3d 42 3d 39 3b 40 38 36 34 30 33 3a 3d 3d 34 37 35 36 3d 38 41 39 32 31 35 33 2b 35 35 30 35 2d 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 29 64 7c 7b 74 78 74 6e 7b 77 7d 78 7a 77 73 76 73 6c 6f 70 73 74 6f 62 68 59 60 56 4a 50 3d 38 22 1e 13 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 09 09 16 19 25 2e 34 33 35 32 3b 38 3a 3a 3a 3b 3e 35 3a 39 35 3c 3a 37 3d 3a 40 3e 38 3f 43 37 3b 41 39 45 36 43 41 3a 3e 37 3f 45 41 3f 3a 3a 3b 3b 41 3b 37 3c 3e 39 46 39 3b 34 2f 3a 39 37 39 3b 37 3f 34 28 25 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 5f 72 84 7e 75 75 76 75 78 72 6e 75 73 7b 74 72 6e 6b 72 6b 69 6a 5e 5e 5a 57 4c 46 3f 33 24 15 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0c 1f 1f 26 2e 2d 3f 38 35 3b 32 35 34 3f 3c 37 35 3c 3c 3f 37 3d 3a 3b 45 41 38 41 41 3f 40 44 40 3f 42 38 3f 45 42 41 3f 3e 41 42 3a 43 3a 3b 43 48 39 3a 41 42 35 39 3e 3c 38 36 3a 3a 39 42 38 39 30 24 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 26 5b 6e 80 78 75 7b 72 75 69 6f 71 71 73 71 71 63 66 65 66 63 5c 60 59 50 4b 3b 38 2b 2a 18 11 07 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 0d 1d 20 2f 39 32 36 31 3c 37 39 33 2a 38 3a 3f 38 31 3e 38 3d 3c 41 41 3e 3b 45 41 3d 44 47 4c 48 4d 4b 41 46 45 4a 44 40 42 3e 42 47 44 39 41 47 49 3e 49 4b 3f 42 43 42 45 3f 44 40 46 46 43 41 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1b 59 78 79 77 65 6e 71 6d 6c 6a 6c 68 62 6a 66 65 61 60 61 60 55 51 49 43 33 34 24 1b 13 0a 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 09 0b 10 1b 25 28 2e 30 34 38 32 32 34 34 38 41 39 3a 37 30 3e 3e 43 49 43 46 48 4b 49 4a 55 45 4f 51 51 4e 4d 4c 50 58 54 5a 4f 56 54 52 59 4e 4e 56 50 52 56 51 55 51 56 52 4e 54 4f 56 5c 59 5a 58 40 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 59 73 78 74 6d 68 72 68 6c 66 65 68 68 68 61 59 5b 57 4d 54 4a 44 39 32 24 1f 12 0c 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 1a 21 21 30 29 2f 2e 32 36 39 39 34 3e 37 40 40 44 49 4a 4b 53 56 4b 58 59 55 56 60 63 64 60 6e 60 65 62 63 6b 68 61 6b 63 64 69 63 65 65 66 5f 61 6e 60 69 69 6c 66 6c 6f 68 62 69 64 4c 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 52 68 75 6a 68 6c 65 68 63 65 66 66 62 60 5b 5b 54 4a 42 3e 39 39 29 1b 0e 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 14 0e 13 20 25 2d 2d 36 34 2f 3d 3b 3c 3a 3e 44 42 51 51 5f 56 5d 65 5b 5c 65 62 68 6d 6d 72 71 6e 75 73 6f 72 6f 75 6f 73 6f 6f 6c 77 74 71 74 70 72 73 71 76 74 73 70 72 73 6e 73 67 56 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 4b 6a 6c 6b 6c 69 63 63 5d 60 5b 59 5b 51 4e 4a 40 42 35 2f 28 1d 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0c 0d 10 19 25 23 2a 29 30 35 3b 38 37 3d 4a 4e 57 52 58 5f 68 60 65 6b 6b 74 6c 73 70 6d 77 75 77 7b 72 7b 75 73 74 79 7e 78 70 7d 7f 85 77 79 77 76 7a 74 77 70 78 71 7e 76 6d 65 53 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 3e 62 6f 69 5f 60 5a 5a 57 5d 5a 59 4c 4f 40 39 3a 34 1d 1b 09 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 04 08 0e 13 19 20 2a 2a 39 30 38 34 3d 49 4d 56 5f 60 62 5c 65 68 6a 65 6c 6d 71 73 76 78 71 71 79 78 73 77 7c 73 7a 73 7a 76 76 80 7d 80 79 75 7a 78 73 74 75 75 7b 77 72 68 6b 4f 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 3d 59 61 61 5c 52 63 5a 49 4d 51 44 43 3f 34 33 29 19 10 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0f 10 1c 23 28 32 28 33 38 39 41 4c 51 54 55 5b 63 63 60 6a 68 62 63 6f 6c 70 74 75 72 6f 6b 71 74 7e 72 6e 79 6f 70 6e 77 7b 77 76 73 70 6e 74 72 6a 76 71 6c 6f 65 4e 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 36 56 5a 56 54 54 52 4d 44 3a 3a 38 31 2b 19 19 10 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 09 12 20 20 1e 24 28 35 40 41 45 48 4d 54 5e 63 5a 5b 63 63 66 6e 6a 6c 60 6a 72 70 75 79 6b 73 6b 6e 72 72 69 6a 6f 71 75 75 73 6f 6e 77 68 6b 76 67 68 61 5e 4e 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 37 52 5d 52 4d 42 42 37 3a 34 2b 21 20 10 06 05 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 0e 0e 14 1c 29 2d 31 32 34 45 45 4f 4c 58 59 59 65 5e 67 63 63 6e 6d 67 71 69 6a 6d 69 69 6c 6a 68 6f 70 74 72 70 71 64 6f 6a 6c 6a 6b 67 72 74 64 6b 66 4d 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2a 46 51 4d 3b 42 30 2f 26 1c 15 13 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0b 13 12 19 1e 27 28 32 37 35 31 4b 45 50 52 52 5a 5e 63 5f 65 5f 62 63 65 6d 65 69 6d 5f 66 60 5f 66 6a 66 5d 60 68 66 72 67 6a 61 6e 6f 60 65 62 48 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 49 45 32 2f 24 1f 23 1c 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 08 0f 0e 18 1b 26 2d 34 31 2f 35 41 47 53 4c 49 52 50 5e 5c 5c 5c 64 5e 64 67 65 59 60 64 69 6c 61 61 65 62 61 62 64 63 5d 64 67 5e 61 58 55 4b 19 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 17 2a 24 28 17 11 11 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 13 12 14 1c 22 26 28 31 33 3a 33 43 44 47 50 53 4f 53 53 59 57 5d 5f 5b 51 5e 5f 66 64 5c 60 5a 60 5e 61 5f 5f 63 65 66 5a 5c 58 5b 4a 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 1f 18 10 0d 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0b 13 13 0c 18 1b 25 2f 2e 2d 3b 39 38 3e 44 4a 50 4d 50 54 55 5c 56 57 56 5d 5a 55 62 59 57 5e 59 56 5b 51 5e 56 5c 55 61 5b 45 1a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0c 0d 0a 10 1a 1b 1c 25 2b 33 26 33 30 39 3b 3c 47 4e 4c 4c 53 51 4c 55 57 5c 53 5b 50 50 55 54 59 54 4e 57 4c 52 4e 44 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0a 0e 15 14 11 1b 16 1f 20 20 26 2f 3a 42 42 40 4a 41 4e 4c 44 4f 4b 52 49 4f 4a 4e 51 48 4d 48 46 42 45 43 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0c 0b 06 05 0f 0f 0d 1d 21 30 30 35 3c 3f 31 3e 3a 3e 42 3a 3d 3c 44 3f 39 41 33 39 37 35 38 2f 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 10 17 1e 1b 23 1e 23 28 1c 2a 2a 2a 27 23 24 28 22 20 25 20 20 19 1b 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 04 09 0e 08 12 0d 0f 0e 12 16 12 0c 0d 0b 09 0e 0d 0b 0e 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
