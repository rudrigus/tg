 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 04 02 06 05 03 02 0d 10 12 11 06 0c 13 10 0a 14 1a 1e 28 22 21 21 21 22 16 1c 1d 11 0b 0d 19 1a 34 2d 28 31 38 34 22 13 13 05 06 05 03 04 06 05 08 02 09 1b 15 15 13 06 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 0a 0d 03 09 06 05 03 06 07 05 08 07 08 0a 14 10 18 0c 14 19 12 10 1d 12 21 24 22 22 19 29 33 32 2c 32 32 3f 64 60 48 3b 22 24 24 37 35 40 50 43 3e 50 5a 51 32 23 11 12 0e 05 05 14 15 09 0d 12 18 1d 17 1b 21 1e 12 14 06 05 03 00 06 0e 0f 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 08 00 06 13 0e 0a 07 05 0c 09 0e 10 0b 16 19 1f 1e 18 14 14 0e 1b 27 26 2d 38 37 3a 43 3c 35 3d 50 5f 5d 49 4f 6e 76 73 58 4f 47 46 46 60 6a 65 76 6d 6a 6a 5b 49 3f 33 2b 26 13 17 19 2b 25 22 1e 1f 12 1a 17 1e 15 1f 17 0f 14 0a 08 01 07 1f 20 1b 07 05 03 02 06 05 03 02 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 07 03 05 06 05 10 0d 0a 13 07 0e 13 15 0f 11 1b 14 18 24 2d 45 3d 30 2b 33 30 41 5f 52 5b 63 6e 69 5f 5b 57 61 6d 73 71 72 7f 84 6b 64 5c 56 66 65 65 65 6f 78 82 95 a8 86 6e 67 68 62 5f 5e 57 53 4e 50 52 49 3b 34 2e 2e 25 1a 1d 1c 20 27 1c 14 12 12 0f 1c 16 21 1d 0d 11 09 06 0b 07 09 0b 05 03 00 06 05 03 04 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 08 06 05 0e 0a 06 09 0e 05 0a 06 09 0c 14 0f 09 12 15 18 21 25 21 26 3c 43 3e 5f 7b 6b 63 65 6b 65 6a 71 7c 69 67 78 73 65 5d 57 65 6d 69 79 72 79 6a 66 65 69 6a 6f 71 62 6f 79 78 8e 8c 80 7c 6f 76 70 72 73 75 6d 77 75 79 6b 64 62 59 4e 4c 40 37 38 34 3b 35 3b 24 1e 1a 1e 1d 1d 16 15 13 11 0f 15 05 0b 06 05 03 03 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 07 00 06 0e 0e 06 15 11 13 0e 09 0e 1e 12 1f 1b 22 2a 29 2c 39 3f 45 45 50 53 50 74 8f 98 a2 94 89 7b 6f 5c 6d 5d 5e 65 5f 60 64 65 64 6f 6e 67 6a 72 72 6a 6f 6d 6e 73 74 75 71 79 75 7f 82 7e 76 77 75 75 6e 84 76 75 78 7a 79 70 6d 6c 6b 6a 65 52 55 54 52 4c 4b 49 3b 48 3d 35 2a 34 25 25 1a 18 06 10 0d 0a 0b 07 0a 0a 0d 05 08 01 08 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 0a 11 0d 0f 19 13 0f 17 18 1f 1b 1c 23 24 41 42 45 46 4b 41 46 57 61 5e 70 69 80 86 9a a9 a8 a0 8e 81 79 68 66 69 64 64 5e 6b 67 6d 6b 70 6e 76 71 73 71 72 72 78 77 77 7b 80 7b 7a 7b 7f 7e 83 7d 80 74 80 7b 7e 7e 82 7a 7b 75 77 77 6c 74 69 60 58 53 56 4e 52 55 53 4b 4e 4a 49 49 46 46 36 3a 39 3e 2e 18 0e 19 13 0c 10 13 0e 09 08 0d 0a 0a 10 12 09 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 03 06 05 04 00 06 05 03 01 0d 08 0b 08 06 16 15 12 10 1b 20 1c 24 2a 29 2f 34 31 40 52 5f 65 6f 74 73 6e 74 84 86 92 8f 90 87 90 a1 91 96 8f 89 8b 86 7c 77 79 6f 73 70 73 6c 77 75 77 78 76 75 75 78 77 79 81 7a 7d 7c 78 7c 82 86 7c 88 78 7c 85 7c 88 83 7c 84 7f 7c 7b 74 73 6d 6f 6e 68 68 5d 5a 59 54 4f 4b 4c 49 50 51 51 4d 51 4d 48 4c 5a 54 4d 48 3b 3d 34 2a 25 2a 25 19 11 13 0a 0d 08 06 0d 14 05 07 05 03 02 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 07 06 05 0d 0b 07 08 0f 12 1c 1e 16 25 2a 29 2b 37 3c 3e 51 56 51 55 54 58 67 6e 80 80 85 96 84 8e 8b 8b 7b 7e 79 74 73 72 80 84 84 84 87 81 85 80 7c 7b 76 72 71 7c 74 78 77 76 6e 71 7c 7b 73 7b 77 73 78 82 7d 7b 84 84 7e 84 7c 7e 82 83 7b 84 7a 82 78 7f 78 69 72 6c 69 64 62 60 5f 59 56 53 5b 53 5d 51 4a 55 4c 4e 4d 4f 52 5c 5e 5b 57 57 4d 46 42 3c 4a 3d 32 27 18 1b 17 0b 16 0b 03 01 06 05 05 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 08 06 05 03 00 06 05 03 02 06 05 03 0e 06 05 09 12 0d 0d 19 11 1b 18 24 2a 29 2f 36 44 42 54 5c 62 68 76 73 7a 70 64 62 61 60 64 68 72 6f 75 7c 79 7a 7f 7a 73 74 75 7c 7d 7b 83 88 7f 85 86 88 86 74 7c 79 7a 7d 7b 7f 7f 7a 80 79 7c 84 79 7a 79 78 81 78 83 80 7e 88 80 85 84 86 85 85 82 7c 85 84 80 7a 78 7a 6d 70 6d 69 6b 67 5f 64 60 59 5f 56 5d 59 56 5b 53 53 59 5a 51 4a 5b 55 59 59 5f 61 4f 55 5a 5e 66 57 41 29 2f 21 2a 22 1a 11 0b 18 0d 03 05 06 05 05 01 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 07 05 03 0c 10 10 0a 0a 14 14 15 17 1e 1d 1d 27 20 31 33 3b 44 4a 58 62 6d 76 85 8b 89 7d 76 76 5f 68 69 66 62 71 70 6e 71 6d 73 73 70 79 7a 7e 77 78 85 7d 7e 79 7b 81 82 85 81 85 7d 82 85 81 7c 84 7f 8a 87 84 81 8b 85 79 7d 7e 7b 7d 82 7e 7d 84 8d 8d 8c 89 90 86 80 8a 87 86 85 7f 71 79 7e 75 70 72 69 71 6e 70 6c 6b 6b 65 66 62 67 62 60 5e 56 5a 5f 56 51 57 54 5e 58 58 57 57 56 60 6b 75 71 4a 4b 35 37 32 2c 17 1e 1f 20 24 21 14 17 15 09 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0d 13 15 18 1d 1f 2e 33 39 46 4b 4d 46 4d 4b 57 6f 7a 83 7e 8a 86 7f 7c 6e 6e 6f 66 67 6a 6a 6c 6c 66 73 6f 6f 65 77 7b 70 78 7e 7e 7a 80 80 84 85 85 86 8f 91 8b 8d 8a 88 8a 87 85 80 83 81 8a 88 8e 87 89 7d 8a 82 86 88 83 87 82 85 88 8c 85 8a 90 8a 83 90 88 8a 90 85 8a 7d 7e 7d 78 6d 6d 71 77 74 78 79 73 74 72 72 75 6e 6e 6d 68 68 62 54 5c 5a 5f 5b 55 5a 4f 53 55 5f 61 5f 68 71 70 60 5b 50 4a 4b 41 2e 2c 25 28 25 1f 1e 1c 14 0b 06 0c 03 03 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 06 09 0c 0a 10 16 11 1e 24 2a 39 37 3c 3d 4c 60 6e 7a 7e 7b 80 84 91 89 7f 7b 72 74 71 6d 6e 70 6b 63 6b 69 69 6e 6e 79 6b 71 74 6d 78 7c 7b 7d 80 88 89 86 8d 85 92 89 92 93 94 95 96 a3 9d 96 9c 92 99 91 9c 98 95 90 95 90 8c 89 84 87 87 8c 85 8b 8d 8c 8a 92 8b 93 8f 8a 85 93 8b 90 89 8d 7a 84 82 7f 80 79 81 7d 84 77 85 82 80 83 85 86 75 7d 79 6e 70 6e 61 68 5d 67 5f 5b 5d 61 65 5e 5d 5e 60 60 6a 69 6d 6d 5f 5e 5e 5d 59 4f 3b 35 2c 30 23 1d 1d 1a 12 13 11 04 0c 05 06 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 01 0b 05 0f 10 13 12 19 2a 25 35 3d 44 4a 4d 50 4e 59 62 6c 7b 85 84 85 7d 7b 71 6d 76 6f 6d 70 70 76 70 6a 71 6e 77 6e 76 73 6b 74 6d 76 75 7f 7f 85 87 8f 95 8f 99 9d 9a 9d 97 9a 9c b0 af bc b6 b8 bd b8 b3 b3 a7 b3 a2 a6 a8 99 98 8e 92 91 98 8f 89 8f 97 85 93 8e 95 9c 8e 8f 90 91 8c 91 8f 85 8c 83 89 91 81 87 88 8a 8b 8c 8c 90 8e 93 9d 94 90 85 80 85 7c 7c 76 66 70 63 64 64 65 5b 61 67 5b 63 60 5d 60 67 5f 58 5b 5e 60 62 61 5e 5d 65 55 44 47 30 29 29 1a 18 11 14 16 0c 11 08 01 06 0a 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0c 08 0d 0d 13 13 1d 1e 2a 33 3b 3b 44 4c 4c 55 54 60 62 55 5c 5c 63 72 72 72 71 6c 6d 6d 6c 69 68 70 70 76 72 6a 6c 6e 6a 6d 6f 75 75 6e 76 75 7b 87 89 89 8c a2 99 9b 9d a0 a6 b3 b6 bc c3 ce d8 db db dc e3 dc d4 db da c9 c6 b6 b9 b1 af ad b0 a3 a0 99 96 9a 95 9e 92 9b 9f 99 a1 8e 93 90 8d 94 95 93 93 94 96 90 92 93 95 91 99 93 9d a6 9d 9e a0 9c 9b 96 89 8a 90 7d 7b 75 6c 69 64 68 6c 62 68 64 62 62 64 5d 63 5e 56 55 63 52 5a 55 52 57 5a 65 6a 64 60 5b 42 32 25 11 14 14 13 12 15 12 08 0b 0d 07 0f 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 06 06 05 03 07 06 06 12 10 16 1f 23 2d 35 40 4e 50 56 54 58 5c 69 5d 5f 5e 5b 5e 62 69 68 6a 73 6f 75 77 77 6d 72 74 72 6d 74 6d 76 72 68 75 77 7a 81 78 7e 88 8d 88 92 89 8a 9c 9a 9b a8 b3 b4 b4 c5 cc e4 e9 fd ff ff ff ff ff ff ff ff ff f5 e9 df dc d4 c9 c2 c2 c0 b9 aa b5 b0 ad a9 a5 a6 a8 a3 a7 91 9c 99 99 a2 9f 96 99 9c a0 9e 97 a8 a4 a5 aa a9 a4 ab b2 ab a9 9e a0 9a 9d 8d 8a 86 7e 7e 6b 79 72 64 6c 69 6c 6e 65 68 5f 59 60 62 55 5b 57 60 5a 5a 54 5a 5f 63 64 6b 73 72 61 5f 42 2b 26 1d 12 1d 1b 12 18 15 15 07 06 07 0d 0a 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 07 0b 0b 14 18 15 22 22 30 31 41 50 4e 55 60 5a 61 5f 5f 68 64 66 5b 62 65 67 74 63 6c 67 6f 6c 82 6f 7c 75 7f 76 70 77 6f 77 73 7d 80 7b 7d 81 7f 90 83 94 8c 92 a0 9d a4 b0 af b6 b9 c6 d2 df f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 f5 e5 e3 d7 d9 d1 cc d0 c9 c3 be b5 a7 a9 a6 9e a4 9f a2 a1 a1 9e b0 a7 ab ab af ad ae b5 b0 b9 b6 b9 b2 bb ad ab a9 a5 99 9c 8f 86 86 79 78 75 74 6c 71 64 66 60 6d 66 61 65 5e 62 5f 60 55 59 62 60 59 55 5c 5a 59 60 5c 59 72 70 64 56 44 2d 2f 26 1c 19 1f 13 0b 11 15 10 15 10 0d 0f 11 0a 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 08 12 15 0f 1e 1b 24 36 33 42 46 51 5d 57 5b 5f 67 63 5d 5d 70 6a 62 6d 6a 68 66 65 69 71 70 70 74 75 6c 74 78 7d 7b 79 73 73 7b 79 7e 81 7a 87 86 8a 88 97 8a 97 9b 96 a8 a3 b7 b6 c3 ce d5 e1 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff ff f4 f5 ed ee de d5 b8 b0 ad a8 a9 a5 a6 a5 a6 a7 a8 b4 b4 b4 b1 b8 b4 b8 bc bb bd c8 c4 c5 be b8 ab ab a4 9f 9e 96 8a 86 80 7c 79 6c 71 71 71 6b 6d 68 5a 63 5a 5d 64 60 5d 60 59 54 58 60 60 56 55 54 55 59 55 65 6b 74 75 67 60 4d 38 2d 1e 20 1b 19 1b 1c 14 16 0e 17 0c 0d 06 01 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 03 05 06 08
 08 0d 0c 13 19 20 27 31 39 45 4c 5b 58 62 63 68 65 5e 64 61 6a 6a 69 60 61 65 6b 71 69 6c 70 6c 73 77 7d 72 6e 74 7b 7c 7e 7e 7c 7b 7b 7c 7e 84 86 85 8f 97 96 9d 9d a3 a9 a6 b1 b2 b5 bf d1 e2 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe e7 d0 ba b6 ae b2 a6 b1 ae b1 b0 b8 b4 b7 bc b8 c3 b9 c8 bf ce ce c6 cc c6 c9 c6 bd b2 aa ac a5 9a 92 8c 7c 7a 78 78 6e 78 73 6c 77 62 6b 64 68 64 6c 5b 60 60 61 5f 5d 58 5d 59 5b 59 54 55 56 5b 5f 62 6d 75 6b 5f 5f 52 3f 32 23 17 13 17 17 15 16 16 12 14 03 09 0c 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 03 0f 0b 14 1c 1e 1a 24 1f 32 39 4b 57 5f 5e 5f 61 66 68 69 68 6b 6a 6a 6b 6b 6d 6b 6d 6e 74 6b 6b 6f 78 73 75 75 79 78 78 7d 78 73 83 7c 84 84 7d 82 86 88 8d 93 99 a4 9a a3 a6 a9 b4 ab ad b9 bc cc e8 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb cd be b6 ba bb b9 ba ba c1 b7 c2 ba bd ba c3 cd ca ce d1 cd d2 cf d5 d3 ce c3 bf ba ab a7 a6 96 90 84 7e 80 7f 7e 78 80 70 79 70 6a 6b 67 68 61 69 66 6a 5e 5b 64 64 5c 62 60 5e 5b 60 52 5b 65 61 6b 6d 6c 66 5f 55 52 44 48 33 20 22 20 13 19 13 11 19 11 10 0c 09 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 07 0d 0b 18 16 21 1f 26 29 40 4e 64 6f 72 69 67 5e 60 60 6a 64 69 5e 62 66 64 67 6a 6d 6f 70 70 76 77 72 76 76 71 74 7c 7e 83 7a 7a 7b 7a 84 84 7f 7e 84 8b 8f 95 9c 9e 9a ac a6 a5 b0 af b1 bc c0 c9 dc ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dc c2 bf bc bf c2 bc b9 c2 bb be c5 be c6 c8 d0 d7 d4 d7 d9 dc dc d1 d6 cb c8 c3 b7 b5 a5 a7 96 92 8b 8d 8a 7e 86 84 85 82 7f 72 70 69 70 6b 68 63 60 6c 64 64 69 64 60 64 60 61 5c 5c 5d 56 5c 59 58 5c 5f 5d 53 50 4f 51 46 3f 43 39 28 26 13 16 0c 13 12 09 0d 12 09 0d 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 06 14 15 1e 21 22
 22 2d 3a 44 55 72 7a 77 66 65 65 65 65 62 60 65 69 60 69 6c 6b 6f 70 72 74 77 6f 79 75 73 75 84 85 85 85 8c 7f 80 7a 84 86 85 85 89 81 8b 88 8d 97 95 a4 a4 aa ae b3 b1 b3 c1 c6 c7 d8 e8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb cc c5 c0 c8 c4 c5 bc c4 c2 c5 c0 c9 cc cd da dc db d5 db da e3 e0 db d5 d1 cd c5 bc ad a9 a2 9a 96 8e 8f 8d 86 87 7e 83 7c 76 79 70 6e 6f 6f 71 69 6d 69 65 68 6b 61 5c 5d 60 52 5f 5f 58 5b 5f 5b 5d 52 57 49 4d 47 4c 4a 4b 4e 4f 49 41 38 26 1c 17 16 16 10 12 0d 07 09 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 0e 0e 14 1a 1d 1b 21 28 31 41 55 68 65 69 6d 71 66 69 61 5c 61 60 66 73 6a 66 69 65 67 73 74 77 81 84 83 81 84 87 84 8b 8b 8b 91 90 83 86 84 8e 8b 86 94 8a 92 90 9b 8e 9f a3 ab b2 aa b0 ab be b8 c1 d4 d9 e7 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe de d0 cc d6 cc c9 ca c9 c1 c7 c6 d1 d3 d8 cf df e4 e4 e1 e2 ed e7 dd e1 d5 ca c9 c3 c2 b2 aa ab 9b 9b 9e 90 94 8d 8e 8d 84 79 70 78 72 75 76 78 6b 6b 70 77 72 6e 6a 6c 68 63 5e 62 5b 5e 5c 57 58 49 55 51 4d 52 53 4c 48 4b 48 60 6a 6b 54 46 29 16 16 18 23 14 1a 14 14 07 0d 0a 06 0a 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 05 03 06 06 0c 0a 13 17 24 20 25 3d 41 58 59 55 69 60 5f 66 64 61 65 5f 5a 63 61 6e 70 69 6e 69 70 66 74 76 79 7e 80 7f 89 86 8d 95 8e 97 96 99 96 92 8f 8d 90 84 8a 8b 8e 93 94 97 a2 9f a6 b0 b4 b2 c0 ba c0 cb ca d6 de f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e3 d5 d0 ce d4 d1 d0 c6 c5 cf cc d6 d4 d8 dc e1 e5 ec e8 ec eb e4 e3 e7 e3 d6 cb c9 c4 be b7 b0 a1 9d 9c a4 a3 9a 9c 85 8d 86 7d 74 82 71 7c 75 7a 7b 75 7b 6d 71 6a 6f 6d 6b 71 60 63 63 5f 5e 5b 5c 50 57 55 4d 58 58 55 4d 4f 5c 75 79 64 58 35 34 20 19 1e 1e 25 18 15 09 08 09 11 07 09 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0f 05 04 0a 08 14 19 1d 1d 29 38 49 52 70
 6f 61 60 5e 5a 5e 64 5e 59 63 5f 65 65 67 6a 67 65 69 68 73 73 74 72 7c 7c 84 88 8a 94 96 8f 9b 9e 9c 97 9e 9e 95 9b 97 9b 98 92 94 8d 9b 9e a0 a7 a4 b0 b3 b5 c2 c7 c7 cf d4 da e8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e1 d3 d9 d5 df ce d7 d0 d1 ce d6 db d2 e0 e4 e4 e4 ee e8 e9 f1 ea e6 d9 d0 d5 d0 ca c4 b8 b5 ad a4 aa a6 a5 9b 92 93 91 89 86 8a 88 82 86 82 71 7d 76 73 7b 74 72 70 65 69 66 67 6d 63 59 5d 57 5f 58 55 4d 4b 55 59 57 51 56 5c 5d 6e 57 4f 4c 44 2f 20 24 25 1c 1d 1e 11 0e 06 09 06 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 05 0a 09 0e 0f 1a 1a 25 2b 30 45 5f 5a 69 6d 65 62 63 5d 68 66 5e 68 63 69 68 62 6a 70 68 6b 72 6f 73 78 6d 76 80 81 85 89 8a 96 9c 99 a1 a3 a6 a0 a5 ac a6 9f 94 a0 a1 a4 a4 a3 9f a0 a4 a6 a6 b1 b6 bc c1 c9 ca c9 d4 dc e2 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ea de e4 e6 e0 d7 df d8 d5 da dc e9 de e5 e5 eb eb ed f5 f0 eb e9 eb e9 e2 e0 da cb c7 c6 c4 b3 ba b5 ad af a9 9c 9e 92 8f 8e 8e 8a 8b 70 84 7d 80 7c 7a 79 77 77 77 6a 68 72 75 6b 67 6b 5b 63 5c 5c 60 61 54 58 5b 57 57 4c 52 5a 62 5e 5c 5d 55 45 35 37 2f 2b 29 25 1b 1a 10 0f 11 0d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 0d 10 16 1b 29 39 3c 41 50 6f 6c 66 6a 64 67 67 63 66 65 69 68 68 6b 68 71 69 70 68 6c 6e 70 71 74 81 75 7b 81 7d 97 8b 96 94 9a a7 a2 ab aa b2 ad b7 b5 ad b2 b4 ae a3 a7 a8 b0 b0 a8 b3 b6 b9 b7 c6 bd cf d9 d6 e3 df ed fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f0 f2 e8 ef e7 e3 eb e3 e7 e6 e7 e9 ea f2 f0 f2 ee eb ee f0 e9 eb e2 df d8 d6 d1 cc c1 ba b8 b9 b9 b1 aa a3 a2 9c 92 8f 9b 8a 89 92 81 88 82 7c 75 7d 76 7c 7f 77 78 76 6e 6d 74 67 62 66 60 62 5c 5f 57 58 5b 57 55 58 5a 5a 5d 62 60 69 5a 58 4b 3a 46 3b 28 1f 24 1b 17 12 0a 16 04 06 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 0d 0a 0d 1e 2a 31 44 45 54 68 79 8b 87 6f 67 64
 6b 68 69 71 6f 6d 70 70 76 7a 6e 7d 6a 73 75 75 73 6e 7c 7f 80 7d 8b 8d 8e 8d 99 a0 a8 a6 ac ad b3 b1 b7 ba b2 b6 b0 ba b9 b8 bd b7 b4 b7 b3 bb bb bc c7 ce c7 cf dd e5 e4 e9 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fd f0 f4 ec f5 e9 f5 f4 ec ed f0 f3 f2 ed f1 f3 f7 f4 f0 ef e6 df df db df d5 d1 cb c2 be ba b9 ad a4 a2 9e 9e 95 96 98 8b 92 8b 87 8a 81 80 76 7d 77 78 75 76 71 71 73 79 6e 6d 66 5d 5b 66 5d 5e 5b 5f 5f 5c 50 5c 5c 66 6a 68 65 5d 57 57 52 54 4c 3d 39 2a 29 14 15 1a 0d 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 07 06 07 12 12 11 1e 39 50 66 77 83 8d 98 a4 8d 70 6b 67 64 71 73 6b 70 76 74 7a 78 80 7a 7c 77 77 7c 7b 82 7e 7b 8d 84 89 89 91 96 95 9a a5 ac b9 b5 ae bb b9 be c3 ba bc c4 bf ca c3 c7 c7 ca c3 c3 cd d0 d2 ce d9 d8 dc e4 ee f6 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f8 fb f6 fb f8 fb f9 f8 f8 f7 f1 f5 f6 f5 f3 f2 f0 ed e8 e4 dc de d8 d5 cb c9 c1 bb bb b1 b0 af a9 a1 9d 95 98 96 8e 88 8b 8a 86 80 7f 79 81 80 7a 78 7d 7c 7c 71 7a 73 6c 76 6a 67 6d 65 66 66 64 65 68 5f 67 63 5e 56 5d 58 4e 5c 61 69 5d 55 45 3a 28 1f 17 1b 13 0d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0f 0b 0c 0d 0e 15 2b 2b 48 64 6d 88 93 9a a5 9c 82 65 67 6d 70 75 76 7b 7b 7f 79 8b 80 8a 88 87 89 85 8a 81 85 82 89 85 8e 95 97 8e a3 9d a3 b2 b2 b1 ba c3 bd bb c4 c2 cb ce ce ca c4 ce cf d0 d4 d4 cd d7 db dd df e2 df df f4 f2 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb ff fa fc fb f4 f4 f8 f8 f0 ed ed e9 ec db e4 db db d9 d1 cc ca c1 b9 b1 ae ac 9d a0 a0 9a 97 93 95 8d 94 83 83 7d 81 7a 7f 82 7e 79 76 79 84 78 6f 6f 6c 6f 63 6f 6f 6a 6a 6e 65 66 62 59 5a 5c 5c 55 54 54 5a 64 79 6e 5f 44 3e 33 25 1e 20 15 0a 0e 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 09 0b 05 10 07 11 20 2c 3b 50 60 6b 6c 80 86 89 84 83 76 6e 6e 6d
 75 72 78 76 79 7f 8c 8a 85 90 91 8d 94 94 90 94 8a 96 8b 92 9a 8f 9a 9a a0 a3 a7 ab b5 b5 bb c2 c3 c4 c3 cc c4 cb d2 d0 d6 de dd d8 e1 de de e6 e9 e6 f0 f2 ef f2 fd fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff fb fb f5 f8 ed ee f3 ee f2 f0 ed ee e9 e6 e3 d9 d8 d4 ca cd bc c0 bc b3 b6 a4 9e 9f a0 a1 9a 89 96 8b 87 85 8b 81 84 80 7a 80 79 82 7a 81 79 75 6e 6f 6e 6c 6a 73 71 6b 69 64 58 5c 55 5f 59 58 61 59 52 5a 60 6b 67 60 5a 45 38 38 2b 24 15 17 14 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 09 0e 07 05 0e 0d 0d 19 22 3b 4e 52 5b 69 6d 75 78 72 75 73 63 72 6d 70 6f 6f 7c 84 86 85 8b 91 93 9b a0 98 a4 92 9a 98 a6 a0 a4 99 a1 9f a8 a7 ae b0 aa bc b7 bb c1 c8 cd c9 cd d1 d2 d6 db d5 dd e0 ec e6 e2 e7 e8 f4 f9 f0 f7 f9 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fe ff ff f5 fb f5 f7 fa eb f0 ee ee f0 e8 ec e2 d3 d9 d8 cf cc c3 c1 bd ba b2 a5 a2 a7 95 9f 99 90 92 84 8a 8b 89 85 7d 83 84 84 8e 82 7d 80 72 77 81 77 78 72 71 72 66 59 5b 54 5d 57 5d 5a 56 5a 5e 52 5c 53 5e 5d 5d 63 5a 4a 3a 37 27 26 1a 1b 18 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 06 05 11 0a 0f 09 0f 0e 1d 28 39 55 62 59 62 65 6b 6c 75 6f 71 6f 73 6e 6f 6f 79 80 7b 82 88 8f 9e 98 9e a3 a6 a3 a6 af a9 af a7 a5 a1 a5 b0 ad b2 b5 b1 b7 ba be ba c3 c5 cd d4 cc d2 d8 d6 de d7 df e9 e9 f0 ed f5 f9 fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa f8 fa f7 f2 f3 f8 f4 f6 ed ef e1 e5 e2 dc da d3 d1 c6 c1 c5 bf b3 ab a0 a4 a7 a6 99 97 93 8e 8e 88 91 85 84 84 8b 86 80 85 84 7a 7d 80 7c 70 70 6f 5f 64 66 60 5e 5b 5b 5f 61 57 5f 56 59 52 52 53 50 5d 54 59 5b 60 51 44 3c 34 23 27 1d 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0e 0f 0b 0a 11 14 1d 1e 34 4a 5f 69 64 61 61 71 70 71 73 71 74 70 70 76 7b
 7f 7d 83 88 8b 8e 95 97 9d a6 a4 ae ae a4 b6 b0 a9 ad b3 ad b2 b2 b9 bf be b6 c4 be c9 c6 c7 c6 d5 d4 da d5 da e7 de eb e8 ef fa fc f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 fb f6 f6 f9 ef ee f5 f4 f0 f1 ea e5 e7 e4 e2 d9 d3 d6 cb bf bf be b7 b1 ae a0 a5 a0 97 94 97 92 8c 93 8b 87 8e 84 82 7e 80 78 83 7d 79 76 73 67 68 6d 65 6a 66 65 5d 5f 5f 55 5c 58 55 5a 56 55 59 50 53 58 51 5c 63 6b 63 50 43 3f 33 26 16 11 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 05 06 10 0d 0e 15 0d 0d 14 16 28 2a 4e 5d 67 5a 65 6a 5f 62 6b 6a 6f 6e 7b 7d 76 7f 81 80 80 83 82 8c 93 9b 9e a0 a8 a4 b1 b1 af af b1 b7 b7 b3 bc b5 be c0 bb c1 c2 c2 c8 c9 ce d3 d1 d3 d6 da e1 e6 e1 e5 e8 f9 f4 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 fb f5 f4 f9 f6 f4 ef f1 ed ec e5 e2 e4 e6 d9 d6 d1 c6 bd bc b9 b6 a9 a1 a4 a3 96 96 97 94 89 90 87 8a 85 81 7e 7c 7a 7c 7c 78 72 75 6f 68 67 66 69 65 66 65 5e 5d 58 50 65 5c 5f 52 53 52 5f 59 59 54 5a 52 54 72 74 62 59 4a 30 22 16 0d 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 09 10 11 0c 16 14 19 13 12 1f 23 2e 44 63 6e 67 5a 61 61 61 69 73 6d 78 7e 7e 7d 85 81 87 8f 8b 89 8e 95 94 9d a5 a4 ad ae ae b7 b3 ba c1 bc bc c0 c4 c1 c0 c6 c1 c4 c4 cd cf d6 d0 d6 d7 d9 da e2 e4 e5 ea ea f4 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f6 fb fd ff f8 f8 f6 f0 f3 f1 f3 f2 f0 e7 e2 ea dc d5 d1 d0 cb c6 b0 b5 ab a8 a6 a3 a0 9b 95 8b 8c 8b 84 83 89 88 83 7f 78 7a 76 7b 74 76 71 68 6f 67 6e 68 66 6a 66 5d 66 5c 64 55 5d 5e 58 54 5a 59 57 58 53 5b 67 79 7a 6c 56 52 3b 2f 22 12 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 08 0b 13 13 1b 17 0e 14 21 2b 3c 50 5d 60 59 60 58 62 60 62 68 6e 6f 79 74 7e 83 8a 86
 92 89 90 95 93 93 a1 a5 aa af b1 b4 b1 c4 be c9 c4 bf c6 c6 c7 cd cd c9 d3 cb cd cd d4 cd da d9 da d9 e0 e4 e9 ef f0 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff f9 f6 f6 f3 f4 f5 ef f1 ef e6 e6 dd de da d6 d1 c9 c2 bb b4 ae ad a6 a1 9d 9b 99 8d 90 8b 84 88 7d 82 7e 85 7a 7b 79 7d 78 78 73 6f 75 73 6d 69 65 69 69 59 64 5c 63 58 5c 5f 64 55 5f 59 57 5a 5d 5c 64 7a 83 7e 6e 51 37 35 23 24 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 0a 0d 1c 17 20 1c 19 20 23 45 4b 53 5a 5e 5f 5a 61 5b 5f 5e 69 64 6d 74 76 7e 88 8c 8f 92 95 9b 96 99 97 9e a2 b0 b5 b0 b7 b4 b3 c1 c2 c9 ca cd d1 d2 d0 d1 d0 d4 d0 d6 d5 da e0 dd db db de dd e7 ec f5 fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f9 f3 ff fb f5 ff ff f9 f8 f9 f6 ef f2 ee eb f0 e2 e2 d8 d6 d1 d0 cc be c2 b1 b1 a8 a9 ad 98 98 99 8c 90 90 8a 83 80 82 83 82 81 7d 84 79 7c 81 7a 71 76 69 6c 6f 6b 6c 64 62 5f 57 55 61 61 58 63 5d 63 59 5d 5e 54 50 5f 77 83 7b 6a 56 43 35 28 1e 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 11 11 10 1f 25 20 25 33 32 2f 3f 4f 5a 5d 58 5e 61 60 5e 5e 6a 6a 73 70 6d 6a 75 78 7a 8b 97 95 98 9c 98 9c a5 a7 aa ad b5 b0 b7 c0 c6 c2 cf c9 cb d0 d1 d6 d8 d8 d8 d6 db dd e4 dc dd e5 e4 ed e5 f0 f4 f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff f9 fe fc f7 ff ff f3 fd fa fd f7 f5 ee ee e9 e2 e1 e4 d5 ce d1 c7 c4 c4 bb b0 ac aa a0 a4 97 90 95 98 91 82 84 83 8a 83 78 7e 7d 87 77 79 7b 7d 76 76 78 74 73 6e 66 65 62 65 68 62 65 66 64 64 60 60 61 5c 59 52 5d 57 74 82 75 60 5b 43 3e 2f 23 1c 07 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0e 0d 15 14 1d 23 31 3b 45 50 4a 58 65 66 5c 5f 4f 5d 6d 6a 5d 6a 65 62 74 65 6e 81 7a 81 86 86
 97 9b 9c 97 a3 a3 a8 af b4 b6 b8 c0 c7 c9 cb d2 d2 d0 dd e5 d4 e0 de df e5 e3 e5 ec e9 ed f1 ef f7 f7 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff fb fa ff fa fe ff f6 f7 fa f8 f6 f4 ec ef e9 e9 e1 da de d7 cb cd c7 c2 b6 b6 b1 b2 b1 9c a6 9e 9a 9a 9a 93 8b 84 84 88 87 85 80 8e 85 80 81 80 77 7a 80 79 74 71 6d 69 75 6b 6e 69 64 65 66 6b 65 6b 5e 58 5f 5e 5d 5e 63 75 7e 73 69 58 45 3e 26 16 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 10 0c 1a 1b 22 30 3d 54 5a 69 6d 7b 87 6e 59 59 5f 63 60 5a 62 61 69 6e 6c 7d 79 79 7d 88 86 8c 90 9e 9d 9f a9 9c a7 ae b2 b1 c1 c1 cb cf cb d3 dc d9 d8 e5 e9 df e9 e9 ea ed f0 ee f7 fb fa f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fa ff ff fa ff fe f6 f5 f9 f9 ef f6 ed ed e9 f4 ec eb e0 e3 e0 d6 d3 d0 cb c3 c4 c0 bd b1 b4 ad a7 a5 a2 98 9e 96 8e 90 88 8a 8d 8c 8a 88 81 88 84 7e 81 7d 7b 78 79 7c 7b 73 70 76 7a 78 6e 6a 70 6f 66 6a 71 60 60 61 60 56 5b 54 60 75 74 73 60 4b 3e 31 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 06 12 12 16 1a 27 3a 3e 4d 56 70 7b 8e 8f 90 74 65 51 5d 5c 64 5f 66 65 6f 76 7d 7b 80 8d 84 86 8d 83 94 a0 9f 9b 9d a9 aa b4 bd b2 bd be cc d3 d7 d4 d9 e0 e6 e4 e8 ed f0 f1 f0 ef f4 fb f4 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb ff ff ff ff ff fc ff fd f6 f3 f9 f5 f9 f1 f4 fa f2 f7 f0 f4 ed e9 e3 e9 eb e2 e2 da da d9 ce c9 c4 c6 be bd b7 b1 b8 b2 ab a3 9d 9d a1 9f 99 8c 8c 89 92 8c 90 8f 86 87 8a 89 86 85 82 82 7b 81 7d 7b 79 7a 73 7c 76 7e 73 7b 68 6e 6d 69 68 60 5e 5e 5b 5e 64 7b 78 63 4e 38 21 20 16 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0a 12 0e 1c 1f 26 35 3f 46 5b 65 7d 8f 96 95 7b 6d 56 59 50 5f 60 64 5f 63 6b 6c 77 80 85 93 8f 89 93 98
 94 9a 9b 9d a4 a4 ad aa b6 bb bb c7 c9 db cd db e5 e7 f0 f1 f5 f8 f3 f9 ff fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ff fa f6 f9 fd fa fa f4 f1 fa f3 f8 f6 ef f1 f1 e8 e6 ef ed df e1 da dd da d9 d2 d1 cb cd c2 c3 c6 b8 bc b7 af ab a5 aa a1 9e a5 9d 96 98 99 97 95 94 94 91 92 89 8a 87 87 87 88 83 83 83 7e 83 7f 83 80 7e 75 7c 76 7a 6f 71 62 6b 60 60 57 56 5a 69 75 75 5e 4a 27 1f 15 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 14 1b 27 2a 32 39 38 54 61 7d 95 99 96 7d 6a 5a 56 50 5a 64 60 5c 61 5f 69 67 72 72 81 92 8b 95 97 99 9e a0 a0 a1 b0 a6 b6 b0 b5 be c6 bf ce d4 de de ea ed e8 ef f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f9 fc fa f0 f9 fe fb f7 f4 f5 f7 ed f2 e8 f1 ef ee ef e9 ea e5 df e1 dd e1 d5 d5 d2 d0 d0 cc be bc b4 bc be bd ae b4 a9 a8 9b aa 99 a1 99 94 99 8e 8a 8e 91 92 8e 99 88 8d 8a 88 8e 90 8d 8d 83 84 82 86 81 84 7c 7d 80 77 73 6b 6c 61 56 58 59 53 50 69 75 66 5b 3d 27 12 12 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 1c 15 20 2a 32 43 49 55 61 7c 8e 98 91 82 64 5f 61 55 5a 5a 59 5a 63 62 65 6b 70 73 75 7b 91 95 97 a5 a0 a8 ae aa ac a8 b1 b9 bf bf d0 c7 cb d3 d6 e1 e5 eb ed f7 f7 f9 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff fb f2 fb f8 f7 f6 f6 e2 ef e9 ef f3 e8 ee f2 eb ed e2 df e8 e5 df d6 da d4 d2 cc d4 ce c1 d0 c3 b9 c2 be bc ad b4 aa a4 a0 a5 9a 9b 9a 9c a1 9a 95 91 96 8e 8d 8d 92 8c 92 8d 89 90 8d 87 92 88 8c 85 88 8a 85 85 87 79 72 6d 66 5f 60 54 63 5e 5a 66 6f 66 48 3c 2c 1c 13 0c 05 06 01 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 06 07 15 17 23 27 2d 3c 4a 50 67 79 8d 91 88 78 69 65 5f 63 5c 63 60 65 5e 62 5b 61 6e 70 73 7c 80 8d 97 a1 a7 ae
 b2 b0 af bb bb c1 ca c8 c8 cb c7 d9 dc db eb e4 ef f3 f8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 fb f6 fd fc f5 ed f0 ed ef f0 e8 ef e9 e7 e6 ef e4 ed e0 de e6 dd da db d7 db dd d6 cf ca ca cd c5 c8 c2 c0 c0 c5 b3 b4 b5 ab ab ad ab aa 95 9e a5 9c 9f 9e 95 97 96 92 92 95 93 8e 97 8e 93 8c 86 8a 96 88 8d 8e 8c 89 85 6f 7a 6e 68 66 5f 60 54 59 58 62 6a 5a 4b 3b 28 24 13 07 08 05 00 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 11 12 15 25 2a 33 42 53 60 70 8d 9c 8b 72 64 61 5a 5e 68 64 5e 5e 5e 64 5f 60 63 75 6d 71 7c 84 8f 91 a3 a4 aa bb be be c7 c4 c7 cc cf cd d3 d6 dc da de e1 e9 f7 f0 f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fd fc fb f5 f4 f4 f2 f0 f2 f3 f1 ed eb e8 e8 e8 dc ea e6 df e2 dc de d8 db df da dc d6 d6 d3 ca d0 c6 bf c3 c3 be b9 bc b5 b6 b7 af ae af aa ad 9b 9c 94 97 9e 9d 9b 97 92 96 8e 89 96 90 93 8d 8f 92 93 8b 8d 96 90 87 89 7c 79 78 6d 69 67 65 60 61 56 52 59 5d 55 50 45 32 27 18 12 10 08 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 0a 14 17 21 1c 34 3e 4b 61 6a 77 97 a0 7b 6a 5f 64 63 5f 60 67 63 64 6a 6a 61 6a 73 75 78 6c 82 87 94 9a 9f aa b5 be c0 c5 cd d0 cb d9 d5 d5 dd e0 dc e3 e7 e8 ef f5 f1 fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f9 fe fb f7 f7 fa f5 f4 f7 f4 ec f1 f1 ec eb e6 e5 e1 e1 e2 e2 e2 e3 de d5 d4 d0 d1 cd cf d0 d1 ce c6 c6 c8 c9 c2 be bc c1 c0 b8 b4 bc a3 ae ac ab a9 a6 9c 9e 9f a3 9a 9d 99 90 92 91 8a 93 94 94 8e 8f 93 96 8e 94 8b 89 90 82 83 76 7a 74 6a 6b 62 61 5f 58 50 57 4f 58 57 4e 3a 32 1b 19 0b 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 10 1b 19 26 20 3f 4d 58 6d 72 8c 9b 90 76 60 5d 5d 60 5c 69 60 73 68 69 6c 65 6b 77 75 81 7e 8e 86 a4 ac a9 b9 c0
 b8 c4 d2 d2 d6 d6 db d2 da eb e6 e6 ee e7 f0 f3 fb ff fb ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff fa fd f9 fa f2 f1 ef ef ea f1 e6 eb ef e6 e1 df e5 e0 dd db d2 d8 d6 de d0 d6 d6 cd d6 d1 d2 cf cd c2 bf bf c5 c2 bc b8 bd b8 ac b3 b3 af aa a8 a5 a3 a1 9d a3 a2 a1 9f 91 93 99 94 91 93 95 8d 9a 90 93 8f 91 94 91 8e 8b 84 7a 7a 75 6e 6b 68 5e 60 5b 59 52 55 53 53 52 4c 37 30 2a 1a 13 05 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0a 17 14 24 2b 34 40 49 5f 6e 81 95 a1 8d 66 61 5c 5c 5e 5e 66 6b 66 6f 6c 6d 75 6b 74 70 80 7d 8c 8f 9a 9e ab b8 ba c7 cb ce d4 d5 d9 db df e4 df e3 eb ed f0 f4 f2 f7 f5 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 ed f1 f2 f3 ee f2 ee ea e7 ea e4 eb e4 df d9 da db d0 d8 d3 d6 d1 d6 d0 cd d2 ce c9 c8 ce c5 c2 c4 c5 bd bb b3 c3 b6 b1 b0 ab ab b0 a7 a8 a1 a3 a0 9c 9e a3 9a 98 95 96 95 8c 8d 91 96 94 94 9c 94 91 8d 8d 8c 87 81 7e 73 79 6e 71 68 63 5b 59 51 54 55 52 51 51 4c 47 3c 2f 16 0a 0c 05 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 12 14 22 27 2e 3d 42 4c 66 6e 8a 95 a4 81 60 5b 5d 67 5f 60 6c 69 68 69 70 74 6f 73 6e 79 84 88 8b 8c a1 a3 ae bf be cb cd d9 d1 d5 e0 e2 df db f3 e8 ea f1 e9 eb f5 f9 f7 ff fd ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fb ff f9 ff fd ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f2 f8 ed f3 f1 e9 e2 ef ea e7 e5 e3 dd e4 de d9 d7 d2 d2 d7 ce cf cc cd ce c1 c7 d1 c9 c5 be c0 bf b8 ba c0 ba c2 c0 b6 b2 ae a9 af b1 a6 a3 a2 9c a5 98 97 9b 9a 9c 94 9d 9a 88 92 8d 9b 9c 92 95 9a 91 8a 8e 89 89 84 7a 76 74 6d 60 64 5c 5e 61 5b 53 55 55 4f 5c 4f 4d 44 32 27 17 0d 04 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 0f 17 17 2b 32 36 48 49 5c 70 85 91 9d 95 6f 64 5d 61 64 68 5f 71 72 74 6c 7c 7b 77 79 75 81 86 85 91 97 9c a4 ac ae b9
 ca c8 d1 da d5 de df de e7 e4 ec ed eb f8 f7 f6 fe f4 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 ff ff ff ff ff ff ff ff fc ff ff ff ff fc f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f8 f2 f1 f2 f0 f1 ea ea ec e9 e3 e1 e0 e1 d4 d2 d4 df db ce d3 c2 c5 d1 cd c8 c6 cd c8 bf c3 be c4 bc bb b6 ba bd b5 b8 b7 ad ad b3 aa aa aa af a9 9d a5 9b 9f a0 a5 9d 97 93 99 96 99 9c 96 99 95 9e 9e 99 a0 87 8c 87 85 7b 7c 73 69 69 65 65 5e 64 55 5b 5f 52 54 58 5c 58 4f 44 29 15 0e 0e 04 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 12 15 1e 22 31 3d 4d 58 70 7e 87 a1 a1 90 69 64 62 60 64 66 6c 76 7b 78 7e 7f 80 79 7d 7d 80 89 8c 8d 8f 9c a6 ae b4 c0 c6 c7 c9 d2 dc d4 da e2 e9 ed ea eb ea ee ee f7 f9 f7 f9 ff fd ff fb f9 fd fc ff fd fa ff fd f8 fc f9 fb ff fe ff ff fb fe fb ff fd ff ff f9 fe f5 f6 ff f6 ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e9 f2 e8 e8 eb e8 e7 ed df e4 da dc e3 d4 e2 d0 d5 d1 ca c8 c3 cb ca cd cb c3 bf be bf c1 c0 bd be c1 b4 bb b5 b1 b5 af b0 ab ae a6 ad a9 aa a7 a7 9a a0 9f 9c 9c 97 97 99 95 94 95 99 9a 9c 9b 99 99 91 91 82 8e 7e 82 77 7c 72 66 61 65 5a 5a 62 5c 5b 53 58 5c 5c 65 60 5a 41 2f 1b 17 10 04 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 0a 0d 1b 25 35 38 46 4d 5f 6a 7e 92 9e a1 86 6d 63 5c 63 68 67 6d 7b 7b 81 89 87 8d 86 85 86 8b 8b 91 90 96 9b 9c ad b6 b7 c5 c1 c3 cb cf cf db df e1 e0 de e7 ea ef f1 f6 f7 fa fa f7 f7 fe ff fa fe fe ff f5 f8 f9 fd f7 fc fa f2 ff f8 f4 fe fc ff f4 fe fa ff f7 f7 f7 fc f4 ff f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 f4 f5 f0 f0 f0 e5 e8 df e5 e4 e4 db de d5 d2 d6 cc cd ca c7 c9 c2 c4 c1 c0 b7 bd bb c5 be bc b4 b7 b2 b8 bd ae b6 b0 ab ab af ac a8 a7 a9 a9 9e a4 a6 9c 9d a1 9e a1 9d 95 98 97 9d 9c 9d 9b 95 9e 97 8f 8b 89 88 8a 80 81 74 6b 74 64 6d 63 67 59 58 55 55 58 5c 57 5f 63 62 59 3b 2b 25 13 0e 07 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 11 17 1b 26 2d 3e 46 57 6a 7b 91 a2 a8 a2 78 6d 67 6d 6b 6d 68 79 7a 84 85 91 94 94 8f 96 91 97 94 8f 99 9e 9e aa af bb b5
 be c5 c8 cb d1 d7 d3 da de e4 e3 e8 ed f0 f1 ed f1 ec f3 f7 f2 f4 f4 fa f9 f6 f8 fe f9 f9 f9 f6 fc fa f3 f5 ed ee fd fa f7 f8 f7 f8 f9 f9 fa fc fc f2 fc f6 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 f5 f2 e8 f1 eb eb e6 e3 e5 e4 de dc da da d1 cd cf cd ca d0 cb ce c6 c4 bc c4 ba bb be be bd b7 b4 b7 b3 ad bb b3 b5 b0 b2 ad af ac ac a9 a6 a7 a9 a4 a6 a4 9d 9c 9c 9c 9b 96 9c a4 95 9b 9a 9d 8f 95 96 8c 8c 87 88 81 77 79 67 6c 6b 69 64 66 60 56 5d 57 5c 58 5a 59 68 73 76 65 52 3c 26 1d 10 06 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0a 14 21 26 31 33 3f 45 5e 6c 81 90 af a8 97 78 66 66 6c 71 71 70 77 7e 83 8e 8b 93 9a a5 9b a0 9b a3 a4 a1 a6 aa b1 b6 bc c0 c2 cb c9 cb d1 d1 d3 d5 d6 de dc d7 e6 ec e9 e6 e3 ec f2 f1 f7 f4 f5 f5 ff f6 fb fb f5 f7 ee f8 fd f5 f6 f4 f3 f5 f6 ef f3 ee f2 f9 f5 fb f1 f9 f3 f5 f4 f7 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 f0 f3 ef e1 f0 eb e2 eb db e1 e2 db d4 d2 cf cc d0 c9 c7 c4 c4 bd c1 c6 b6 bc bd b2 bb ba af af b3 b4 af b9 af af a4 ac b4 ae ad a6 ae b1 a8 ad a7 ad b0 a7 ab a6 9f a2 a5 a1 a0 a1 99 95 9a 92 94 96 8f 8f 84 87 89 8b 84 7a 72 6b 75 6b 64 69 5f 61 5d 60 59 5b 5b 5e 62 72 7c 73 5f 4e 38 2a 27 1c 10 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 1a 1f 2c 40 3b 53 64 7e 8d a0 a6 9f 85 6c 69 61 6b 6c 74 7a 77 7f 86 8c 92 a3 a2 99 ab a7 a4 a7 a4 af ac b5 bb b1 bf c1 cc c4 d3 ce d3 cf ce cc d7 d9 d8 dd dd e2 e6 e9 e8 e6 f1 ec f2 f6 f5 f0 f1 f3 f6 f8 f3 f6 f2 f4 ef e9 ee f0 f8 f3 f2 f0 f0 ec f6 f5 f7 f2 fb f2 f0 eb f2 ea fb fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 f3 f5 ed f1 e9 e4 e6 e1 e7 e5 da d9 d4 cf d3 cb cd c6 c7 ca c6 be c3 c0 bd b2 b5 b9 b6 b0 b1 b2 b6 ae b3 b1 b2 b0 b1 aa a9 ab ac ad ac a6 a8 a2 ad aa a9 ab a6 ab a9 a1 a5 9e a5 a1 9d 9e 9d 96 8f 95 98 8b 91 8e 83 7d 7e 84 75 6a 71 6d 6b 62 63 5c 5f 61 60 5c 5a 51 55 60 65 76 81 6c 66 47 45 33 2a 1e 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 16 1c 28 36 42 4e 59 6e 7b 8f a0 a8 94 7a 6a 60 68 70 78 78 78 82 81 8b 91 9a 9a a5 9d 9f a6 ad b2 af b2 b0 b5 b3 bb bf c1
 cd cf c8 ce d5 d4 cf d2 d6 dc d9 db e2 dd e7 e2 e7 e0 ee f2 f3 ef f5 f4 ee ef f2 f7 e6 eb e7 ea ed f0 f3 f3 ed e7 ee ea ee ea e2 f0 f0 ed f2 ee f3 f3 fa f1 ee f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec f0 ee f5 e1 e3 d3 e0 dd dc e1 db d6 d5 d1 cb c4 ca c9 c6 c3 b9 b6 bd ba b8 b0 b8 b9 b2 b6 b1 b5 b4 ab b0 aa b1 ac b0 af a9 ac b1 b7 ae ae af aa b3 b7 b4 b4 ab af a7 ab a4 a7 aa a6 9e 96 98 8a 86 90 91 93 93 89 7f 7a 80 7b 70 78 71 6f 6f 65 63 61 58 62 62 55 55 5d 50 5b 6a 7e 87 7e 67 5c 4a 3b 2b 1e 0f 0b 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 0b 08 15 20 20 38 43 52 5e 72 84 97 a0 a4 8f 7a 69 68 6f 72 77 73 77 7a 86 8e 93 98 9f a0 a6 a9 a9 b4 b2 b5 b3 b6 b7 bc c1 be c3 c6 cc c3 c5 cb d1 d0 d2 d1 d6 dc d9 db e4 d8 e6 e4 df eb ee e9 f3 ee f0 e9 eb f4 ee ef e5 ed e7 e4 e2 e5 e9 e8 e7 f0 e9 ed e8 ea f1 f0 ee ec ef f4 f0 f5 f4 f8 fc fe fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 ec ec e2 e9 e5 df d9 dd d2 d8 da d1 d0 d3 c6 cd c6 be c4 be b8 ba bc b4 ae b3 ae b3 ae b4 ae b5 b7 b2 af b2 b0 b6 aa ae af b9 b2 b4 a7 af b5 b1 b1 ac ae af aa a2 a8 ab a0 a5 a3 99 9b 8c 92 89 92 8e 85 8a 87 87 88 7b 7b 7f 70 6f 74 69 71 61 61 6a 5d 61 58 58 60 57 5d 5f 6b 83 88 7b 71 5d 50 36 2f 24 10 0b 06 07 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0c 1e 29 30 46 58 65 6f 84 99 9c 95 7b 6e 6a 69 73 70 70 6e 73 7b 84 8b 8d 94 9a 9c a7 ab af ad ae b0 af b1 bc be b5 b0 c1 c1 c2 c2 c1 c4 ce c6 d1 d5 cb d7 d0 d2 d9 d7 d9 e3 de e9 e4 e7 e9 e8 e4 e9 ec ec ea e7 e4 e8 e2 e4 e7 e6 e4 e4 f0 e7 ea f0 e6 e6 e8 eb ed f0 f1 f2 f1 f6 f4 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe e9 df e0 db de da d7 dc cc d5 cd d3 cb cc c1 c9 c0 bb b6 b2 bb b6 b2 b3 b1 b0 b4 a5 ac a8 ad ab b5 b5 b4 b2 b3 ae b2 b5 ad b0 ab ae b7 a6 aa a6 a8 a6 a2 a8 a0 a0 9d 9e 9a 9d 90 9c 90 94 89 84 87 87 8b 84 87 89 83 82 7e 78 73 72 6f 76 69 6d 62 64 57 62 5a 60 59 61 5e 5b 5b 68 87 89 79 73 59 47 39 31 21 19 0c 05 03 02 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 06 0e 14 1c 27 3a 46 55 6e 79 84 97 9a 84 6d 62 6e 68 72 7d 6f 79 7b 73 7e 78 8a 96 8e a3 9e 95 a1 aa ad ae af b3 b5 b4 b6 b5 ba
 bc bd bd bb cf c5 ca cd c8 d2 d3 cf da dd d9 e4 df e0 e4 de e6 ea e5 e0 ea e3 e5 e7 e0 e0 e5 e6 e4 e5 e4 e2 e3 e1 e2 e0 e6 e5 e9 ea ed e8 ed eb e3 e7 ee f5 f4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed e1 d7 da e1 d9 de d1 ce c8 cd cc c3 c3 c3 c5 b6 b1 b1 b4 b2 b0 b5 b3 a9 ac b3 ad ad b4 b3 b0 b8 b5 b9 b5 ba ae b1 a9 ac ac a8 ae ac 9b a7 9e 98 9a a4 a3 9b 9f a0 9c 95 94 9b 9c 8b 91 8f 8d 87 8a 8b 80 83 84 85 7f 7b 80 73 78 6b 6f 64 66 62 5e 5b 57 5b 5a 5e 62 58 58 67 69 8d 8f 85 72 59 5a 44 31 25 12 0c 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 05 08 06 17 21 1f 34 42 55 69 71 8a 9a 91 79 6a 69 68 70 72 73 72 6e 78 79 86 7d 8e 87 90 9a 92 9a a0 a8 a6 a7 aa ac b1 af b3 a7 be bc bb b6 ba c3 bf c7 bf ce ce d2 cb d8 da d9 df e2 dd e3 e0 e6 e8 e7 e2 e4 e5 e2 e8 e4 df d7 e2 e2 e0 de e7 e1 e4 e0 e7 e7 e2 e5 e2 e2 ee e4 e4 ec e7 f0 f0 ef fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e2 cd dc d7 d7 cb ce c9 cf c2 c5 c3 ba bc b3 ae b6 b5 b3 ae b3 b0 b8 b1 a7 af b1 b2 b6 ba b7 b5 b0 b5 af a7 a7 a6 a6 a6 a6 9d 9d a7 9a 9b a0 97 96 99 9a 9d 9f 8f 93 97 8f 93 8d 97 8b 87 8a 89 83 83 8d 85 79 82 7d 7b 7e 74 6c 6d 70 6e 6b 61 66 5f 5e 5d 60 5a 61 5e 5d 5c 6e 87 9c 85 78 62 49 3e 36 1e 13 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0e 0d 19 25 35 4d 53 6a 77 7c 8f 91 6f 63 65 6c 6c 6a 73 7a 76 7b 7a 83 7d 7f 8b 82 8f 8f 95 a3 9d a7 a7 a5 ab a9 b8 ae ae b5 b4 b1 ba c2 c4 be c6 c7 c9 c3 ce d2 d3 d7 d6 e4 de d9 d7 d9 e1 e0 de d8 d8 e0 e4 d6 dd da d6 da e0 dd df db dc d8 d6 d6 db dc de e5 e3 e1 e1 df ea eb f0 ea ed f0 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e7 d2 d1 d3 d0 c6 be c9 c1 be c3 c0 ba b8 b8 b3 b5 ab a9 ad b0 b3 af b2 a8 aa b7 b8 b6 b4 af b2 ad a9 a4 a3 a0 9c a4 9e 96 a0 a0 96 98 94 a1 8d 9b 95 8f 91 93 98 94 93 98 91 91 90 8b 93 87 80 7e 83 80 8e 7f 7e 7e 73 7b 77 75 70 71 6a 63 66 67 66 62 67 5b 5c 61 5d 5f 5c 75 8b 99 89 7b 5e 50 3e 2a 1c 11 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 07 0b 24 2d 35 45 57 6b 75 7e 94 8a 70 62 59 66 6d 6e 7a 6f 7b 7d 76 7f 84 7d 7f 86 92 95 93 97 95 a5 a5 a1 a0 9a ae a9 b5 b8
 bc ba b9 bb c4 c4 c8 c4 ca cd c8 dd d5 cf db dc d8 d9 da d9 de dd d7 da e1 db df db d9 d8 d9 dd db dd d2 d5 d9 db db de dd dc df dd e5 e0 e0 d9 e4 e0 e4 e8 ec f0 f7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 d9 d5 c3 ce bf c0 c1 bf be b8 b9 b9 af b4 a5 af b4 ae ad af b5 af ae b0 a9 b5 af ad aa ae ac a5 aa 9f a2 9e 9a 98 a1 94 a1 95 9a 93 97 9c 91 96 94 8d 8a 91 88 96 8f 8f 8e 94 97 91 8d 90 88 86 81 7c 84 78 80 72 6e 78 78 78 6b 74 6b 71 6b 67 66 6c 62 5d 62 5e 54 59 63 65 88 8f 90 77 6c 5b 42 3a 1f 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 06 0a 17 25 2d 3c 51 5a 70 7c 7f 86 7c 68 64 5b 69 69 66 71 70 73 7e 78 7c 82 83 80 88 8b 92 97 9a 99 a5 a3 9f ac ad ae ac b6 aa b3 bb b3 b2 c4 be c3 cd d2 c2 d4 d1 d4 d0 d4 cd d2 d6 d2 e3 df dc df e1 d8 de da d2 dc db db d5 d4 d3 db d6 da db d5 d2 e0 d7 de d9 dd de d2 db e1 db e6 e8 e4 ea ee f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff de cc bc c4 b8 bc b9 b1 ad b2 b4 bd b6 b5 a7 a6 a8 a5 aa aa a7 ac b4 a7 a5 af af b0 a4 a9 a3 a4 a1 9b a0 a0 a0 9c 97 9a 98 96 93 8d 96 91 8d 98 8d 94 95 87 91 8b 90 8d 95 95 89 92 87 88 86 7f 87 88 86 84 7f 7e 70 79 73 79 7e 6a 6f 71 68 69 67 69 63 65 62 69 56 5c 62 63 78 9c 8d 86 62 51 49 30 22 1a 07 05 06 05 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 0a 12 1e 26 33 4c 5b 6a 83 8a 82 70 61 53 5c 5d 64 64 6f 71 76 78 7c 6f 79 7a 87 8e 89 84 91 99 99 9e 9f 9f a2 aa a7 b4 b4 b0 b6 b1 b6 b5 c4 c4 c5 ca cb c5 c9 ce d1 d2 d1 d4 cb d8 d3 d4 da d9 d4 d6 d5 d1 d6 da dc d8 cf d9 d5 d3 d3 cf cd d3 ce ce d3 d6 df d9 dc db d5 d7 dc df e3 de e1 ea e5 ed ee f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dc cb b8 ba b7 b7 b4 bb ac a5 ae a5 af ad a4 ac a1 a1 a8 a1 a2 ad a8 a3 a5 ad 9f a2 a8 9e a2 9f a3 94 9a 9e 96 94 90 9a 8e 9a 98 90 9a 93 8b 93 8d 94 8d 8b 8e 8c 90 92 92 8a 8e 93 8d 87 82 80 82 7e 7f 81 7d 83 78 79 73 75 6d 74 72 6a 64 61 61 67 60 67 5b 5a 57 59 63 6a 79 92 91 83 63 53 4c 29 22 0e 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 07 11 1c 24 3a 45 61 75 81 7d 73 6c 67 5a 5b 63 64 65 5f 6c 71 71 73 7d 75 79 86 89 8c 8a 85 91 94 a0 a1 a5 a6 ab ac ac b7 af
 ba b3 b9 c1 bd c1 c0 c6 be ca cc ce d3 d0 d6 cd da d6 ca db d2 d2 da d4 da d8 d5 cf d5 d3 d7 db d4 d1 d5 d3 d4 cf cd d2 d0 d0 d4 cf d0 cf d0 ce d7 dc d1 de d8 df e2 e1 e5 f9 fc f1 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 ea df da c6 c5 d0 cd e0 e2 e1 fc ff ff ff ff ff ff ff ff ff ff ff dd c3 b3 ae b4 b2 af ad b0 ae b1 a8 a5 ac a3 a7 a1 a5 a2 ac 9d b2 a8 9f 9f 9a a0 a0 97 9a 98 99 a6 97 93 97 95 98 9a 9f 92 9b 8f 93 97 94 90 8e 93 92 8c 8b 94 91 90 91 8f 88 8c 90 87 8c 88 84 83 87 85 81 81 7f 70 76 72 70 75 6f 67 70 6d 66 66 67 5e 62 61 63 60 60 5e 63 74 86 8b 82 6c 59 40 36 1e 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 03 06 0a 0e 21 31 3c 50 64 79 83 80 6b 62 61 60 5b 5c 59 64 6e 69 67 72 6f 77 79 7e 7c 8c 8a 84 85 93 95 99 99 9f 9d a1 a5 af b6 b8 b4 b5 ba c5 c7 bd c1 c8 ca c8 c2 c7 ca cf d7 cd d5 d4 d6 d4 d0 cf d5 d0 d1 d7 cc cf cf d0 d6 d1 d1 d2 d1 d3 cc cc d4 d5 d5 cd c7 ce d1 ca d4 ca ca d0 d2 d2 d8 d7 d9 dd e3 e3 ec ec e8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dc d9 cc c0 c1 be b3 ad b3 bc bd cc db e8 f2 ff ff ff ff ff ff ff ff ff fc bd b2 af a7 b3 ae ab b1 a5 a9 ab a0 a5 a9 9e a6 9d a0 a3 96 a3 a1 9a 9a 9a 9a 9d a1 97 9f 96 9b 95 95 95 95 9c 98 8f 9b 97 9a 95 8d 92 8e 92 92 9a 88 92 95 8d 88 90 89 8f 88 83 82 83 8c 86 89 81 7f 7e 7f 77 78 75 72 76 76 77 6c 73 6b 6d 67 69 61 61 62 5b 59 63 64 66 70 8e 8a 88 6a 60 3e 38 2a 0b 0a 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0e 1c 28 3b 51 69 7f 8a 7f 70 63 5d 61 5d 5f 5c 63 65 6b 67 64 6c 70 79 75 79 86 84 8c 8c 87 8c 97 92 9c a4 a6 a9 a5 a7 aa bb b1 bc bb c7 ba c5 c4 c8 d1 d0 cd cc c7 cb d4 cf d2 cf cb cf cd d0 cc d8 d2 c8 d2 ca ca ce d2 cf d0 cc d0 ce cf ce c4 c8 c8 d1 c5 c0 ca c6 c5 cf c7 ce c7 ce d0 d2 cb d7 da e1 de eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e4 c6 b9 ac a6 9a 9d a1 9c 9d a2 a6 b4 c3 dd e4 f4 ff ff ff ff ff ff ff ff c6 b3 b1 a6 a5 a9 ab a6 a4 a8 a8 9b 9d a2 9a 93 97 97 9f 9b 9d 97 9a 93 9b 93 9d 94 99 9b 9a 94 96 91 90 8f 90 92 98 94 94 97 94 92 93 89 90 8d 8e 8c 8b 8d 91 8d 92 86 91 87 85 8d 8b 84 84 85 83 7c 80 7f 82 7d 79 77 74 73 74 74 70 69 6d 67 64 65 5d 5f 60 5e 5d 51 5b 71 8b 8f 83 65 59 3c 38 1a 10 09 05 09 06 06 05 03 00 06 05 03 00 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 03 0c 06 15 27 30 3c 53 60 74 85 83 66 61 5f 5d 64 69 6a 69 65 67 6d 6e 70 6d 75 75 76 7a 7d 81 8c 8c 97 97 9c 9b a6 a3 a1 ab ae a8
 ae b2 b8 bc b7 c9 bc c5 c8 cb c5 ca c3 cb cb c9 c6 c5 c9 ca d1 cd c8 c7 cb cb c3 c9 c5 bf c0 cc cb c9 c3 c4 c7 ca c6 c5 c6 c3 c1 c7 c0 c9 c6 bd c5 c3 cb c7 c4 c5 ba c7 d3 ca d2 ce df ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 d7 ce b6 ab 9f 97 89 8a 8b 8a 81 8f 8f 98 a0 b6 c4 d0 f0 ff ff ff ff ff ff ff c4 ab a0 9c a6 a3 a2 9e a2 9a 93 9d 96 92 96 99 95 9d 9b 8b 95 97 92 92 96 91 9b 92 94 91 90 93 98 91 93 8b 8e 95 91 91 8d 93 94 8e 93 8f 88 88 89 8c 8a 8c 8a 8a 85 88 86 86 87 8d 87 83 80 89 7e 80 74 72 75 71 7a 70 70 6f 75 74 6f 62 64 64 64 68 62 65 61 5d 5e 61 5e 72 87 8d 7b 6d 59 46 32 1b 06 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 09 06 0f 23 2e 44 4d 6a 71 7e 87 6e 64 5f 56 5c 63 6b 6b 6d 66 67 6a 74 70 6e 72 75 7e 80 84 81 8a 8c 98 9a 9b 9f a2 a4 a7 ac a9 ad ae ba b3 c3 bc c0 c3 cb c4 c7 c5 c9 c2 bd c9 c8 ca c6 c8 c3 c8 c9 cf c0 c3 c2 c9 c6 c9 c1 c7 c5 be c6 ca cd ce b9 c8 c9 c6 c4 c7 c0 bf b5 bc bf c2 c1 c5 c4 c0 c5 c9 c2 ca cd d1 dc ff ff ff ff ff ff ff ff ff ff ff ff ff f8 db cc c9 b1 9d 97 8e 7f 7d 74 6f 78 74 6d 74 84 8b 92 a1 b6 cb f0 ff ff ff ff ff ff ce ad 9e 9f 99 99 a2 98 9e 9b a1 95 9c 97 94 97 92 99 99 95 9a 93 8f 94 94 91 9d 90 95 95 9c 93 94 95 91 88 94 88 91 93 88 97 8f 88 92 8f 8b 88 8e 89 8b 90 84 8f 83 82 86 86 84 89 7b 84 80 86 7b 7e 79 7d 79 79 76 7a 6f 6d 73 67 71 6b 6e 63 58 66 63 68 63 5e 5e 5a 5c 73 7f 88 84 71 57 4a 36 1a 0b 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 08 00 09 16 23 28 3c 51 5c 6a 7c 82 67 68 65 5f 63 5f 65 64 69 71 69 68 6e 72 70 6f 70 6e 74 83 81 85 92 91 93 8f 98 9e 98 a0 a9 ae b0 ad b5 bc c1 bc c6 c1 c4 cc be c0 c5 c5 c5 c6 c7 cd c6 c5 c1 c4 bf c6 c5 c3 c0 c3 c7 c0 c6 c6 cc c4 c2 c6 c7 ca bf bc bc c0 c0 c2 b3 b7 b6 b7 c0 b9 b8 c1 bf c5 c6 c7 c0 c2 c6 c2 d6 ff ff ff ff ff ff ff ff ff ff ff ff e4 cc b3 a2 95 80 84 77 6a 6d 60 59 58 59 5d 5d 66 5f 69 73 82 94 ab cc f2 ff ff ff ff ff e5 aa a0 8d 95 94 9c 9c 93 95 93 91 96 91 93 91 92 98 94 96 91 8f 9f 92 93 91 9a 8d 8f 90 93 8c 8f 8b 91 94 90 8c 88 85 8e 95 84 8d 8f 88 8b 8d 87 88 8e 84 8b 88 86 85 83 8b 7f 88 81 7b 78 76 74 7b 73 75 76 6d 78 6d 6b 72 6f 70 73 61 6f 71 64 64 60 61 5b 5d 60 5c 64 63 8b 8d 7f 72 61 42 2b 1d 0d 08 05 03 03 06 08 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0e 1e 2f 37 4d 5a 72 7d 78 6a 5a 60 57 5d 64 64 67 69 69 6d 71 6c 67 71 75 6b 74 79 74 83 7a 8c 8a 8a 90 8d 97 9d 9d 9c aa
 a8 a9 b2 b0 b9 be b8 c0 c0 b8 bf c1 be c3 c2 c2 c1 ba c5 c0 bf c4 c0 be c0 c6 bc b5 be c0 b6 bb bd b7 c1 bc bc be bf ba bc b8 bb ba b3 af ad b5 ab b0 b5 b6 c1 bf bd b2 bb b6 be ba cd ee ff ff ff ff ff ff ff ff ff ff c8 a9 99 80 72 6f 59 62 53 59 52 54 52 51 47 4a 43 4c 4e 5c 60 69 76 89 9b bd e9 ff ff ff ff f4 a3 99 8d 90 98 95 93 8f 95 92 93 8f 92 8b 8d 95 8f 92 89 8c 8e 90 95 8f 8d 92 8e 88 88 90 86 8f 85 8a 89 8c 90 8f 8e 81 8e 84 86 8b 7f 8b 89 83 88 84 7f 87 83 85 81 7d 85 76 79 7d 7d 77 7a 79 79 70 71 71 6d 70 77 6c 73 71 6c 67 6f 67 63 5c 61 59 55 5b 59 51 58 62 68 7f 89 82 72 59 3b 23 11 10 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0f 24 24 38 4f 5a 6d 78 76 66 5f 5f 60 56 5b 60 65 65 6e 6a 69 74 71 6d 73 77 79 79 81 81 82 89 80 8a 8e 95 94 99 96 9f a0 a7 ab a7 b4 b8 b2 b9 bc ba bb be bd c1 bc bc c5 c4 be c4 c2 bb c4 c3 bd c2 b2 bf b4 ba b9 b6 ba bf b8 bf c1 b7 bc bc b9 c5 b5 b5 b4 ad ad a3 ac ae a9 a8 b1 b4 be b6 b5 b8 aa b4 b9 bf da ff ff ff ff ff ff f9 ef e8 c3 9d 83 77 64 5e 57 56 57 4c 4d 41 41 49 46 44 4d 44 49 50 53 55 54 5c 69 78 90 b6 e9 ff ff ff ff a2 93 8b 94 93 91 99 93 90 93 92 91 8e 92 8d 88 8a 95 8c 8b 8d 91 98 8a 89 97 8e 8f 8e 8d 93 8e 84 88 8c 8e 84 88 88 85 82 8c 8b 8b 87 89 81 83 8c 8a 82 89 81 80 7b 7a 80 77 7c 7d 7b 76 7e 70 78 72 75 77 6e 77 6b 6d 68 6f 6d 6e 6d 68 64 60 5c 5e 56 59 59 52 56 63 6c 7f 85 82 6d 56 40 32 10 11 09 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 06 06 15 1e 2b 3b 47 5a 6f 6e 7a 60 5c 66 5f 58 5e 62 5c 6a 6a 67 6e 6e 73 70 73 75 75 7f 78 7e 82 7f 84 8b 8e 8e 9c 92 98 97 9c a6 a9 a9 ad ad b3 b5 ae b4 b9 b5 bc bb c4 bd c4 bc b2 bf bf b5 b8 ba b7 be bc b2 b6 b8 b4 b9 b6 b7 bf b6 bd b0 b9 bf b5 ba b8 b6 b2 b0 aa b0 ae ae ad b4 b4 b3 b0 b8 b0 b0 b4 af b4 bc d4 ff ff ff ff ff fd d6 c3 b3 9a 7b 64 55 50 49 4d 48 4b 4b 45 3a 3d 3d 41 40 3f 3f 3e 44 43 4f 50 50 59 5c 70 92 b9 fc ff ff ff a4 89 85 8d 92 8e 9a 8a 8f 90 87 8e 8b 91 94 8f 8d 89 8d 91 89 8a 86 8e 86 8e 8a 86 8b 86 8d 8f 8a 8c 8b 8d 8a 8b 85 88 90 8b 86 89 88 89 8c 82 89 80 7e 83 7b 7a 7d 7a 7c 77 7a 84 73 72 78 77 79 70 70 74 6f 71 77 71 70 6d 6d 69 68 66 69 67 57 5f 5f 5c 5e 61 56 62 6d 7d 85 83 6d 58 37 1f 17 0d 06 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 16 2a 35 4a 62 67 70 62 61 5d 55 54 5a 60 56 5c 61 61 65 64 71 71 7b 75 72 78 7d 79 84 7d 7e 89 8a 86 8a 90 93 97 97 9c
 a6 9e a9 a3 a4 ae aa b3 b7 b5 ba bb c0 b9 bc bf b7 b7 bc b6 b3 bb b6 b9 b2 b4 b9 b3 ad b9 b5 b4 b2 b5 b7 b7 b6 b6 b9 b6 b9 a9 a4 a9 a5 a7 a2 aa a4 ad b0 b0 b0 ad af 9f ac ad a1 b0 af c7 ff ff ff ff ff e5 ba 9d 8d 7a 63 53 47 45 48 44 3f 3d 3e 3d 39 38 33 34 36 3c 27 31 37 36 3f 42 3c 43 4f 59 6a 93 c8 ff ff ff a5 8a 84 84 8a 8d 97 95 8f 8a 8a 84 88 85 84 87 8e 87 87 8f 8c 89 86 8a 8c 88 8d 88 8a 8a 89 84 86 83 8a 8c 89 83 8e 8b 86 85 86 84 7d 84 85 7d 8b 83 77 7f 7a 79 76 78 7c 73 75 75 6d 72 71 73 7a 78 73 73 65 6a 75 69 72 6b 6b 6d 62 6b 5b 62 60 60 5b 4f 5d 60 62 5e 6b 73 80 7a 66 52 3a 29 1e 10 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0f 1c 23 42 4c 5b 69 6a 5d 5e 5c 57 5d 5d 5f 58 5c 60 5f 69 65 6e 73 70 78 72 76 7a 75 7d 7e 7d 82 89 84 8b 96 8e 9b a0 9a 9f 9c a4 a5 a5 a6 ae b1 b2 ae b7 b8 b3 b7 b3 ba c1 b4 b6 b2 b0 b6 b8 b4 b3 af af b5 b9 b2 b2 ad b5 ba b2 b9 b0 ad b1 a9 ad a5 9f aa a1 a9 a5 a0 a6 ad a9 ab a0 a2 a2 a6 9e a5 a7 a6 b3 bf e7 ff ff ff ff da b2 91 71 58 50 4f 4c 3e 3d 31 37 34 2b 2a 2a 2a 1f 2f 29 2b 30 2b 2a 32 35 42 45 41 3f 49 54 70 a3 eb ff ff a9 89 80 86 88 98 90 91 8d 8e 88 91 8a 8f 8d 8b 8f 8b 8a 88 86 90 85 86 86 88 81 8d 90 8a 89 88 7f 85 88 84 8b 7f 78 8a 8c 82 8d 84 85 7e 85 89 7c 81 7d 74 78 78 76 75 77 67 72 78 6c 71 77 6c 73 6c 74 72 6b 6f 6d 6d 6e 6b 67 6b 64 5f 67 5b 60 57 52 60 57 5c 60 67 6a 6a 82 7c 68 55 3e 25 23 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 05 00 0a 0e 1d 25 3d 47 5a 66 65 5e 53 58 5b 54 5c 59 5a 5a 62 66 66 61 6b 70 72 75 78 7d 7f 84 81 85 78 7d 7a 80 86 8e 93 93 95 98 a2 9b a1 a1 a3 a1 a6 ab b0 b1 b1 b4 b2 bb b6 b0 b4 aa b1 b4 b0 af b2 b1 a9 ae b5 a3 ac b0 a5 b9 b5 b2 b0 ba b2 b1 af ab af a6 ab a6 9f a0 9a a7 9d 94 9f 9d a3 a6 a2 99 a3 9f a2 a1 aa b1 d2 ff ff ff ff c3 91 77 5c 50 4a 42 3c 2c 32 27 2d 28 20 26 20 29 25 22 21 27 1d 2b 29 2f 2a 31 35 39 39 44 50 6a 85 c7 ff f8 a9 8e 85 8c 8b 8a 93 87 8a 91 8d 89 86 8a 8f 84 88 86 87 90 8a 8c 8b 8f 7d 8b 7f 79 7f 82 83 89 85 8b 86 87 83 85 86 83 8a 82 84 84 84 81 85 80 7d 7d 7b 7c 75 70 78 6f 75 79 76 80 71 6d 71 78 6c 77 71 6e 6a 71 6d 73 6a 6c 69 6d 63 62 64 52 56 5d 51 58 62 5d 5e 5e 5f 62 7a 7d 65 56 37 26 13 11 0d 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 12 06 0e 20 23 36 47 5a 67 5e 57 53 4f 59 50 55 55 54 5f 62 62 62 65 63 6a 75 75 7d 85 7e 81 83 86 84 80 7e 85 89 88 89 87 92 88
 9a 99 95 9c a0 a1 a8 a6 a7 ae aa a5 ac af ae af b7 b0 aa a9 b1 aa b1 af b5 b1 a6 ab a8 a7 a7 a6 a6 a5 af ba b1 ae b0 a7 a2 a2 a0 ab 9f 94 9b 9b 9a 9f a2 99 9a 9c 9c 9b 9d 9f 9d a5 9e ac c1 ff ff ff ff b0 8a 64 4c 41 47 35 30 28 2e 2b 20 23 1b 1e 16 1a 1b 20 1b 1e 1a 1f 1f 24 28 1d 24 25 31 3a 48 52 77 a8 ea e4 a0 89 86 85 89 88 8a 8f 8a 88 85 7f 88 7f 8d 84 82 8c 88 82 85 87 84 85 86 84 84 7b 7b 83 7f 84 84 84 7f 80 7d 7f 8b 83 89 7f 81 84 83 7f 86 7c 7b 7c 7a 7d 78 72 75 73 6e 74 6b 6c 6d 6c 74 60 69 67 70 6d 67 6c 6b 65 6a 6e 6f 6a 65 5d 60 59 5a 5c 5d 58 55 59 5f 56 5f 63 78 79 61 48 39 1c 17 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0d 08 16 1a 30 33 49 58 67 65 5c 52 4b 4d 56 55 5b 5a 59 5e 62 65 67 65 70 70 74 70 80 7c 84 7c 84 83 83 84 83 86 88 87 8d 9b 96 97 94 95 93 9d 9c 9b 9f a3 a1 a3 ae a9 a7 ac b2 b3 b2 a4 ad a1 aa b0 a8 b0 ad a3 a5 ac aa a9 a7 b3 ad af ad b1 a9 ab a6 a2 a0 a3 96 9f 9f 93 9c 93 8f 9a 97 99 9d a2 9d 9b 9c 9a 9b 9d a7 b9 eb ff ff ea 9b 77 56 49 40 2f 26 23 2e 21 18 19 20 20 1a 13 17 17 13 14 11 1a 1a 21 17 18 20 25 25 2b 28 36 4f 6a 99 d0 cd 9d 96 85 8a 8c 86 95 89 8b 89 8c 88 85 8a 82 8a 8a 8a 8b 84 81 86 80 7c 79 8b 83 82 79 7b 7a 7a 84 85 80 86 7e 7d 7d 7e 85 7f 7f 7e 7f 7d 7b 76 7f 79 77 7e 78 82 75 7b 74 6f 72 6b 6b 6f 6d 6e 72 61 69 66 63 6a 67 6f 73 6f 6a 6a 6d 60 57 5e 55 58 5a 5b 57 61 60 68 5f 66 70 78 5c 50 37 24 1c 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 05 03 0b 0f 17 1e 21 3c 46 59 69 65 55 48 4f 51 4c 52 5a 54 5d 5d 63 63 5c 61 66 68 73 78 7a 83 87 87 86 92 8d 87 89 8d 8a 83 90 8e 8c 8c 8e 96 95 98 9a 9f a5 a1 9f a7 a6 a4 a7 aa a8 ab af ad ad ac ac b0 a7 ab a1 a9 a7 ac a7 a7 b0 a6 af a8 a7 ac a0 9b a0 a8 9e 9b a0 9b 99 94 92 9b 92 92 99 9b 9a 97 96 a0 99 97 96 94 a0 a8 cb ff ff d9 9b 64 54 41 34 26 27 14 1d 19 1a 1c 1a 12 17 18 1a 16 19 14 13 18 14 16 16 16 14 1e 29 2a 24 2e 44 66 85 c2 be 97 97 89 84 89 89 8d 88 85 8c 89 83 87 8a 85 84 85 8a 85 89 83 80 7e 80 84 82 81 79 7f 75 7c 81 7a 83 7a 7c 86 7e 7a 87 87 80 7c 84 7e 7c 76 73 73 78 79 74 76 74 76 74 6c 72 76 73 66 74 69 6a 67 6d 6b 68 6f 65 67 70 75 70 72 67 5c 5f 60 56 55 54 62 60 65 66 6a 6a 67 69 75 7a 62 4c 3b 2b 26 0d 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 1c 26 2c 33 49 59 6d 5a 53 53 4e 4c 4a 53 4e 53 4e 53 5d 5f 59 62 60 66 70 71 72 7c 80 7a 7e 90 8b 90 90 8d 90 90 8a 92 8f
 96 90 90 96 96 96 90 9a 9a a1 a5 ac a2 ab a4 aa ac a4 a5 aa ad a6 a9 aa a8 9d a5 ab a6 a9 b0 a4 a8 a2 9d a8 a1 98 94 98 94 90 96 91 8d 8f 93 90 8f 94 8b 93 92 98 95 97 98 93 9a 9e 9a 9e 9c aa ee ff da 99 5f 4e 34 21 22 18 15 16 0a 13 0a 0d 0c 10 09 13 12 06 0c 14 0f 12 16 09 18 1a 1b 1e 18 19 24 40 5e 85 b5 a5 93 8d 88 89 85 91 8a 86 80 80 7e 89 89 8c 87 84 88 80 82 8c 80 81 7e 75 84 84 88 75 79 83 76 81 70 77 7a 7c 78 82 7e 81 82 7b 7d 7b 80 7e 76 75 78 79 78 73 72 74 72 74 6c 69 6e 68 65 67 6d 6f 61 65 67 64 66 5f 68 66 6e 6a 70 6f 5e 60 53 56 59 5f 59 63 64 69 6a 6a 66 66 6d 79 62 51 3d 28 1b 09 14 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 0d 0b 14 24 20 3c 4e 57 69 5a 52 51 47 4b 4f 50 58 57 56 5b 59 58 5f 5f 5f 65 65 6f 73 77 7f 86 83 89 8b 91 92 95 a3 8e 93 96 8c 94 8f 90 92 96 95 9d a1 a2 9c a4 9f a6 a2 a9 ab a9 a5 a5 aa ab a6 a4 9c a8 a3 9b a5 a0 a5 a7 ac a6 a0 9c 9d 98 8f 8a 96 94 8e 93 95 8c 8f 90 8e 8e 8f 89 94 92 8f 96 93 99 90 9d 9d 9a 98 9e 9d c9 ff ea 94 61 55 34 22 1e 19 11 0f 0c 15 0b 0e 0d 05 0c 0f 0d 0f 0b 0c 07 09 07 0d 0e 10 13 0d 1f 1f 1f 2f 57 81 a7 a2 97 8b 88 90 84 87 8a 86 89 84 83 7f 8c 8b 85 8b 83 8d 82 87 7d 7f 7f 84 85 7c 7a 7b 78 7e 79 82 7d 76 80 7e 75 7a 7f 84 83 79 84 70 76 7a 74 75 70 79 75 75 76 78 75 6d 6e 63 6d 6d 6f 6e 72 6c 60 74 5e 68 5b 63 68 6a 73 6a 6e 69 64 5f 59 54 59 52 5d 64 64 67 70 72 5c 5e 6c 70 62 55 3b 2b 1c 15 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 05 16 18 1f 2f 38 46 5f 65 60 5a 56 4e 50 4d 4e 50 54 4b 57 59 5b 58 5a 5e 62 66 65 6a 72 78 7e 78 82 85 8a 8e 8d 9d 94 90 96 98 97 92 9b 9a 92 99 95 a0 a8 9c 9e a0 a1 9c a8 a9 ac a6 a5 a7 a6 9e a3 a5 a1 a4 a4 a3 a6 ae aa a2 a0 9c 98 9a 98 8b 90 8e 90 90 96 86 90 89 8a 92 8d 8e 8a 8c 8a 94 97 94 97 90 94 96 97 9b 96 9e b2 ef ff a6 66 42 2e 1b 13 1b 16 14 0f 05 08 0a 0f 0e 07 09 0f 0e 0a 13 0c 09 09 11 0f 15 17 22 17 1a 14 2d 4f 89 a9 a0 93 90 84 8b 82 85 8d 84 80 83 83 93 83 86 89 81 84 86 8a 88 89 85 85 81 7f 7f 7c 84 7d 72 76 76 79 73 74 7a 6e 74 79 78 83 76 72 7a 7a 73 72 77 73 71 75 73 6c 76 76 72 70 6a 74 6b 69 6c 63 66 68 66 6b 6e 5e 6e 61 62 66 70 72 6a 5f 64 5f 62 63 5c 61 64 67 62 67 67 67 61 6d 77 62 60 43 2f 23 0e 11 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0e 0d 22 2d 34 56 62 69 65 55 51 4f 51 4d 4f 52 51 52 54 55 51 54 58 60 5e 62 67 65 68 70 71 7c 82 82 87 90 8a 95 8f 95 97 9e
 99 94 96 97 93 9c 9d 97 9e 9c 9f 9c a3 a0 9f a3 9f 9d a8 a7 a3 9f 99 9a a1 9f a7 a2 aa a9 94 9a 9b 97 88 8e 85 86 85 8a 96 89 8e 88 8b 80 8f 8f 8e 8f 8f 88 8c 8a 8c 94 8f 8f 8b 91 93 98 9b 99 a4 bf f6 c0 70 4d 2d 1a 10 10 06 09 09 07 07 08 03 0f 0d 05 0a 02 06 05 08 0c 06 05 08 10 0b 1d 13 0f 12 25 59 85 9c 93 8c 8a 8a 84 80 8a 81 83 7d 8e 86 85 8f 88 84 86 87 7d 82 84 83 80 7e 84 83 7e 78 7c 78 79 75 7a 77 78 73 76 75 78 7c 7b 75 7b 7e 74 6d 74 70 75 78 72 6d 79 69 74 6b 74 79 6e 6a 66 66 6a 65 61 66 67 68 65 67 61 62 61 5f 60 67 60 65 5f 60 60 67 62 5e 65 60 5d 5e 58 5c 61 72 7c 69 5d 49 32 17 13 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 1b 22 2e 38 50 5c 64 6d 5b 53 56 50 50 4e 4d 4a 49 54 52 4c 52 54 53 59 5e 62 61 6d 6c 68 77 7b 81 82 7f 83 8b 95 88 95 98 99 93 9a 9a 97 98 9e 94 99 94 a0 a1 9a a2 a3 a3 a3 a0 a4 a4 a1 9b 9b a0 a2 90 9d a1 a6 9b 96 99 8b 8b 85 8d 89 89 83 89 88 7c 82 7f 8f 83 86 83 8f 89 89 87 81 86 88 88 8a 8d 8d 96 8f 9d 99 99 96 a3 d3 c6 75 4a 28 12 0a 07 0f 06 08 02 06 05 05 06 06 05 04 03 06 05 03 07 07 0a 0d 06 0d 0f 13 0e 11 1e 54 91 96 98 93 8e 8b 8e 82 84 84 89 87 8f 8a 87 85 7d 8b 82 84 85 82 84 8c 7b 82 7a 79 7b 7a 7f 78 74 74 71 72 7a 72 77 74 77 74 7c 7a 72 75 7a 6e 6f 72 71 68 6c 75 6f 74 6d 6e 71 73 6a 70 6e 66 64 65 62 61 61 61 5d 61 62 5d 5e 5d 63 5e 63 5e 59 53 5b 5e 59 5c 55 4d 54 56 61 5c 54 6c 73 6d 5f 3f 2e 23 07 0c 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 07 09 17 1a 2e 44 49 62 68 68 60 51 53 4f 54 51 50 49 4c 46 54 52 54 58 5a 57 5b 60 60 65 6e 74 6f 77 7c 85 84 82 86 8e 8f 9a 9f 9c 9c 97 9d 9e 9b 92 9c 98 9d 9e a4 9f a0 a2 a5 aa a7 97 9c 9d 9f 9c 9b 9d 9b 99 9f 9e 90 93 92 8a 89 87 8a 84 7d 87 85 90 87 84 7b 89 8f 83 89 8c 82 87 87 85 82 83 8f 81 8d 8a 85 8b 96 96 97 a1 a1 ac be 82 49 2e 14 11 04 06 05 03 03 0a 0d 07 04 0b 05 08 09 07 05 04 06 08 0a 03 00 08 13 16 13 1b 1b 4a 7e 92 96 93 90 90 8f 85 8b 84 8a 80 84 8d 88 7a 80 81 84 84 80 7e 89 76 7c 84 84 7e 78 80 72 72 75 73 76 71 76 70 75 76 6b 73 70 70 74 79 73 79 6a 69 70 74 71 72 75 6f 71 6e 6d 74 6d 70 64 6a 67 70 6f 60 64 5d 64 5e 67 68 69 66 65 51 5a 4f 50 58 56 53 58 56 56 55 51 53 57 55 59 6b 7f 73 66 45 31 25 18 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 07 0d 17 20 28 3a 53 66 76 66 5f 57 59 57 50 4c 52 4a 52 52 4d 50 53 51 57 53 5e 61 5f 68 64 6c 6d 6b 79 81 7c 85 93 8d 90 90 98
 98 9a 9f 9b 9f 99 98 9b a0 a3 a1 9e a0 9f 9d a0 9e a0 9e a4 9d 9c 9c 95 92 9b 95 94 9a 91 8a 88 87 88 83 83 79 80 83 7d 88 81 88 86 81 82 83 79 86 7d 82 8b 83 85 88 85 89 8f 89 8e 91 8f 90 93 96 9a a8 a4 8e 50 30 12 06 0a 0c 05 09 01 06 0b 03 01 06 05 03 0f 0a 09 03 03 06 05 0f 10 0b 13 0e 10 11 1f 48 7c 96 91 98 96 8f 88 8b 83 89 83 87 8b 82 88 88 83 8c 83 85 81 81 83 7d 7e 7b 84 73 7c 77 76 77 78 73 76 77 79 72 6b 71 65 72 7a 75 6f 76 71 74 6a 77 69 6f 6d 72 68 73 74 6a 77 6f 6c 71 69 63 69 64 64 62 6c 62 5f 62 6b 6a 66 62 65 5a 5a 4d 54 50 54 56 4f 55 59 58 5c 58 54 59 56 65 7c 72 64 4f 45 28 11 09 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 08 14 22 2d 4a 52 64 64 66 57 51 5a 58 54 55 48 47 46 52 4b 4d 58 4b 4e 51 51 5d 59 58 64 63 66 74 75 79 78 75 84 84 8d 90 93 8f 8e 92 95 99 98 99 9a 8c 94 94 9e 92 9d a4 9c 9e 9f 98 9e 9a 96 96 95 94 8e 98 98 93 90 8a 84 8d 7a 79 76 78 78 7f 84 82 8c 82 82 80 89 7c 83 82 83 7a 83 7f 88 7d 8e 87 86 87 90 8b 9e 93 98 9d 97 9b 9a 7f 4e 34 12 05 06 08 05 03 03 06 05 03 00 06 05 03 01 06 05 03 07 06 05 07 00 07 05 0a 0f 10 21 47 77 94 95 9b 9e 98 95 8e 84 85 85 84 89 87 8c 84 85 80 82 81 7f 81 83 7a 7c 7e 7c 7e 7c 72 76 73 78 7a 69 71 6e 76 73 6a 66 6d 6c 6f 70 6f 76 67 69 65 74 72 69 6a 62 6b 70 71 74 6f 6c 72 63 65 5d 66 65 64 68 60 68 63 5c 63 58 59 5b 59 56 56 4f 51 53 4e 49 56 50 59 50 5b 54 59 52 62 72 72 6f 53 42 24 17 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 05 08 13 12 24 32 3d 50 5e 70 69 65 55 5c 5c 5a 4e 4f 4f 52 4e 58 4a 4d 49 55 51 5b 55 5e 5f 64 63 63 6a 6a 7c 7a 77 84 81 8c 8e 8b 98 96 8d 95 96 96 98 9b 98 9f 96 9a 9a 9a a0 9c a3 9f 93 a0 98 91 95 91 93 90 8c 98 93 90 88 82 81 75 7b 7a 7f 78 81 80 7f 8a 7a 7f 7d 77 85 82 7d 86 81 84 80 82 82 84 84 89 91 84 8a 90 8e 93 9a 99 93 96 87 57 34 1c 08 07 06 05 06 06 07 05 03 00 06 05 03 01 06 05 03 05 08 05 03 06 0b 05 0b 11 0b 21 42 7c 99 96 ad ad 9b 94 89 8d 8b 8c 8d 84 86 83 84 80 87 86 83 86 7e 77 88 7a 7e 82 7f 82 72 77 79 6f 70 73 73 73 70 74 6d 6e 6f 70 7b 73 6f 73 67 6b 6f 74 6b 72 74 70 6e 6f 73 6c 69 66 6b 6a 68 66 67 66 60 60 61 62 65 60 64 56 56 50 52 56 54 50 4f 52 51 51 53 5c 5c 56 5e 56 52 51 62 75 79 69 56 43 2b 1d 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 01 0c 14 1d 30 42 5a 62 76 65 5b 5f 53 54 56 50 5b 4f 51 4e 4f 59 4b 49 52 59 57 60 5b 5e 67 61 64 69 6e 78 73 7f 84 7a 87 90 89
 97 95 94 94 97 92 96 97 94 a1 93 95 9b a2 9e a2 99 a0 95 99 97 9a 98 92 93 89 8d 93 8b 86 89 87 74 7a 78 7b 7d 7c 79 7d 88 79 85 7f 7d 81 79 7b 83 88 7d 7e 86 81 80 89 84 81 88 84 8c 94 95 9c 95 9d 9f 95 7f 5f 3c 13 0d 09 06 05 03 07 09 05 03 00 06 05 06 00 06 05 03 00 06 05 03 06 09 0b 10 08 0c 1e 48 84 9c a9 af a7 98 8b 8c 8d 8d 8d 85 91 86 8c 8d 89 84 8c 81 8a 85 81 7d 7e 7c 82 7f 79 75 71 7a 74 71 6d 6e 6f 70 71 6a 70 6e 73 73 6b 72 72 63 69 6c 6c 6e 71 6b 74 71 70 72 70 72 6e 69 6a 62 61 6a 60 5d 5f 62 6f 5e 57 57 57 58 57 50 53 52 4a 49 56 55 51 56 53 54 57 55 56 5a 5d 62 72 7b 6f 5f 41 35 10 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 18 22 32 47 59 6a 67 6d 59 5c 4f 56 5a 50 58 52 50 58 50 57 4f 4c 4d 4d 5a 5c 5b 61 5d 61 65 61 67 66 71 75 75 7c 76 88 85 8f 92 98 91 8d 91 98 97 9d 9f 96 9a a0 9a 9e 9c 95 9b 97 93 8b 95 90 93 8c 8a 8b 8a 85 85 89 7d 7e 78 73 7c 7a 7a 7d 7c 7b 83 7c 7e 7b 7d 7e 82 81 7f 7d 81 7b 81 86 86 88 7a 8b 8c 8d 91 8d 91 92 9c 94 9b 86 5f 3f 0d 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 0a 06 08 0c 09 11 15 3f 7e 95 a4 ae a7 8a 90 81 8f 92 91 89 8d 84 85 88 88 7e 7d 87 7e 80 82 77 77 7c 74 78 78 71 77 7b 73 6e 71 6b 67 6d 6d 6d 6b 6e 70 66 6f 69 6a 6c 6d 62 6a 66 6c 71 72 67 66 64 76 6c 6d 71 63 62 62 60 66 64 66 64 64 53 51 54 4d 59 50 50 5c 4b 50 53 4e 4e 53 51 55 5d 54 65 57 5b 5b 62 7c 73 6f 65 47 2a 19 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0b 0f 1e 32 45 54 67 73 6f 5f 52 51 4e 53 59 54 56 4e 59 51 54 54 52 4f 50 4f 57 57 5a 62 59 62 65 6a 72 72 79 7d 77 7d 85 86 89 89 8d 93 91 9c 95 98 92 92 96 96 97 9b 97 92 95 94 9a 9d 92 92 96 87 96 89 8c 8d 8b 88 83 82 76 74 7d 75 7c 7a 78 80 7f 7e 85 7f 7e 79 7c 7e 7e 76 7e 7f 7f 7f 7e 79 7e 8b 86 8a 85 8d 96 94 8b 95 92 91 87 68 44 16 04 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 02 06 05 03 07 08 08 03 06 0b 1d 46 81 91 99 9c 93 86 8d 8c 8b 89 85 91 8f 85 82 81 87 82 87 7e 7b 71 7e 82 75 78 79 75 70 69 72 69 75 70 70 6d 68 6a 6d 6e 61 66 6e 68 63 6e 67 5f 65 73 64 71 74 6d 6c 68 6f 78 6a 6a 63 64 64 64 66 66 65 5a 60 64 62 5e 55 60 4d 55 52 59 52 4e 53 55 5c 57 5a 4d 52 55 5e 5b 5a 57 54 64 6f 77 77 5e 4f 36 1f 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 05 03 08 08 19 21 2d 45 60 68 74 72 61 4d 56 54 56 56 57 5e 53 51 5b 56 55 50 51 57 5a 5d 55 5d 5c 5c 60 63 6b 6a 6f 7c 77 84 77 80 87
 88 8a 8e 93 9a 8b 96 90 96 94 96 96 92 9b 8d 96 93 95 9e 91 92 99 98 89 8c 8c 85 88 8b 92 84 85 7b 76 76 7e 79 7d 84 82 85 7f 83 7b 7b 7b 7e 7b 83 73 80 7e 7c 84 81 8b 87 85 8a 8a 7f 87 91 93 90 97 97 88 82 65 49 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 0b 0a 05 09 06 18 3e 74 8f 9b 95 91 87 8e 8f 8d 8e 8d 8f 8f 84 7f 89 8a 82 82 7a 7c 7a 7b 7b 79 76 75 7a 6f 79 71 71 6f 73 6d 6b 6e 6b 68 67 67 67 6c 6b 71 6c 6f 68 64 70 66 70 6e 66 6c 6a 78 75 74 72 6b 6b 67 66 60 65 67 56 6b 5d 5e 5d 5a 51 57 53 5b 54 55 51 56 4d 4b 4d 55 55 55 55 51 5f 54 55 53 59 69 7a 72 6b 56 3d 20 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 06 06 0f 1f 2c 41 59 66 70 70 56 4e 53 49 51 51 51 54 58 53 51 51 4b 44 49 53 59 61 59 59 56 58 5e 5e 62 68 65 76 75 70 80 7d 82 87 8a 93 8c 8c 91 90 94 9d 90 99 96 92 90 8b 98 8d 91 8f 91 8a 92 93 89 8b 84 89 88 91 89 84 84 81 7a 79 75 7e 72 70 80 7b 7c 84 81 7e 73 7d 7c 75 77 77 7c 73 80 79 75 7e 7e 83 7f 8b 8f 92 91 97 9c 92 8d 7e 61 40 0f 0c 05 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 07 06 0a 14 39 79 9a 9b 94 91 8c 8f 8e 8a 8a 8a 84 8c 86 83 81 7a 81 7f 7f 7a 76 7a 77 73 76 76 77 75 76 6a 6c 74 73 6d 60 68 68 5f 5e 67 5f 67 67 66 62 6a 61 63 6a 65 6b 6e 72 71 71 6d 79 6b 6e 6d 65 64 64 67 64 5a 61 5e 65 62 51 5c 4b 57 57 54 5d 50 4d 50 51 54 52 52 59 5b 58 53 51 5b 58 58 58 65 73 73 69 51 3b 1f 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 06 0b 12 25 32 4c 5c 6e 74 76 63 52 55 4e 52 52 56 5a 55 56 56 50 5c 4d 50 52 54 56 52 5d 5c 5b 60 67 6a 69 68 72 73 76 7c 80 7e 86 88 8b 87 94 93 8e 8e 93 95 95 94 90 92 8d 91 8f 90 91 8e 8e 90 94 91 88 82 88 89 80 86 8c 8d 86 7d 7e 7e 77 7b 75 83 7d 7c 77 7b 73 76 79 76 7c 70 75 7c 7a 79 75 80 7d 82 86 89 88 87 8b 89 91 90 8a 90 7f 65 4e 1c 0b 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0b 06 05 10 0a 0d 13 3a 78 94 9a 94 95 8a 93 88 94 8e 8a 87 85 83 89 7c 7f 78 7c 78 79 76 79 77 74 78 78 6d 71 6f 66 6d 69 6b 70 64 65 6c 66 66 65 6b 6a 70 60 65 6d 63 5f 67 68 6e 6f 6a 72 66 72 6b 72 6e 68 6e 67 62 63 65 64 60 5c 57 5a 58 59 59 57 5f 5b 59 53 51 4f 4f 50 52 5a 52 5a 53 4f 59 5b 59 52 62 5d 67 75 65 5c 3c 24 14 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0b 19 22 36 3d 53 74 78 6c 62 58 4a 56 4c 51 55 59 54 58 59 51 53 56 55 58 59 58 51 5e 5a 5a 55 64 65 66 6a 6c 75 73 71 7d 84
 81 89 89 89 90 89 8d 98 8e 97 94 90 92 94 96 94 91 8e 92 90 90 89 86 88 87 83 87 83 7b 8d 83 86 80 72 77 75 71 75 75 78 76 75 73 77 79 76 6d 70 74 75 79 76 77 74 78 75 7d 80 83 86 84 8d 88 8d 92 8c 8d 8a 87 67 47 1a 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 07 0b 0f 11 39 75 89 95 8e 8f 86 96 89 92 8f 84 8d 84 85 7c 81 7c 76 7d 73 6f 76 79 70 72 6f 6e 67 6f 6e 68 62 69 6c 73 66 67 63 65 64 65 6b 65 6f 5f 60 62 5b 6a 61 62 66 6c 71 71 71 78 72 72 6a 6c 68 6e 60 67 68 6a 61 61 58 5e 54 5a 5e 5b 52 54 5b 61 55 53 52 54 59 58 56 56 5f 57 5f 52 53 55 57 67 69 76 65 5f 47 2c 19 0b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 15 0f 23 33 45 55 6e 75 69 60 52 56 53 51 4d 52 53 53 58 56 4e 55 55 53 59 5f 5c 50 58 59 59 60 64 67 5e 5d 6e 69 71 76 79 78 84 7f 91 83 8b 8c 94 8d 88 90 89 8c 94 8f 8d 90 8b 87 93 8d 8f 86 8a 81 81 84 87 7d 83 83 85 8a 7e 7d 6d 7b 77 73 6e 6f 73 73 6e 75 6b 74 74 7c 75 74 78 78 74 70 79 7d 7b 7d 7e 82 80 8a 85 82 8f 8a 85 8b 79 6a 44 1a 05 04 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 06 05 06 11 32 64 8e 8a 8d 90 87 93 8e 84 87 8b 86 8b 7e 80 77 79 7f 75 72 72 6d 75 6c 73 6d 6d 6b 6a 67 67 6a 66 5e 62 68 5f 65 64 5e 61 68 5f 5f 62 62 68 5e 62 6a 67 66 6a 70 71 7a 74 6e 72 6a 6e 6a 65 66 63 62 59 5d 5d 58 60 55 57 50 59 4f 54 5d 52 51 55 51 52 52 54 53 5a 55 50 56 59 57 51 58 5c 67 70 6b 5b 40 2a 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 17 1d 3f 52 61 6e 6f 6a 5c 53 4b 49 54 48 50 55 54 5a 5f 53 58 4d 54 57 55 59 5a 57 54 56 58 60 5f 63 6a 62 6e 6f 73 79 7d 7b 80 86 83 8c 95 90 93 8f 91 8e 89 92 8f 8d 90 85 8e 86 8d 80 8d 8b 8a 8e 87 79 7d 7e 83 7c 75 7e 7c 71 6a 67 6a 70 67 75 75 70 6c 6f 6f 74 76 7b 79 74 6d 73 75 76 7a 7a 76 7c 80 7d 7e 87 88 82 85 85 88 80 6c 4a 1f 07 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 03 00 06 05 2b 67 8d 95 8f 8b 86 8b 87 85 83 84 7e 81 85 82 6a 75 76 71 74 6e 6e 68 6e 64 67 6b 69 66 66 66 69 67 67 64 65 6b 65 62 61 64 69 66 65 64 60 5c 5d 65 62 62 63 60 6d 78 78 7a 76 73 68 66 62 6c 62 65 6b 64 59 53 51 5a 5c 60 58 55 54 59 58 55 54 4b 56 55 57 4f 59 57 55 58 55 5b 4e 58 58 58 60 6b 70 57 47 22 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 0a 0f 18 21 32 4a 60 6d 74 79 66 54 4b 54 4f 50 57 4f 5d 52 5a 59 5b 5d 5c 5d 58 5c 60 5e 5d 53 57 55 5f 64 6a 6e 75 73 75 76 79
 84 83 81 8b 80 88 93 8a 8d 8c 8c 8c 89 8b 87 8c 91 8a 8b 8b 87 88 90 87 86 7e 7c 7a 85 7b 7d 7c 7e 76 75 77 75 68 6a 66 72 6b 6f 69 6c 70 6c 71 7b 70 76 71 78 6c 7a 80 73 72 75 7d 82 87 7d 81 7d 87 84 7c 7f 69 4e 1e 03 02 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 07 09 07 09 0c 2a 65 88 90 8f 92 88 8b 84 8d 88 84 87 72 79 77 81 71 7a 72 77 73 6a 6e 71 6d 68 73 65 6e 70 6a 65 64 67 5f 65 5f 64 5d 65 66 67 64 61 67 68 69 68 5f 64 60 69 68 64 7a 79 7a 6d 6e 6e 6c 6b 69 64 6b 65 5a 5a 5d 5f 64 56 5c 5d 5a 66 57 5e 58 54 5c 5a 53 5c 54 54 5a 60 5e 60 51 52 5a 5d 55 58 66 68 52 49 30 19 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 11 14 2a 39 42 65 64 77 76 5e 51 53 53 4c 53 4f 4e 56 58 52 56 5b 51 5b 5e 60 5c 60 5e 61 5c 63 5a 63 5e 5b 68 6c 6d 72 72 7a 81 81 85 84 80 86 86 8c 89 8e 91 8a 83 8c 84 88 90 8a 8c 82 85 81 85 7c 86 80 78 80 72 78 7d 80 7c 75 6a 68 69 60 69 6b 6d 6d 67 68 6d 6a 6c 6d 72 6b 6e 6f 6e 74 72 78 73 76 7c 82 77 78 76 7c 7f 85 85 7d 80 65 52 1d 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 07 14 1e 66 81 8f 8c 94 88 8b 86 85 80 78 7d 7e 7a 7c 78 76 75 72 72 66 68 6c 65 67 5c 6c 65 69 6a 63 6b 6b 67 67 60 65 64 61 5b 5e 64 64 63 60 66 65 63 61 65 61 5a 61 68 78 6e 72 6c 69 62 62 69 65 62 60 60 5d 5e 5c 56 59 59 53 5b 57 5f 52 51 5d 4d 53 59 55 54 55 56 59 51 53 55 56 59 50 57 4f 52 60 63 54 4a 2e 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 0b 1a 2d 3e 4a 54 63 75 6b 5c 5c 52 54 4d 48 54 52 55 59 56 61 4f 59 5f 5d 60 61 5f 5e 59 56 5a 5b 62 5e 67 6b 6c 66 73 76 7a 7c 79 81 7f 7e 80 7b 89 8b 86 7e 87 83 83 85 84 88 84 83 84 82 84 80 87 87 85 73 7e 76 76 80 7e 75 70 6a 6e 67 68 60 64 6c 60 69 65 62 6c 69 6f 66 6a 69 6e 73 71 6e 7a 73 76 71 80 7e 7e 82 73 83 7e 75 84 71 63 48 22 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0a 0c 26 5f 85 94 8f 8e 83 85 7d 84 75 77 75 7f 79 79 71 76 76 75 73 68 69 6a 6b 69 67 65 62 60 65 61 63 5e 60 62 61 60 59 67 62 5d 62 53 62 5d 61 5e 65 65 64 5b 54 6b 69 6e 6b 71 71 67 69 5c 6a 67 60 62 5a 5b 55 57 56 51 50 5d 57 55 5a 56 5d 54 59 56 5c 53 5b 52 57 54 4e 54 4d 4d 4f 4c 51 55 54 58 59 54 46 38 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 14 23 28 36 52 5f 69 72 6b 5f 54 4c 5c 52 4d 56 4c 55 54 60 5e 5e 5e 5a 54 5c 5b 60 63 5d 67 5e 5d 5d 66 60 65 6b 69 70 6d 76
 77 76 7a 81 81 84 8a 83 81 86 87 86 86 82 83 85 7c 75 7e 85 7d 81 85 74 7f 79 7d 77 7a 72 79 7e 78 72 6e 65 60 63 61 6a 69 61 68 68 62 70 67 6b 6e 65 6a 70 65 6f 6c 6e 6b 78 79 77 78 77 75 75 72 7b 84 79 79 69 4a 1e 0d 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 01 09 05 1b 56 86 8d 97 8e 83 88 86 7f 7c 78 76 7b 76 7c 6e 73 6e 73 6c 6b 71 5f 69 69 66 69 61 61 5b 5e 64 69 66 60 5c 5f 63 5f 5f 5f 63 64 6b 5b 66 69 61 64 62 69 63 66 6e 72 6c 72 6d 67 69 60 67 60 5a 5e 65 61 58 56 53 5a 57 59 59 59 5c 55 56 5e 54 53 53 51 59 54 50 4a 50 46 59 4f 55 50 56 4f 4c 56 5e 51 48 32 1a 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 03 10 18 24 32 32 4e 65 60 72 74 65 56 4f 50 55 51 53 55 4d 53 57 56 53 58 5e 59 64 59 59 64 5e 5a 60 5e 63 6c 6c 6c 6d 6d 6a 6f 7d 7a 80 7e 79 81 85 86 7c 90 86 7a 82 86 81 84 87 79 7c 7f 81 7d 7f 80 7c 7f 78 72 76 75 76 79 78 77 73 67 6b 65 66 60 60 66 6d 62 69 69 67 62 66 69 62 69 66 6b 70 66 6e 72 6f 76 73 78 78 78 7e 7f 7a 76 82 71 62 4e 22 03 05 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 00 06 0b 1c 59 81 84 8a 84 83 87 78 7e 7c 7d 78 80 76 6d 6f 70 66 70 6a 6d 69 6b 62 5f 6b 64 67 64 60 64 61 5c 60 56 5c 55 58 5f 5d 65 64 5b 61 5e 68 61 57 5a 67 67 67 67 64 72 74 66 69 6b 66 66 60 60 5d 60 5a 5d 5e 51 5a 58 57 5b 5c 59 59 59 5c 56 57 5d 5d 4e 53 59 4f 5a 57 4c 58 58 50 51 47 55 4b 54 55 54 4e 36 1d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 10 17 1e 27 44 56 60 74 73 74 66 50 4a 48 52 50 58 4b 54 53 49 5a 5a 58 5d 53 64 5b 5e 5d 63 62 5f 64 64 5b 65 67 6c 68 69 71 6c 73 79 72 7c 83 7b 7b 7c 7c 80 7a 7e 7c 7d 7b 79 76 80 76 7d 7b 7e 81 7c 7d 75 75 74 6f 71 76 72 78 71 6f 70 58 62 64 5f 61 60 59 64 62 65 62 67 67 69 66 68 60 63 6b 70 79 70 71 6f 74 74 76 6f 76 78 77 7a 75 6d 50 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 06 05 18 51 7e 8a 8f 88 82 81 79 7d 7d 76 75 7b 73 75 71 6f 76 6a 61 69 6b 68 62 66 64 66 64 68 65 66 61 63 60 5d 60 5a 58 61 5d 5a 5c 5c 66 5a 65 64 5d 5c 62 64 64 6a 67 6b 6e 6a 6b 69 5c 5b 60 63 60 5c 5d 54 53 57 54 53 4e 55 55 54 59 4b 55 5b 59 52 51 50 5a 4d 55 5b 50 50 4f 52 46 51 4a 44 50 4c 50 50 43 3b 19 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 14 15 22 37 3b 4e 5e 68 76 74 63 57 5b 51 4f 49 5b 53 5e 51 53 59 4f 59 56 58 5a 5f 5e 5f 61 5a 5d 67 62 66 6d 6a 65 70 68 75 70
 73 77 73 74 7e 81 79 83 79 75 7d 7c 7b 79 78 78 71 79 7d 6f 77 7f 7b 77 73 78 78 75 79 77 74 74 71 78 71 69 60 5f 5c 5c 5d 61 5a 62 65 62 57 64 67 61 62 67 5e 66 6b 66 6d 62 74 73 73 70 72 72 77 71 75 89 74 64 51 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 06 06 05 03 00 0d 09 14 4b 76 81 86 87 84 7e 7d 81 7e 7b 74 76 6a 70 68 75 6b 6e 6a 66 67 69 63 64 5f 63 67 67 65 62 62 5f 67 5e 62 5c 56 5b 5b 5d 62 5c 66 5d 5c 6b 66 5f 5f 60 6a 64 78 75 66 66 64 6d 5e 63 64 5a 5a 5f 5c 54 56 5d 5b 54 52 50 56 5c 53 5f 53 5c 55 4f 54 4c 5a 55 59 51 4f 4f 56 48 4f 4c 53 4d 44 50 52 4b 47 32 16 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 13 14 1a 27 30 3b 4e 66 71 74 6d 62 4f 51 5d 54 57 54 4d 55 57 53 56 49 50 5d 55 5e 5c 59 62 5d 60 64 5e 60 6c 63 6e 69 64 69 71 71 70 76 74 78 7c 72 72 78 81 7b 78 7b 79 72 75 76 70 77 74 7c 73 74 77 70 76 6f 79 75 6d 77 72 72 77 6f 71 71 65 69 61 61 64 5b 56 60 58 63 62 5e 5b 5b 5f 68 62 65 6d 6b 67 6b 6c 6e 6e 70 6f 79 71 70 75 7b 6c 60 4b 2a 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 07 13 48 85 88 88 85 81 7f 79 84 77 76 73 7b 72 73 6c 6e 75 6b 6b 66 66 6b 5e 66 68 64 5d 66 62 59 65 5e 65 5f 59 5c 60 60 64 5e 64 5c 62 5e 60 64 5d 60 68 69 64 6b 70 6f 6e 6a 69 65 60 5f 65 63 5c 55 50 56 53 5b 54 56 52 5f 50 5a 56 51 57 58 53 50 50 4f 52 55 4b 51 4f 4c 55 44 47 47 46 4b 4a 4a 4e 52 47 2f 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 07 1b 1c 21 35 44 5e 64 6b 74 6e 62 58 53 50 58 51 55 55 4c 5d 55 4c 53 4e 5c 5e 5f 60 5d 64 5f 5b 5b 67 6f 5f 6b 69 6a 5e 65 76 74 71 76 76 72 73 75 78 6d 79 75 72 71 74 75 76 6f 71 70 77 74 71 75 69 72 74 78 76 74 69 63 6e 6a 72 71 6f 76 65 5f 66 5e 5b 5e 56 56 60 53 60 64 62 62 62 65 61 65 65 65 62 6a 6d 70 71 6e 6c 66 6c 6f 70 6c 64 5f 49 21 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 12 41 72 84 89 84 82 80 76 75 78 7c 77 71 76 72 67 6e 68 67 69 63 65 63 62 66 62 66 5b 60 5d 5c 5a 64 57 5b 5d 5b 57 56 59 57 57 64 56 5f 60 65 5d 64 6a 60 65 6c 68 6e 69 66 64 62 62 60 66 58 53 59 55 5a 5e 54 58 5a 54 5a 50 56 53 5b 54 53 4a 4d 50 52 53 59 54 49 4c 50 4a 4e 4f 4c 47 49 45 4a 52 4f 42 29 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 04 09 0a 0b 1b 1c 24 36 41 51 61 6a 71 69 61 59 51 55 51 46 4f 4e 54 58 52 54 55 55 58 56 5d 61 5f 65 5c 59 5f 61 66 5f 64 5d 6d 6b 6c 79 67
 6b 72 70 6d 7a 6d 78 75 75 81 6a 6f 7b 76 76 6c 6d 71 71 71 6d 68 71 68 6f 70 74 79 6e 74 6d 66 70 6f 75 73 6a 64 62 57 65 60 60 5d 62 5f 58 5b 5f 67 64 63 62 5c 5b 66 67 62 74 65 68 66 66 69 74 6e 69 65 70 5f 53 24 0a 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 0a 00 06 06 12 3d 75 7f 91 81 7e 7d 79 7b 82 6e 77 76 79 6d 6f 65 67 6d 69 70 67 67 6c 5d 5e 62 62 5a 63 61 5c 5c 5b 60 63 60 5f 5b 60 5f 58 5f 5a 5f 66 63 66 60 68 71 6e 69 6d 6b 69 66 68 5c 6b 61 5c 5b 51 55 53 5a 56 58 52 52 4f 4f 56 4f 56 51 52 5e 53 54 52 47 56 4e 55 4e 4f 53 4d 50 49 43 4a 49 46 48 4e 4b 40 23 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 09 07 09 07 10 1e 33 3a 41 56 61 6d 6d 6a 57 55 50 54 4f 53 55 54 4a 55 4f 5a 5b 52 5a 59 59 60 5a 54 5c 62 5c 67 64 6b 62 63 6a 65 64 6d 6a 6f 72 6f 6f 6b 71 6a 70 73 71 75 71 71 70 6e 6b 70 73 75 6a 69 6a 63 6b 6a 6b 71 6f 6f 6a 6a 69 6d 70 75 73 69 66 65 60 61 59 64 5f 57 5e 5e 5b 62 54 64 5c 6d 63 61 62 67 65 65 64 69 6a 69 6d 6c 72 6b 68 61 5d 48 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 15 39 78 86 86 8a 85 7d 75 7c 7d 74 73 77 69 76 67 6c 6d 64 6e 6f 65 68 61 6a 62 64 62 5f 68 62 5e 60 60 63 5c 5d 64 5b 64 5f 5a 60 63 5c 61 67 5c 5b 6d 6b 6c 70 6a 6a 6b 66 61 6d 6b 67 65 5e 5b 50 57 58 53 5b 54 4d 55 5f 4e 54 51 58 4a 4f 4c 53 55 4f 50 51 5d 55 4c 4b 4b 4a 4c 47 49 3e 44 49 45 47 3d 2f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 08 0d 0e 25 25 3a 4e 54 64 75 68 5f 4d 4d 51 4b 45 53 51 55 58 55 53 51 5c 53 4c 5a 58 57 60 5c 5b 5a 5d 5d 5e 61 63 66 6c 6a 5f 66 6d 6a 69 6a 6d 6a 70 6a 74 6b 6d 74 70 6b 6e 70 6c 6f 6a 66 6b 66 6e 66 5e 67 64 64 66 63 69 6b 6d 69 64 6b 6c 6f 68 5d 5b 62 54 5a 5c 53 5e 5a 60 63 5e 5a 60 5c 5c 5f 60 61 60 65 62 63 60 61 60 61 66 66 64 60 5e 48 21 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 30 79 7b 8b 7d 77 76 6e 7a 77 75 75 73 73 65 69 67 69 6e 67 61 63 5e 64 65 61 63 5d 5c 5e 5d 5c 5a 5f 60 5d 54 61 62 5c 5f 64 58 60 5c 56 65 5f 69 6d 70 70 6d 6b 6c 60 6e 60 63 68 64 66 5c 50 56 4f 59 51 52 57 58 53 54 4e 4c 4f 50 51 4d 4c 50 4d 48 49 4e 50 52 48 4c 48 47 42 46 47 42 41 44 43 3e 31 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0d 05 0a 17 1c 2e 35 41 52 64 6f 68 5a 51 52 4c 5a 52 52 59 50 53 5f 52 55 53 51 4f 56 53 63 5f 58 5c 5d 60 5b 64 5c 5f 5a 63 5f 6c 6b 65
 67 6d 6d 6b 72 64 6f 64 68 70 69 6a 6e 6a 65 6f 6b 69 6f 64 71 69 64 62 65 65 63 69 62 6b 6f 70 69 68 6b 70 71 6a 67 64 5e 5d 5a 5a 5b 57 57 56 5d 65 60 5c 59 62 58 5b 5a 5f 69 63 5e 64 5b 57 58 61 60 5d 6b 53 4d 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 0f 30 6f 84 81 77 75 7c 73 81 76 75 75 70 70 73 6a 60 68 5f 6a 6c 65 69 66 63 5e 64 65 5d 65 64 5b 62 64 59 62 61 65 5c 60 5b 5f 5b 5f 5c 60 64 64 61 6a 70 71 6f 65 6b 6a 68 61 6d 6e 79 6e 61 56 57 51 4b 53 55 53 53 4c 56 50 50 50 50 4d 50 4e 4f 4c 4f 4f 49 53 50 4c 4b 49 41 45 3e 45 40 43 46 3f 3e 30 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0d 10 16 22 39 3b 48 59 6c 67 70 5a 54 53 56 4f 4f 49 52 50 53 5c 53 55 5a 57 4e 4f 5b 5b 5a 55 5a 53 58 67 5e 5a 69 65 69 66 69 6c 6d 63 65 6c 63 6d 6b 65 68 65 6a 6e 67 6c 66 6b 69 6f 68 68 65 5c 66 65 63 62 62 5f 68 64 5f 62 66 62 5c 6a 6e 6b 67 6a 65 63 61 58 5e 5a 62 55 59 60 5e 64 5c 5a 5f 59 5f 66 5a 64 61 62 5f 5c 5c 69 60 56 60 5b 53 3e 27 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 0d 11 2d 68 7d 88 83 7a 72 73 7a 76 71 75 7a 7a 76 6d 66 69 6e 67 67 64 63 64 68 6e 60 64 66 64 67 59 65 61 64 67 62 69 65 60 5f 62 64 62 5f 63 68 63 6b 6f 78 6e 6c 73 64 65 60 69 6e 7b 81 74 68 60 58 5c 53 4f 55 57 50 4f 52 4d 51 54 4f 4e 52 50 52 4f 50 54 51 51 54 4e 4c 47 42 44 44 45 4a 3c 42 40 32 24 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 05 06 0c 14 10 2b 27 38 4e 54 67 71 72 68 53 52 53 4a 53 4d 59 52 58 5a 57 5b 5b 54 4f 55 54 57 5b 59 53 54 55 5b 63 5f 62 65 64 5e 63 69 63 5f 6f 64 5f 66 6e 63 6a 6d 6c 62 60 65 67 63 65 69 5f 5d 63 62 60 60 64 61 5e 60 62 60 63 64 5f 61 67 62 68 6b 67 68 68 5e 55 51 57 5c 52 5f 5a 61 5d 59 4c 55 5e 55 5a 5f 57 5d 5d 54 5e 62 64 56 5a 5e 55 66 51 3f 23 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0f 0c 23 66 7f 7d 7f 79 7e 78 7d 79 74 74 74 70 6e 6c 71 6f 6a 73 6e 63 64 60 63 68 64 68 6a 65 62 69 66 69 65 60 6a 61 65 64 5e 65 5f 5e 58 5d 6a 65 6c 74 64 6a 6a 65 69 58 5f 69 77 75 86 6b 63 51 4e 57 53 4e 4f 53 53 4f 4f 44 4d 4a 50 4c 4d 50 4e 52 51 4d 49 4d 4f 49 48 40 44 43 45 44 49 3a 38 38 2c 1f 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 08 10 1f 22 33 46 4f 5c 6a 65 6f 66 5b 4e 50 53 50 51 52 54 56 59 57 55 4e 54 5b 5c 56 58 54 56 54 5b 59 5d 5d 5e 60 64 62 61 63 5b 64
 61 5f 65 63 61 64 61 65 66 64 65 5f 64 69 66 6a 66 5a 60 68 5d 63 61 53 64 56 62 57 5f 5f 5d 5e 64 62 63 64 5b 60 6f 64 5b 62 5a 64 58 5f 57 4d 5c 58 5b 5d 5d 5f 5e 58 56 59 58 5b 5f 56 61 60 5f 5e 5c 59 5b 53 48 22 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 23 66 78 86 7c 72 76 76 7d 70 6e 6d 6f 78 6f 72 67 72 72 68 61 69 70 64 69 59 68 64 69 66 67 71 60 64 65 68 6e 6c 70 6a 66 60 6a 5e 62 64 64 68 63 6b 6d 6c 6f 5d 65 5d 67 6d 7e 7f 71 6e 5e 52 53 56 4f 52 4f 4b 50 46 51 4e 4e 4f 4f 54 49 54 41 47 53 49 42 4e 44 3a 46 4a 3b 44 44 48 45 3b 45 37 26 13 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 0d 0e 1c 21 2c 47 4a 65 6f 71 6e 64 5d 4c 53 49 4d 51 4b 59 55 51 55 55 59 4e 56 5c 56 56 56 56 58 54 5b 5d 5d 5b 5c 62 5d 5b 60 62 60 61 64 64 5e 67 68 6e 63 66 64 66 65 62 66 5a 5e 60 6b 68 63 5a 5e 5d 68 5c 60 63 5a 5b 63 5e 63 5c 62 67 64 63 66 6a 68 64 5d 65 5d 60 60 53 56 5c 53 57 57 5c 60 55 56 5b 5f 5c 5a 5c 58 59 5c 57 5a 5a 55 54 50 45 20 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 2a 58 73 7d 7c 76 75 72 7b 75 75 75 70 71 76 6a 6e 6e 6b 6b 65 66 65 62 64 62 6e 65 67 6b 64 6b 6f 70 66 68 6c 67 71 70 70 6c 6c 6b 65 6a 66 66 6f 70 65 6e 61 6b 5e 5f 69 69 75 71 6d 66 5e 57 4f 57 53 57 5a 54 53 43 51 4d 50 48 4e 47 49 48 48 4a 4c 4b 4d 48 4b 4a 4c 50 45 4a 44 4b 46 40 39 28 20 17 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0f 13 17 2b 35 44 4f 5b 69 6e 7a 6b 5c 47 52 4c 55 47 51 50 54 59 57 55 52 52 54 59 58 5b 56 57 5b 59 54 5b 58 5a 61 5a 5f 5e 56 5a 5b 5b 5a 62 5d 5d 65 5b 63 65 6a 66 60 60 61 65 60 62 5e 62 5e 58 5f 5f 64 59 51 5b 56 57 52 5b 60 63 62 5d 61 5e 6b 5f 70 66 5d 5b 5c 5a 5c 5c 5d 5e 5a 5b 53 54 54 55 5a 56 54 5d 56 59 61 59 55 57 5a 5c 56 54 53 38 20 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 04 06 05 03 16 5e 78 7c 75 76 75 70 72 72 73 72 71 75 70 6f 6a 69 6d 6b 67 67 6c 6a 6a 62 6e 62 6e 6d 5e 6d 69 6e 71 6f 6c 6e 75 74 74 75 64 6f 69 70 6c 6e 6f 6f 6d 6e 60 5e 53 59 64 67 6d 68 64 5e 53 4e 4e 4f 55 4e 4b 4e 49 4d 46 52 4c 4f 4d 4d 54 47 4f 4f 47 47 4a 49 45 49 46 49 43 45 44 45 47 43 37 29 1b 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 06 0d 16 1d 2f 30 41 50 5e 67 69 7b 6a 5e 51 4a 50 49 4d 55 44 4b 51 50 4e 57 58 56 4e 57 52 4d 60 53 58 51 55 5a 59 5f 59 5e 62 5a 57 5a
 56 64 5e 5d 54 60 5c 56 61 5c 5d 64 62 55 65 62 5c 62 60 67 5c 5e 5f 59 5a 60 55 51 5b 58 57 59 5d 58 61 62 5c 64 6b 66 65 5d 5f 64 55 60 59 5e 54 4e 5a 5a 4f 57 5b 50 57 5b 5e 5d 57 5d 58 56 5b 54 57 58 4c 51 42 22 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 05 1a 57 75 7f 7b 79 75 77 6a 6d 73 72 78 75 6f 71 77 6d 70 66 6f 63 6b 5f 6e 64 68 62 6b 6e 67 71 6c 6a 72 63 6e 75 74 7e 74 83 7a 73 70 76 70 71 71 74 70 69 63 57 5d 5b 60 63 70 62 54 53 51 50 53 4c 4b 50 50 51 4a 48 4c 4c 48 52 54 49 48 45 48 48 4a 45 4e 44 41 46 44 43 47 43 45 3b 44 36 36 1e 0d 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 20 2b 35 44 4f 60 72 71 7d 72 62 55 55 46 47 4c 48 4d 51 50 4f 58 4d 5b 50 4e 4e 52 5b 59 54 58 58 4e 5e 56 52 5e 5b 58 58 5b 62 57 62 5a 58 5d 5e 65 60 5a 5b 5e 5a 5e 69 5f 61 58 5e 5f 5b 5a 59 5c 54 5c 5c 54 5c 59 59 5b 5f 5d 63 59 5a 58 61 6c 71 6d 64 65 69 54 59 5a 4f 57 58 59 50 51 4f 53 58 5c 54 5e 53 62 58 5c 5a 5a 5e 5c 5d 58 52 3d 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 16 4b 78 7d 7c 76 74 75 75 75 6b 72 6e 70 75 6b 6a 67 69 6d 6a 68 72 65 70 6a 69 6d 6c 6b 6a 62 6c 69 6b 62 6a 72 72 77 85 81 8a 89 7a 77 79 75 78 79 6c 67 69 61 60 64 62 5f 5f 5f 60 54 56 4b 4c 4e 54 55 4f 52 4a 49 4c 4f 4f 4d 57 44 52 4b 47 4f 45 4c 4a 43 4b 49 4f 48 4d 4e 46 44 40 39 2b 18 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0c 19 1b 2d 4d 53 66 71 6f 7b 73 6b 59 52 4b 52 4f 4f 53 52 55 5c 5a 4d 52 52 4f 5b 58 58 56 53 55 57 52 59 5e 50 52 54 5e 58 5e 55 56 5a 5b 60 5b 56 5d 62 5c 60 5b 59 61 5b 5e 5b 59 60 5d 5b 59 56 60 4f 58 58 54 59 58 51 5e 5f 59 60 60 5f 58 63 6f 6d 66 5d 62 64 68 60 5c 59 53 53 53 5f 58 5b 5a 5e 58 52 61 54 53 5e 64 60 5c 56 5a 51 51 53 42 20 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 19 55 78 79 82 75 74 6e 71 78 72 73 6c 72 6c 74 74 73 6f 65 69 68 69 6c 64 66 69 6a 6e 6a 64 69 63 63 64 71 6a 71 71 75 79 83 7b 83 7a 74 81 69 78 74 6f 70 66 63 62 5e 5c 64 64 60 5e 5b 51 4c 50 57 52 4d 4e 4f 46 45 54 4b 47 4b 52 4c 47 46 4b 4e 41 4a 49 45 4a 45 49 46 48 4e 43 46 3e 29 29 12 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 08 0e 19 1c 34 38 49 5f 6c 69 73 78 6d 54 48 4e 44 44 50 4a 4b 48 56 51 4d 54 4f 52 55 51 58 4f 52 53 4c 54 53 57 5a 55 56 5b 59 59 57
 5d 57 55 55 55 5a 59 5e 56 5e 54 64 5a 58 57 5d 54 54 59 5a 57 55 5a 5a 61 5a 4f 55 57 59 5a 5b 5a 54 51 64 62 63 6b 6c 72 55 6c 5f 55 5d 54 5b 50 4e 54 53 4e 56 52 53 5c 54 59 57 57 59 4f 59 5c 5b 53 55 4c 4f 39 1d 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 49 74 7c 76 71 70 6e 75 72 74 73 71 70 6e 6b 75 6d 6c 6e 72 65 6d 6d 6d 61 62 6b 6b 67 65 66 6d 71 6c 65 61 6a 6c 6c 75 7a 7f 78 6e 70 71 6c 70 77 73 6b 6b 6b 64 5b 61 62 5d 5f 54 50 58 47 46 4f 50 55 4c 42 4a 44 4d 46 4c 48 4f 44 53 3c 49 43 45 48 4d 43 4a 43 47 4a 47 44 3e 44 43 24 18 08 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 04 18 22 32 36 4c 5b 6a 6e 7f 76 6c 5a 54 45 4a 44 4f 47 4e 49 50 54 54 4a 52 55 55 58 51 4e 4a 50 50 53 5a 54 54 51 55 59 5b 5a 5a 55 5d 4e 5a 5f 53 61 5a 5e 5a 56 5d 59 59 60 5a 51 59 57 54 53 51 53 57 54 56 5e 58 58 56 4f 56 5a 5a 61 62 62 69 70 64 6a 67 62 60 58 62 62 5b 58 58 4d 5c 59 4c 55 58 51 52 55 56 4d 59 59 61 55 54 58 55 52 54 42 21 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 10 50 77 83 80 79 76 75 78 76 6c 69 6e 6e 73 72 6e 6e 6d 6b 65 65 69 6c 6f 6a 6f 62 6c 65 71 6a 66 65 6c 6d 6b 69 61 68 76 72 72 75 6e 70 6d 64 69 6d 75 75 6e 63 65 65 64 62 62 5b 53 53 4f 57 50 57 51 50 4d 53 54 4d 49 50 4d 48 46 53 4b 3f 44 47 4b 4e 46 4a 49 41 43 47 41 43 40 43 36 2b 1a 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 13 20 2e 2a 42 59 62 67 78 70 6d 52 4f 4c 48 4c 4b 49 46 4e 45 4b 4d 4a 50 4e 50 53 53 53 51 4a 53 55 56 5b 59 54 54 57 50 54 54 57 59 5c 54 51 58 58 52 52 5d 57 57 5c 61 58 54 56 58 59 57 55 53 55 54 51 54 56 50 4c 52 5a 59 5f 59 5d 5f 66 70 73 6e 69 63 65 5f 59 5c 55 53 56 52 53 4f 4e 54 56 58 52 55 55 54 51 5d 59 56 53 55 56 4d 4d 4f 3b 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 07 0f 4e 73 7c 87 75 75 6f 6f 72 78 74 75 70 74 68 69 71 70 66 6f 6b 6f 69 6d 6b 6d 65 6a 64 6e 70 6a 65 6e 73 6f 6f 6b 67 64 6b 68 69 64 68 62 6f 6b 6d 77 72 6f 69 5a 60 60 5f 5a 55 52 51 50 50 58 57 48 48 51 51 5a 4c 51 47 48 43 50 50 54 4e 41 45 41 47 46 43 4d 48 4d 49 45 4d 3e 3d 36 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 03 11 12 29 29 40 57 5e 6b 71 7d 65 5a 51 42 3e 3b 43 4a 49 4d 49 53 44 4f 44 4e 4a 4f 57 4f 52 4f 50 55 54 52 55 5d 5f 5a 56 5e 55
 54 51 51 51 54 4e 55 58 56 58 57 54 52 5a 51 58 5c 55 4e 56 50 50 55 54 5a 52 53 49 4f 53 55 52 54 52 55 63 69 72 65 66 65 5e 5c 5d 56 58 4e 54 55 53 52 50 4b 54 4f 51 4d 4a 56 54 5c 51 59 57 50 53 5d 54 4a 50 42 26 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 43 79 7e 7b 7c 78 74 74 76 71 73 73 76 73 74 67 6b 69 6f 72 72 70 73 66 6d 71 62 71 6a 70 6e 6b 72 74 6e 70 71 72 65 66 62 63 64 5e 65 60 65 66 72 75 73 6f 65 5f 5e 57 4e 57 55 51 5a 51 4f 4f 4b 49 4e 50 46 49 46 46 3e 46 4d 46 44 44 41 44 4d 40 44 44 4c 3d 4d 50 44 47 43 3f 3b 27 12 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 12 1a 25 2b 38 4b 55 66 72 79 72 5a 4b 46 3f 46 44 46 49 47 50 47 4a 4b 4f 58 4e 52 53 4e 54 4f 4f 59 54 55 57 57 5b 5b 5b 55 59 5b 5a 5b 53 59 54 58 5f 52 5b 56 57 5b 5c 4c 54 59 51 5e 56 4c 4f 50 50 56 5b 4c 59 51 51 58 59 5d 64 65 69 64 6b 66 63 60 5f 5c 5c 53 53 54 55 58 53 52 55 4f 51 4b 48 52 50 47 55 52 52 55 50 54 4c 58 5f 52 4e 47 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 3c 6c 7d 78 77 72 6d 77 75 71 76 7a 76 7b 70 74 76 6a 73 67 6a 6a 6e 70 6d 70 6c 6c 6b 6d 69 6e 66 6b 6a 69 76 73 70 71 6a 6e 65 66 69 5d 5e 64 69 6c 78 6d 68 5c 58 54 50 50 51 50 56 48 49 4c 4e 48 52 4f 4e 4d 47 4b 49 4b 53 4b 45 46 48 41 4a 46 4d 4b 4a 42 46 46 49 50 44 43 36 2a 0d 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0b 1a 1a 29 2b 44 52 65 6f 6b 64 5b 48 3f 3f 44 4a 4b 4d 51 4e 4c 43 52 47 54 44 4d 54 57 4b 4c 51 4b 55 57 58 56 54 53 56 53 5b 55 5a 57 54 57 51 57 51 5e 57 4d 54 53 59 4f 59 57 59 54 59 53 58 52 51 49 4e 55 55 57 52 58 5d 56 5a 67 69 6f 6f 63 62 66 5c 61 58 56 53 57 59 4f 51 48 4f 54 56 52 50 57 58 60 55 53 58 51 53 55 4f 53 54 4d 42 40 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 02 3a 6f 79 81 74 7c 6f 79 7a 77 6e 75 79 70 70 70 76 75 68 70 71 71 6c 74 6e 72 6d 70 6d 71 6a 6e 77 6c 6d 6f 6f 65 6b 68 67 67 66 61 5f 6f 6d 66 6e 70 6a 67 67 52 52 56 53 55 54 55 51 49 48 4e 52 4b 4b 4f 4d 43 49 49 4a 45 43 4f 4b 53 4b 4f 49 4d 4d 4a 47 49 47 4a 4c 4b 46 3d 28 22 18 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 14 1c 22 2f 31 4e 54 5f 6d 64 55 49 45 3e 3e 45 47 49 49 45 4e 3c 3a 43 44 4c 50 43 50 4b 4c 4a 4c 54 55 54 56 60 4c 4b 51 56
 4f 5a 51 53 56 5b 54 58 56 56 4c 5a 50 48 56 55 53 54 54 55 54 49 52 4e 52 4a 4b 4e 4b 53 5b 59 5a 5c 60 6d 62 63 5f 5b 67 51 56 57 59 58 51 55 54 4c 4e 4e 4f 54 53 4e 54 49 52 52 4d 51 55 50 52 50 56 52 50 45 43 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 2f 65 76 75 7c 74 6a 70 72 70 77 76 6a 75 76 6d 70 6a 75 71 6e 73 73 6a 6d 6f 66 73 6c 71 6f 6a 6e 70 6b 70 67 67 65 64 5c 60 59 60 63 61 65 66 6e 70 64 60 55 54 44 50 4c 4a 4b 48 49 56 47 4a 53 45 4c 4b 4b 47 4d 47 51 47 46 50 4a 45 4b 43 44 47 4e 46 4b 43 4a 4c 47 47 40 2d 2e 17 10 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 1b 1c 27 2f 36 50 54 63 60 4f 42 3b 3f 48 3d 4a 45 48 40 45 48 47 49 45 4e 53 4c 45 4a 59 4f 4e 57 4d 58 57 5a 58 58 5b 57 58 4f 51 54 4a 53 4d 53 57 55 53 53 52 56 48 53 54 49 53 50 4d 56 49 51 4d 54 4f 51 4e 55 58 58 57 5f 61 68 5b 58 5d 5d 58 5e 61 54 4e 51 4a 4e 55 4b 51 52 51 4c 4d 4c 52 56 58 54 4e 52 4a 56 54 58 56 46 4b 49 3e 21 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 2f 63 79 74 6f 7a 6d 79 77 6f 76 71 72 75 6d 6f 73 71 77 72 6d 70 6b 74 67 6e 72 75 6a 74 69 6f 6c 67 61 6c 64 65 63 65 5e 60 5e 55 5a 5a 5b 5e 62 5c 5e 5a 51 4b 52 51 4d 51 4a 45 4f 4a 49 4d 4d 49 50 4d 47 41 4a 41 45 51 45 4c 4a 45 51 48 45 44 46 47 43 44 3f 43 4c 45 41 27 1e 17 09 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0c 14 1a 1f 28 35 42 4c 5b 54 47 50 44 43 45 46 42 4b 47 4b 44 4a 4c 4b 49 47 46 53 53 48 50 45 4c 55 54 55 5a 5c 52 55 55 56 58 5f 5b 53 52 50 58 56 52 5d 5a 54 51 53 4f 4a 4d 56 50 57 4d 53 58 51 5a 4b 4c 50 59 52 58 5f 5c 67 5e 66 61 5e 55 60 59 60 56 59 56 50 52 54 48 56 55 48 4c 4e 50 51 4d 51 58 59 52 55 53 52 52 51 51 53 4e 4f 40 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0e 20 5f 79 73 6f 75 6b 74 78 7b 6e 75 79 77 74 76 7e 75 77 7c 76 73 77 73 70 74 72 69 79 75 6d 70 73 70 66 67 65 62 60 5c 5b 5c 5c 5e 5e 66 60 5c 64 59 5a 56 50 4b 45 4f 4e 4d 51 4b 49 4f 47 4d 50 50 4f 4c 4e 4a 4f 4f 59 58 4a 4e 42 52 4d 4c 4e 53 41 4b 4c 49 51 44 4b 43 33 27 16 10 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 13 18 27 27 31 46 4a 42 41 3f 47 44 41 49 3f 41 49 46 3c 4b 46 4a 48 4a 4c 4c 4a 4c 4a 4a 4e 47 4b 4f 55 5d 4e 4f 4c 54
 5c 5f 55 54 56 4e 54 56 52 54 4a 55 56 4f 51 52 46 53 4a 54 48 51 50 4c 4e 45 4d 53 48 4f 58 61 5a 5b 57 54 5c 5d 4c 5b 57 5b 5c 54 53 50 4b 3f 55 4a 4e 54 4f 4f 50 53 53 51 44 46 4a 4b 4f 54 55 4e 4d 48 4a 4d 3c 20 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 19 64 6d 80 7a 73 73 78 71 6b 74 70 73 76 73 6d 74 69 73 74 77 78 76 71 6d 75 6c 74 72 74 73 6f 6c 69 69 60 65 5f 64 62 59 56 5b 55 5f 5c 58 59 59 56 51 4f 4a 49 4b 42 4f 4d 4d 4a 4a 4e 4c 45 42 47 54 4e 52 46 49 45 4a 4f 4e 4d 4d 4b 45 46 4f 42 45 4a 4e 4d 4e 45 47 41 39 1f 15 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 05 12 1a 23 2d 31 3a 3f 45 44 43 47 3d 48 45 43 44 3a 45 40 46 4a 44 4e 4b 4d 4a 55 49 4e 4f 4b 46 52 49 54 55 59 5e 54 50 58 4f 54 55 55 52 52 56 57 50 4c 4c 4c 51 51 52 4c 52 4e 4e 46 49 45 4c 44 4a 4c 4f 53 56 57 60 61 5b 63 59 54 52 5d 5a 5c 59 47 4c 4d 47 50 4b 45 47 54 4d 50 4b 4e 4a 55 51 4c 4d 50 56 4a 4c 4e 53 47 45 40 3f 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 22 55 75 79 70 6f 6b 69 70 75 6e 6d 6e 6e 75 6d 72 72 73 72 77 74 7a 72 74 74 6f 6f 79 6e 6e 71 6e 6e 67 64 6c 64 5d 5a 5d 5b 5b 5a 64 56 53 53 57 52 52 4c 4e 53 4d 50 4d 4b 49 46 4e 45 48 4c 52 43 43 44 4d 45 45 4e 4a 47 4b 4a 4a 50 49 4e 48 46 4e 40 48 45 48 46 41 3a 26 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 1d 28 30 34 3c 3c 41 43 3b 46 40 45 3c 46 3f 4b 3c 44 41 41 48 44 46 4f 4a 45 47 4b 4f 50 5c 53 51 53 4a 56 5d 53 58 5c 59 53 4e 4d 4b 52 4a 5a 4d 51 57 4f 55 4b 4c 51 56 52 4c 4a 49 50 4a 4a 54 4d 57 5b 51 5f 60 58 5a 5b 4f 55 59 5a 5b 50 50 4f 51 46 4d 4d 4f 4f 4e 45 4d 56 58 4c 55 55 4f 54 53 56 4e 53 45 4d 4e 46 42 4f 3b 1a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 5e 75 70 78 69 64 6d 70 71 73 76 6a 6a 6e 75 76 75 79 77 72 77 70 72 6f 78 75 73 6b 72 6d 6a 75 64 64 62 5e 5a 5a 5f 5b 51 5a 5b 61 57 55 59 4d 5a 54 54 4e 4b 45 4b 4d 4f 54 4a 48 47 45 47 4d 47 4a 52 50 53 44 49 4b 49 4e 57 4f 51 46 4a 43 4c 4a 4e 4b 47 47 40 47 39 29 12 13 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 13 14 1e 27 2e 40 3d 3f 45 40 42 41 46 3b 46 42 48 45 3a 3d 46 40 4c 4a 4f 50 4b 4c 4f 51 50 53 4c 4b 4c 4d 51 54 56
 52 5b 55 52 57 55 52 50 56 49 50 4a 51 54 4a 4a 56 4d 4c 4a 4e 4d 48 4f 51 4a 44 46 52 54 56 64 65 60 53 54 43 52 56 54 5c 4f 54 4e 53 46 45 48 4e 50 4a 53 4a 4b 50 44 53 50 49 46 4a 58 4e 4b 4d 53 49 4b 41 44 3f 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 1a 5a 6a 73 75 6e 61 70 75 64 77 6d 78 71 6e 70 6a 70 6d 6a 6f 69 6b 6b 6d 70 67 70 6a 73 6e 6d 68 61 62 61 5d 5e 58 58 55 56 59 5d 5b 5a 50 4b 50 54 4d 50 4a 4a 4f 4b 4e 49 4b 47 46 50 47 4d 4d 52 4a 4f 4d 42 41 45 49 44 49 51 4b 4b 43 49 44 46 49 4a 47 45 3f 4a 3b 37 1f 14 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 08 11 22 22 2c 36 3d 39 44 3e 45 3a 3c 45 47 45 4d 48 42 46 47 47 45 47 4c 4c 4e 49 54 4f 48 52 48 4e 54 54 59 56 4a 51 56 50 48 52 51 4e 49 4b 4f 53 45 4a 49 44 4f 4d 4d 49 48 4c 48 55 42 4c 47 4b 4d 53 58 5d 67 5f 5a 5a 4c 55 54 56 53 5b 52 58 54 45 45 47 4b 4a 4e 42 3d 47 45 4a 4d 4b 50 4b 4b 43 50 50 52 4c 48 44 42 40 42 38 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 16 53 6d 6b 73 6a 67 70 67 6c 65 70 68 6f 6c 70 70 6b 71 76 71 75 6f 73 6a 6c 69 67 6c 69 62 67 6b 69 65 62 5b 57 4e 5d 52 5a 52 53 5a 5a 52 4c 4f 4f 4a 43 43 46 4b 4f 4b 50 48 4b 42 49 48 4f 43 44 4b 49 44 49 44 4d 51 50 53 4c 4d 47 4a 4c 4d 47 49 4a 45 49 46 3b 3b 27 16 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 14 18 27 27 2f 3e 41 41 3d 44 46 3c 39 3f 46 45 41 40 3e 42 49 47 48 4e 4c 49 46 42 50 4d 4e 4f 4a 4d 53 57 52 52 59 54 51 53 52 55 4c 55 4e 4f 4a 4c 4d 4c 47 45 50 4a 4f 47 48 4f 48 50 4a 4c 4c 47 4f 62 5d 60 5c 4e 4b 54 51 53 57 49 54 5c 5a 54 4a 4f 42 49 48 41 49 50 45 46 4f 45 4a 46 50 4d 45 4a 47 47 46 4d 4a 4e 47 40 3f 21 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 4d 6e 6d 77 70 6e 6c 69 6c 65 70 6b 6e 6f 68 6c 6f 6d 71 69 66 71 69 66 6f 67 69 63 72 61 6f 6d 64 67 61 5e 5d 51 56 51 59 53 56 54 4d 4c 50 52 4d 47 4d 4c 52 50 4d 48 47 48 44 45 4b 45 50 49 4b 4a 4f 47 48 4c 49 4c 45 50 4f 45 4f 49 4c 4a 4b 4e 46 4a 49 3b 46 2c 27 19 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 12 1d 30 35 34 36 3f 41 49 44 3e 47 3e 46 4f 40 44 47 42 42 48 4b 4a 49 40 4b 47 4d 54 54 4f 54 50 4f 4d 4f 54
 51 53 56 53 51 50 52 54 4b 4e 4b 52 52 4c 4b 41 4f 47 44 4e 45 47 3f 46 45 4b 4a 57 54 5b 5c 5a 5b 51 48 4c 4c 4a 48 50 5c 53 56 59 51 41 4b 4b 48 4a 47 4f 44 4b 53 4a 44 4e 4e 4e 4b 4e 48 4b 48 53 4d 41 47 42 46 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 19 49 69 70 6f 69 60 65 69 6c 69 6b 65 68 69 64 6f 6e 6f 70 6e 6f 69 66 6a 6b 5e 67 73 64 68 60 5d 64 56 58 5f 54 5e 5f 5b 5b 5a 56 56 53 4c 43 52 4e 48 4d 45 50 4f 4d 41 4d 4b 46 4e 46 46 46 45 46 4a 4e 47 4c 4b 50 4a 4b 4c 4f 4a 48 54 47 42 44 4c 4f 48 4a 39 37 2e 22 1b 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0d 0f 20 2f 35 3f 47 44 41 3c 42 3a 43 3d 42 3c 48 3e 47 4e 49 48 49 42 40 46 43 4f 4e 4c 3e 42 4f 53 4e 4d 58 54 56 51 4c 50 54 4b 47 4b 4c 4d 42 4e 47 55 49 43 43 51 45 4a 49 45 4d 4f 50 47 56 50 59 5d 55 4f 4d 4a 4b 4c 50 52 4d 59 55 5a 50 47 4e 4d 44 42 4f 4d 43 48 4a 4f 4a 44 44 4a 4d 45 4a 47 46 49 42 47 47 4a 3f 3f 1f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 48 5f 71 66 62 60 63 6b 67 6c 68 66 67 6e 64 71 6d 63 6e 6d 6a 69 67 66 68 6c 62 66 60 62 60 65 63 5d 5f 5c 50 54 55 53 53 4f 50 4d 4b 4c 4f 47 4b 45 45 49 4c 4d 43 3e 48 48 4d 49 44 45 4a 46 4b 4c 4e 43 47 4a 4f 4b 49 44 4b 4c 4b 4b 45 40 45 4b 42 42 42 37 39 2e 17 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 15 25 2c 2b 48 45 45 45 3d 3d 3e 45 42 3e 43 42 44 41 44 45 43 46 48 49 41 45 49 4a 4f 4c 52 54 46 51 4e 53 5e 53 52 50 4e 52 51 4c 52 50 49 4f 3e 55 4a 47 4b 47 43 4c 44 3f 4b 44 49 4b 58 5c 5e 5f 59 54 4e 4e 4d 4a 47 45 4b 54 5c 5d 56 4e 4b 4b 4b 41 49 40 47 47 48 3f 44 41 3d 4b 4a 47 49 4b 49 46 45 48 48 41 40 42 3e 21 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 14 47 6b 68 70 65 63 6b 64 64 6c 6a 6a 69 6d 68 6d 66 72 68 65 6a 6e 69 69 6a 67 6c 66 6b 6e 61 5f 59 58 52 50 4f 57 51 53 55 57 54 55 4a 53 56 4e 4a 47 45 42 4b 4a 3f 4b 48 46 42 44 49 44 46 48 49 4b 4e 55 48 4a 4c 46 44 48 5a 45 48 47 50 4c 46 4a 48 48 3c 35 2c 23 10 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 18 1d 2b 33 38 49 44 4a 3f 42 3d 40 47 46 45 44 37 41 43 51 44 4f 4b 48 44 42 4e 4a 49 4b 4f 4c 51 4c 47 53
 56 4a 4d 4d 4e 50 44 48 50 4b 4f 52 49 45 4b 43 48 47 43 4f 47 44 4b 3f 4d 50 55 62 5d 64 62 54 52 4d 51 4c 4a 50 4f 55 5a 5a 55 52 4d 42 49 45 48 49 4a 43 48 4a 41 47 42 4f 4c 4f 44 4b 44 44 4d 4e 47 3d 43 43 3e 26 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 43 62 76 66 66 54 5c 61 61 62 64 69 68 68 6a 6a 68 68 6f 6f 66 6a 66 67 6d 68 62 5f 5f 62 5f 61 5b 55 55 5d 54 57 4e 52 4d 54 4b 4e 4d 41 51 49 54 46 47 4b 46 4c 44 4d 4b 47 44 43 43 47 4a 48 47 4d 50 4c 54 4e 4d 43 45 50 51 53 4f 4a 4f 44 47 42 3f 3e 45 37 29 1e 0e 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0a 17 22 31 38 3c 40 43 40 3f 44 40 43 47 47 48 46 42 42 43 3e 49 45 44 42 3d 3d 4e 40 44 4a 46 48 48 50 50 4e 53 4b 4a 45 47 46 4c 45 47 3d 4d 49 40 42 45 40 46 40 48 3d 43 49 50 51 54 61 5f 5b 51 56 4f 4b 50 45 45 4c 46 44 4d 56 57 54 4f 47 50 4e 47 48 43 47 47 45 41 48 40 42 45 4b 4e 4a 4e 42 48 45 49 4a 42 44 3b 45 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0a 36 5f 63 6b 6a 62 5f 68 5c 65 66 63 64 62 66 65 63 6d 65 69 64 62 6d 64 68 67 5f 5d 65 59 64 59 52 57 52 55 4f 4c 51 52 4f 4d 42 3f 4f 45 46 44 4a 48 41 50 50 43 4d 47 46 45 48 42 3f 48 4a 4c 4d 4e 45 42 4e 47 4c 4a 49 4b 4a 40 4c 48 50 4e 49 4c 45 46 48 35 2b 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0b 19 1a 21 3c 39 3d 44 3f 3e 42 47 46 43 3a 44 40 3f 43 41 45 41 4d 40 45 48 46 41 43 4e 4b 4d 52 44 51 50 4f 4e 4d 4a 48 4c 45 48 4c 46 4e 43 41 43 49 42 3c 43 45 46 42 45 49 49 48 4c 55 55 59 54 55 51 50 4f 44 47 45 4a 50 51 5d 54 55 4e 46 48 4a 46 3f 41 45 46 3e 4f 43 41 4a 43 44 41 4f 44 4f 47 40 43 44 4a 40 48 3a 26 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 37 61 5f 65 64 54 60 64 62 56 5c 5e 64 64 61 66 5e 64 6c 66 65 5d 6c 65 64 65 63 5c 60 5f 5c 5a 51 53 55 5a 52 42 58 51 4d 4d 46 3f 51 48 43 47 49 42 45 4e 45 44 4b 40 46 4a 46 45 44 4d 47 4a 47 47 4a 44 3f 4f 52 4a 49 4b 4f 4d 4c 4b 4a 4a 47 4d 42 4a 38 33 1e 16 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 14 26 2c 46 42 3e 46 46 41 3d 44 43 41 42 3c 3f 3d 3a 4a 46 47 44 3a 3e 45 44 4e 49 4d 4d 47 4f 53 54
 54 50 4d 4f 53 4d 48 4e 4e 4f 45 44 49 4b 45 51 46 46 43 46 49 42 3e 45 4b 4e 4a 53 56 57 56 47 4a 45 41 51 43 4e 43 4e 55 55 56 53 4c 4a 49 44 4c 48 45 44 49 46 3d 41 47 42 4d 4c 3d 4c 47 45 4c 49 4c 46 41 40 3f 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 37 59 66 65 64 57 5d 5e 5d 61 60 5a 64 68 5f 62 63 61 63 5f 63 65 6c 59 6e 5c 68 5f 64 5b 5d 5b 5a 55 4b 52 54 4c 4e 4a 47 47 49 45 46 49 4a 50 45 4d 49 44 4c 46 49 3a 41 51 45 48 41 4c 4b 48 44 4a 47 4f 4d 44 4a 4c 43 4d 55 43 4d 4f 4a 4e 40 49 49 49 38 2b 18 12 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 07 10 1d 2e 36 37 3d 42 41 3c 3f 45 41 3d 3a 43 45 3e 37 3b 42 45 45 43 3f 47 49 44 45 4a 3f 46 44 44 4d 4d 53 4d 4f 49 46 45 4e 51 41 4f 46 43 4d 45 48 4a 45 4c 47 3a 4c 47 46 42 4a 56 58 5a 56 51 46 4d 48 4b 48 44 4d 4b 47 55 52 53 59 57 4c 4b 48 49 42 4e 44 41 45 4b 44 4a 42 48 45 4e 43 4b 4d 4d 41 3b 48 48 46 41 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 30 5b 5d 65 68 58 5f 5e 61 59 62 62 66 5e 5d 60 5b 63 67 67 6c 5d 64 5e 65 65 61 5f 58 58 56 57 55 48 51 4c 4c 4f 4d 47 4a 53 46 49 4e 44 48 47 41 3f 46 50 50 47 42 3f 42 46 47 40 48 44 47 45 45 4a 48 4e 4b 44 46 4d 4e 4f 42 4e 49 41 4f 4f 45 4d 45 42 33 22 16 0a 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 12 1e 2b 30 42 40 3d 38 41 40 47 48 3c 41 3a 44 3d 3a 3e 4c 42 45 45 44 47 45 41 44 47 48 45 49 4a 4e 4b 52 4d 46 49 4d 52 4b 44 4d 3b 46 47 44 50 4b 4a 46 48 42 3c 41 45 41 44 4f 59 60 5d 5c 5a 57 54 4f 47 46 43 44 4e 4c 4f 52 51 54 53 50 41 4b 4c 40 49 46 47 3e 41 46 47 4b 4c 51 4a 52 41 48 40 49 45 44 44 48 4b 2d 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2b 57 5e 62 58 56 62 62 5b 5a 54 60 5f 5b 61 58 5e 5c 64 65 66 62 60 60 6b 5b 5f 57 5d 54 55 50 5d 55 50 55 44 4e 4e 4b 51 4e 4d 47 4a 4c 48 4a 49 42 47 41 47 44 48 4a 46 46 41 46 4a 44 4a 45 46 4c 41 4b 44 47 46 55 4b 4b 4c 51 46 54 54 4e 4d 3e 41 33 2b 1e 0f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 10 25 30 41 3d 42 3e 3e 40 46 41 39 40 47 41 3f 45 3d 3b 41 42 45 40 47 41 44 48 47 42 49 47 4c 4c
 51 49 4b 48 54 49 41 4c 44 49 4d 4a 47 4f 45 3c 49 46 44 45 46 40 47 3c 4a 4f 5d 5b 5e 5e 53 55 45 46 44 47 42 49 49 46 4c 4a 4f 50 53 50 51 4b 49 48 49 41 4d 42 48 49 46 49 4e 47 44 4b 4b 4a 42 47 40 4b 43 52 44 2f 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 21 58 68 5f 5a 58 5d 5c 55 5c 5c 61 61 5f 5f 63 64 64 62 5f 65 63 5f 5f 5f 5f 60 5b 55 5a 5a 56 56 56 4b 46 50 4c 50 4e 45 49 47 47 48 4b 4f 4e 46 41 46 4a 4a 4a 50 43 46 52 50 4c 42 43 47 48 47 4a 45 4a 47 4d 5d 4b 46 48 50 50 56 47 56 4d 44 4a 39 38 21 18 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 1c 27 3a 3d 38 46 40 3a 45 41 3f 3d 3b 45 3b 3b 3e 47 41 41 3e 3f 45 44 41 45 41 45 3d 43 43 4f 46 47 4b 45 4a 4d 46 52 49 4b 4e 4a 45 3a 4c 44 40 40 40 46 46 3b 42 41 40 4a 47 50 4c 53 5c 52 4f 49 3f 41 53 4b 4d 44 4a 4f 54 53 4f 4b 4f 4c 4f 4a 48 49 46 41 49 48 45 46 48 43 45 47 4a 4d 4a 3d 43 41 40 3c 45 32 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 29 50 61 5f 5b 59 5e 5f 56 5f 58 5a 63 5c 5e 60 59 56 62 61 62 52 64 56 60 55 59 53 50 4b 52 56 4e 4f 4f 4e 47 43 4e 40 40 50 43 43 4d 47 49 49 49 4e 41 47 43 4a 4d 4e 48 45 4e 4a 49 43 44 44 49 4a 4e 49 47 4b 41 4d 46 4a 54 52 4e 51 4e 53 45 3e 3b 2f 23 12 06 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 1a 25 3e 3b 39 44 35 43 3e 3f 3a 3a 3d 39 40 48 39 40 3e 3e 46 3d 44 42 3c 43 46 43 48 4b 4c 47 4e 47 42 49 44 47 4a 45 4f 45 44 47 42 45 46 46 4b 46 46 38 47 3b 3f 45 42 44 46 44 4f 47 4d 4a 3e 4b 4c 45 45 49 41 42 45 48 4c 56 47 4d 4a 4a 42 46 46 42 45 42 4b 46 3c 47 46 44 49 43 45 45 44 4b 3c 37 41 43 2b 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1e 4f 5d 57 59 5d 5e 59 5a 55 62 59 5d 5a 5d 5c 5a 5d 5f 63 5c 5e 5c 56 54 56 55 4e 51 49 58 4d 4d 4c 48 47 47 48 3c 3f 45 47 4a 41 45 44 4a 48 43 4f 3e 4a 50 42 4b 44 4b 48 4a 47 45 47 4d 47 44 46 4d 4a 4e 48 47 48 4d 4f 54 53 56 47 4d 42 41 40 30 2c 17 0b 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 18 24 37 3c 3b 3e 3d 40 39 3f 3e 3b 3e 45 42 37 40 41 3b 43 43 44 4d 42 46 47 48 3e 46 46 45
 43 4a 4b 51 4e 4d 49 49 4a 4a 45 49 4b 42 43 44 4a 4b 43 45 41 43 4b 3d 4c 41 45 45 3f 47 4a 4f 4d 41 44 48 46 4d 43 44 4b 47 44 4f 50 49 4d 4f 50 48 4a 45 45 42 4f 46 44 47 4c 4a 47 45 43 3b 4c 49 44 46 3d 41 3b 30 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1d 4e 54 5b 5b 5b 5c 5a 4f 5f 5a 65 62 5a 61 63 5e 60 62 59 61 5b 56 5a 54 53 51 50 51 4b 4a 4c 4a 4a 4d 4a 49 47 3c 4a 3f 46 4f 49 47 46 4d 4b 4f 47 4d 4b 44 4b 4f 44 51 48 46 4d 4b 4f 48 49 50 49 4d 49 4b 4b 50 47 54 58 4f 5a 52 4a 4e 4d 4b 40 2e 2c 19 07 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 13 22 2a 32 39 40 3d 40 3e 39 36 38 42 3a 35 3c 3c 3f 42 40 3d 3e 42 42 47 44 48 44 4a 48 45 46 4a 3d 48 46 4b 46 47 47 43 40 3f 41 4c 44 46 44 42 45 44 43 41 42 42 42 43 4c 45 3b 3d 4a 4a 42 44 47 45 47 42 4b 45 4b 4a 47 4a 47 4f 55 52 52 49 44 46 44 48 46 44 42 4a 4b 47 40 4d 43 45 44 42 3a 3d 38 3b 35 2f 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 4b 53 5c 62 58 5e 60 5e 5f 5d 5a 5a 58 64 59 5a 64 60 5c 58 53 5c 52 57 53 4c 50 49 46 4a 49 44 46 46 45 49 49 4b 43 44 4a 49 44 46 49 47 4b 4e 46 4e 41 45 44 4d 45 52 44 4b 4b 46 49 49 50 50 4d 4a 4c 50 4e 4c 55 5b 56 56 56 58 4f 49 49 40 41 2f 1c 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 1c 23 2f 30 32 3a 40 40 3d 42 37 37 42 36 35 40 3d 3f 3a 3d 37 37 46 46 3b 4b 42 45 43 48 48 45 3e 44 47 49 39 47 41 55 3f 42 4a 51 44 41 3d 43 40 45 46 3c 3f 3e 43 43 4b 32 44 44 4c 4d 40 3f 40 4e 41 40 41 47 4f 48 43 4c 4a 54 4b 57 57 4a 46 49 3c 48 41 46 49 45 45 47 45 3e 44 43 41 41 3b 3a 37 34 3e 2c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1b 44 54 5c 59 4b 5f 54 53 5e 5e 5b 5d 52 57 5b 5e 5e 5a 5b 5f 57 4f 4a 52 4b 53 55 4f 50 4b 4e 44 53 44 48 4d 48 4a 45 46 47 47 4d 4d 3c 3d 44 40 4a 3e 4d 4a 47 4e 52 4e 47 44 41 4a 46 4c 4e 49 4e 4d 4d 50 4b 4f 50 50 57 58 55 59 46 4a 45 40 37 24 1d 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0d 1c 28 36 35 3b 3e 3e 3e 3b 39 42 43 3e 3a 3f 38 40 43 3d 41 40 41 42 42 47 3b 3b 3e 47
 43 47 47 45 45 48 44 52 43 42 4e 49 3f 46 47 49 45 48 3d 4d 45 49 40 38 44 41 3e 43 43 47 4c 4e 4a 43 3b 44 3b 45 4a 45 48 42 48 47 45 4f 4f 55 55 52 4e 4d 41 4f 44 42 43 3e 4a 42 46 3b 41 3e 3d 3c 43 3c 45 3c 35 2e 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 4d 60 54 54 51 5b 59 54 58 59 59 5f 57 57 59 5c 5c 58 4f 58 52 5a 4c 4f 50 4e 4d 53 4e 4b 4b 48 47 46 44 48 45 44 45 4d 46 46 4b 4d 47 47 4d 44 45 3c 4d 48 42 45 47 4f 50 4d 51 4e 4b 4b 4e 49 4a 54 55 56 52 53 54 56 4f 53 54 50 4b 4b 3a 3a 33 1d 0f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 16 25 2c 2d 39 45 3e 39 3e 3a 38 38 41 42 38 41 43 3a 3b 3a 43 40 47 40 42 3f 3d 46 41 44 4b 47 45 45 3d 3e 4c 43 49 43 49 44 46 4a 43 49 42 3f 41 3d 46 42 43 43 3c 3b 48 47 47 4f 46 4a 46 44 48 48 3e 41 44 4c 46 49 4b 40 4e 4d 50 5d 52 4c 48 39 46 45 48 39 42 48 44 45 3e 3c 3f 36 41 3e 3a 37 38 3b 31 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 45 4f 51 56 50 59 56 52 52 5c 52 5c 5a 5d 59 59 60 58 54 57 55 50 49 50 50 53 52 4d 4a 4d 4a 45 42 44 48 4a 46 46 45 44 45 4a 47 49 44 42 4d 49 49 48 4b 44 44 4a 49 49 53 4b 4b 49 4c 4f 46 50 52 50 55 51 56 54 57 54 52 5b 54 54 41 40 40 37 24 1e 0f 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0a 1c 2c 2e 3e 37 32 3b 39 37 3f 35 3e 30 33 3e 37 48 40 40 37 3c 3c 3d 42 3b 41 3d 45 3c 4c 3f 46 3f 3a 3f 43 41 44 48 41 43 40 3a 4c 42 44 44 49 3d 44 41 43 43 41 37 48 3b 3f 44 47 3f 3e 49 45 4f 3e 43 4a 47 46 40 3f 42 4a 53 53 5f 50 4f 45 3f 44 3d 3c 41 42 49 46 41 38 3b 42 3e 40 3b 3b 3a 36 41 27 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 3c 54 4b 5e 4a 54 4f 4d 55 52 57 5b 5a 54 5a 52 53 52 4c 59 52 51 4f 4c 53 47 4e 4d 4d 4b 4a 42 44 43 43 51 4a 46 4d 51 43 45 4d 4c 46 49 4b 45 48 46 4f 49 47 4a 47 4e 4c 4f 56 53 4b 4f 5b 53 58 57 56 56 4a 52 52 4d 52 4f 43 4f 3a 3b 3f 30 22 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 0c 18 26 28 34 3b 32 3b 37 35 3d 39 44 32 3b 39 3b 41 42 39 37 47 3c 39 3e 3c 4b 46 4c
 39 41 41 45 48 46 3c 45 4a 45 4d 44 45 47 47 47 46 40 3f 43 47 43 3e 4b 48 40 41 3d 44 45 4b 3e 42 44 3e 46 3c 41 46 4b 4c 42 44 40 49 4c 50 59 60 58 52 49 43 4a 46 3d 41 48 43 40 3e 46 49 43 38 3a 3d 3d 3e 3c 3b 33 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 42 54 52 52 4d 53 58 55 55 55 5f 5a 5e 59 53 5c 50 51 4f 51 4c 4f 4c 54 4b 4c 48 46 52 4c 41 48 46 40 49 4c 48 42 4a 4e 55 4f 4d 49 49 47 53 54 4b 48 42 4c 4c 4a 4a 53 4e 4c 53 49 4b 56 56 4e 54 5e 50 59 58 5c 53 54 52 54 49 4f 43 3e 3b 28 1f 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 20 2b 2c 34 32 35 39 3a 38 2c 31 39 3b 39 3c 33 3c 3b 42 3b 47 3e 44 44 45 46 3c 44 45 3f 42 49 41 3c 44 3f 3f 40 46 46 3d 45 46 45 40 4a 3e 3f 46 46 46 44 43 43 42 3f 3c 48 44 4a 42 3c 3e 40 44 4b 45 46 43 4a 4a 4a 52 57 5d 63 52 51 53 48 43 44 44 3e 41 45 4b 40 42 41 3c 42 37 36 37 3a 33 34 38 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 37 4e 4e 51 50 50 5a 4c 53 56 4f 60 58 54 51 5a 52 52 4e 4d 4f 4f 48 48 49 4f 47 43 4e 4c 47 4a 43 4a 49 51 4a 4d 44 50 4f 45 49 4e 4a 40 47 49 46 47 54 53 4f 4a 4c 54 4c 4b 57 50 47 4a 59 59 5a 50 57 5a 48 52 4e 4e 4f 55 4d 50 3c 3c 27 1e 1e 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 1e 2d 2d 2d 32 3a 3b 31 3d 3a 3c 33 41 3d 37 38 40 44 3d 3d 46 49 3d 41 3f 3b 41 3f 40 43 3d 3d 47 3e 4a 45 41 40 44 44 40 47 46 46 45 42 37 48 49 44 4e 4a 41 3f 42 45 49 4e 4a 36 3e 44 45 38 3e 3f 3c 47 47 46 4d 56 52 64 68 5b 51 4a 4b 48 44 48 3d 44 3b 3f 40 40 3c 3f 3a 3d 3c 3a 3c 3a 37 33 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 3f 4c 4d 47 4d 50 50 52 54 50 5b 4f 58 58 54 51 51 4d 4f 47 50 48 4b 51 4e 50 47 4a 49 3c 4a 46 3e 45 46 44 43 4a 47 47 4a 49 4a 47 4a 4e 4d 41 4d 50 52 48 4e 55 49 5a 56 54 54 5a 57 54 59 54 5a 53 54 53 4a 50 50 51 4a 49 46 43 42 30 2d 18 0c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 19 25 2f 27 2d 35 32 38 36 38 3e 36 37 2e 36 38 3b 42 45 41 42 43 4a 3f 45 46
 3d 45 4a 36 41 3d 42 46 45 3e 48 46 4a 44 40 44 44 45 44 45 3e 42 45 3e 46 41 41 3e 42 41 50 3a 23 2f 48 46 41 3c 38 3f 40 45 41 41 41 51 58 63 6a 59 57 4a 42 41 44 3d 46 40 3e 3e 44 49 38 3b 44 3b 3e 3d 37 3f 30 37 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 3b 47 54 54 4f 4b 54 4f 50 53 50 56 4e 54 58 54 45 52 55 49 4a 4f 4b 4c 44 4a 4e 44 46 46 40 42 49 42 4e 48 43 3e 3f 4c 51 46 45 52 49 4c 51 4f 51 51 51 51 50 50 52 5a 50 55 58 5c 5e 57 58 52 4e 4e 57 51 53 4f 50 55 49 40 4a 42 37 30 24 13 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 11 1d 27 30 2e 36 2e 32 39 37 38 3b 35 3e 3a 3f 3e 3e 40 41 3d 41 44 40 43 3f 3f 41 40 44 42 42 41 44 41 43 48 40 4c 43 3a 44 45 3b 46 41 47 46 41 3c 48 3e 3c 46 3e 46 42 41 45 46 48 40 3c 41 40 40 44 3e 3c 44 42 4d 55 54 55 50 47 4d 51 4c 47 4b 41 45 45 43 38 40 3e 41 3d 3c 3f 3f 35 37 39 2e 1a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 32 4c 4a 4e 47 50 54 44 52 50 4d 55 50 57 54 4b 4c 46 45 43 48 4e 50 46 4a 4d 49 42 43 4b 51 4a 3f 47 4c 48 49 4b 52 53 4d 4d 4e 45 43 51 52 4e 4a 4f 49 5b 4c 4f 57 61 4f 59 5b 5d 5e 58 5d 54 4c 4f 4a 58 45 50 3d 4f 45 4b 50 41 33 2b 22 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0a 16 2a 2f 2c 37 36 2a 34 34 39 37 3d 3c 3b 36 3e 3a 3f 32 41 42 3d 46 3c 40 3d 3b 3d 3c 40 49 3e 43 44 3e 3d 39 44 4b 3e 40 45 43 42 3e 44 48 3f 44 46 49 3f 45 41 3d 4d 45 3e 3a 3d 44 37 3d 40 35 42 42 40 43 3d 4a 4b 52 57 4f 48 44 4c 47 3f 47 3c 3d 40 3a 40 45 36 42 40 3c 40 37 30 3a 30 2e 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 36 41 4c 57 47 50 4a 4e 4a 50 4c 53 49 50 4a 49 49 49 4a 47 47 50 41 4b 49 49 48 45 3c 44 43 46 48 44 4d 43 49 46 46 45 4e 53 47 4d 41 4e 52 53 4f 50 51 53 4e 4e 52 5b 52 5b 55 59 53 5b 4e 54 45 4f 4e 46 48 4a 46 46 44 4a 46 3d 28 21 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 04 06 11 20 23 30 30 2e 2c 36 31 38 32 39 32 2f 3b 3e 44 3e 42 3f 3c 3f 39 45 44
 3b 3e 4a 3b 45 3d 42 40 3f 42 40 41 3a 47 46 46 3e 40 40 4b 3a 40 3a 3e 44 4a 3f 3b 43 3b 41 45 44 3d 3f 45 3d 3c 3b 3e 38 40 48 45 40 42 3c 45 4c 4f 4c 4b 49 4c 3e 44 44 3d 40 46 44 3e 43 3b 3b 38 30 3d 3c 30 47 2f 18 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2e 4c 4c 4e 46 51 50 53 4e 4d 47 48 4f 4f 4d 46 4a 4d 4a 44 44 47 41 45 46 44 3f 44 47 4b 49 47 48 4c 4a 46 43 47 4b 4a 42 50 53 4e 4a 4f 4c 4c 52 58 4e 53 5c 59 60 56 5c 5f 5d 5b 51 4b 52 50 4c 4d 50 4c 40 4d 44 45 48 49 44 3d 2d 18 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 1b 20 2c 2a 31 36 30 2f 37 33 34 35 32 3d 3a 42 36 41 40 3e 43 3b 43 44 43 3d 45 40 40 3d 41 46 41 40 40 47 42 43 40 44 3f 47 3e 44 43 3f 42 44 44 38 42 45 42 42 44 44 44 42 4e 45 3c 46 3f 48 4a 3d 43 40 3e 3e 4c 41 3e 3f 4a 4f 52 50 49 44 42 3d 3f 43 36 3c 41 3f 3c 41 37 3e 3c 38 39 3a 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 33 49 42 50 4c 53 49 56 4c 4e 4d 5b 49 47 4b 4b 41 45 42 44 48 4d 4b 4e 41 47 4c 44 4a 46 45 47 49 4b 49 49 4a 41 4d 4a 4a 54 4d 4a 4d 54 49 52 57 52 5f 55 52 5c 5b 5d 55 5c 59 57 52 51 53 4b 52 50 54 4e 43 4c 40 49 44 45 37 2d 22 1a 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 10 17 19 2a 24 30 39 32 38 33 3b 33 3b 34 39 36 3c 3a 40 43 40 42 3b 47 45 3b 3b 40 3e 41 44 44 3a 41 45 40 3f 42 3d 3d 45 3b 4b 44 41 45 44 41 3f 46 48 4c 3c 36 3e 3f 45 42 42 42 3d 3c 3e 3e 49 3c 36 3c 3d 45 42 46 42 47 4c 45 42 41 40 39 3c 3d 44 48 41 44 36 3f 3f 3c 31 3f 3d 3d 41 37 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2c 42 42 4c 4d 54 4a 48 48 46 47 4a 48 47 41 4c 40 43 44 49 46 4b 46 44 3d 46 3b 47 4e 4a 4f 4a 43 51 49 44 4d 4c 51 50 51 50 4d 54 54 50 59 55 4e 52 56 5e 50 55 55 5e 56 54 53 4f 4b 50 49 4c 49 4a 45 4f 45 46 47 3f 49 3d 2f 2f 16 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 22 32 2b 33 2d 30 33 33 36 3a 38 2f 3b 35 45 37 3c 40 3f 3c 3b 3a
 3b 40 44 37 42 3e 3d 3d 42 3f 41 42 3a 3e 3e 40 50 41 3e 48 41 43 4a 44 4d 3e 3d 41 40 3e 3d 3d 49 3d 40 45 44 3a 3e 46 42 37 44 38 37 41 37 44 3f 3d 45 4b 4e 46 45 42 45 3a 38 3f 3f 3f 37 40 3e 43 40 3a 34 2e 34 31 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 41 49 54 47 55 55 4f 44 47 49 48 50 47 49 45 42 4e 41 47 44 43 44 44 45 46 48 42 4c 46 3e 45 47 4e 52 50 41 49 57 4a 4f 4f 46 54 51 4a 57 4d 58 56 59 5d 54 5f 59 5a 55 54 58 4f 4c 4c 48 48 4b 50 3e 48 41 41 40 3d 37 33 38 27 16 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 15 16 24 2e 38 2e 35 34 41 32 34 3b 31 3b 3d 44 43 42 43 40 40 3e 3a 42 45 40 45 40 42 41 42 3d 3f 44 3c 3f 47 40 42 40 3d 46 48 42 4c 4e 46 46 42 43 42 47 3c 40 3f 42 3e 3e 42 3f 3e 3f 43 42 3a 40 44 3e 3d 3e 48 40 48 41 46 41 50 45 43 3e 44 40 43 43 42 3f 42 39 36 3a 40 41 38 38 34 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2f 49 4a 50 47 48 48 47 4c 4c 4d 43 47 4d 47 49 40 4f 4a 53 3f 3f 49 47 43 4b 4a 4f 4b 45 4b 4c 4c 51 4c 56 4b 57 4c 54 58 54 55 50 5c 53 52 55 5e 58 60 56 57 5e 4e 5a 52 50 5e 51 45 4a 4b 57 52 51 49 44 3c 45 40 3c 3b 2d 28 20 0e 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 10 25 2d 30 34 2c 3c 3c 3d 3f 36 3e 3b 3e 3f 3b 43 40 3e 3e 47 3a 3b 4b 41 43 45 44 40 43 46 41 40 47 47 46 3e 46 40 3b 3e 3f 3b 44 43 49 43 40 4a 44 42 42 3d 42 49 47 49 47 4b 3e 3b 3d 3c 39 46 3b 3f 3a 3d 3f 3c 42 44 44 40 47 3c 44 41 40 3f 43 41 3e 40 44 40 3d 3e 35 38 39 43 3a 23 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 25 41 4a 55 4b 4b 4c 48 4e 43 47 49 44 4c 49 4c 42 4d 47 4c 47 3d 4a 46 44 45 45 4f 42 51 4a 54 4f 54 53 50 54 51 48 52 52 53 54 54 4e 4c 5d 5a 5d 61 5d 57 58 59 55 52 51 4a 45 51 4e 5c 4a 51 4d 4b 43 4d 40 39 38 37 3f 29 24 1e 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 1a 26 32 37 37 2f 3f 3a 43 3c 43 3e 37 3e 3a 41 42 41 3f 3a 40
 49 43 3e 41 3e 47 41 42 3d 3c 43 47 39 3c 40 4b 3c 44 42 47 3d 47 45 43 45 40 42 46 43 3f 3f 43 3f 45 42 45 3e 3c 40 40 3c 3a 3f 3c 39 37 3b 41 3f 39 3f 3f 3c 3f 49 40 42 42 47 49 42 46 35 3d 38 41 41 39 33 3c 32 35 26 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 1f 43 49 4d 49 46 46 46 44 4e 40 51 3d 47 47 46 47 41 42 40 40 4a 45 43 47 4a 46 43 44 46 51 49 4b 4d 50 49 54 4c 4f 54 4f 4e 4e 4f 52 51 58 5b 5c 58 50 4f 4c 55 51 50 58 51 51 54 4a 49 44 4a 4c 4f 4a 48 45 3e 37 3c 34 23 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 10 26 2f 39 3b 37 3a 3b 45 4b 47 3f 3d 37 35 40 3e 3d 3f 41 4a 3e 3c 3f 3c 39 42 3f 40 40 47 43 3c 37 44 47 46 47 3b 42 4d 42 3d 49 41 41 47 44 49 42 42 41 4b 45 45 3e 3c 41 40 3e 43 40 3b 3f 39 38 41 33 42 3f 38 38 41 41 42 44 3e 39 46 40 4a 43 45 43 41 42 45 3c 41 3a 3f 3a 34 22 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1e 40 4c 52 46 41 45 42 47 49 47 46 3f 46 3f 47 47 45 4b 3e 43 4b 4a 4e 49 59 41 47 4a 4d 53 52 4d 4a 50 49 4e 52 55 55 55 59 4a 55 52 58 61 5c 59 5e 5a 5b 52 4f 4e 56 55 48 4d 4d 49 51 4a 50 53 53 4b 53 42 3c 3d 2c 1e 21 11 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 11 27 2e 3b 33 30 3e 47 47 45 43 40 35 3d 3d 3d 3f 3a 3a 47 49 4b 3b 3d 42 44 3f 3f 42 48 3e 47 46 46 47 45 47 45 43 49 3f 48 48 43 45 42 40 4a 45 4d 4c 47 45 46 46 3e 3f 3b 3e 44 41 38 3f 42 3c 45 35 40 3e 39 3a 3e 32 47 3d 44 3d 47 4a 4d 50 43 3a 35 3c 39 3e 3f 3d 42 38 3d 2b 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 3f 48 4c 45 44 4a 4a 42 47 43 49 41 44 48 44 43 42 47 4d 45 47 4f 4a 47 52 4b 4c 49 52 4d 55 49 55 52 4b 50 50 4d 55 51 56 5c 54 58 59 5e 5c 51 55 55 52 52 51 4d 4a 53 4f 50 4c 48 56 53 4d 57 54 47 4e 43 3f 34 32 21 12 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 1a 2c 33 35 36 37 44 3f 45 3f 3d 36 35 39 40 41 3e 3f 3a
 36 44 39 3f 3a 3e 3f 43 42 4b 44 43 45 45 43 40 3f 3e 4c 49 43 45 44 40 3d 41 39 43 3e 45 40 43 42 3f 3f 43 3e 45 41 44 3e 3a 3c 3e 38 3c 3b 3f 3b 36 3c 38 3d 3d 37 3b 40 42 4f 4e 4f 4c 47 3b 40 37 48 37 3b 3d 3e 33 24 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 23 38 3b 4b 3f 45 41 48 47 47 50 4c 4c 47 41 49 49 46 46 45 44 48 49 46 4d 4e 41 53 4d 4c 49 4f 4e 4f 51 51 4d 4d 56 50 52 52 58 5c 56 53 4e 62 51 4d 52 53 4b 4e 4e 53 55 50 4d 44 49 45 51 51 52 53 4b 49 36 35 2e 24 16 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 12 27 25 2f 36 3a 3e 4d 45 41 3f 3a 37 40 43 37 39 3a 34 3d 40 39 3a 39 3c 42 39 45 3c 41 3f 3f 44 44 3e 42 41 48 45 47 42 45 40 42 40 47 43 42 45 49 3c 47 48 46 4a 38 42 44 43 43 3f 45 3e 36 3c 43 3e 47 39 3f 40 40 3b 39 35 3d 4d 4e 56 59 4b 41 42 3b 3a 48 3f 42 45 3f 3c 26 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 40 4a 4a 40 40 51 47 4b 52 55 4e 4c 40 42 4b 42 44 47 45 44 49 40 46 43 46 4d 41 4e 49 54 53 46 4f 4c 56 4a 4c 53 4f 55 51 5a 5a 5d 58 52 51 51 4f 4d 4d 4d 59 50 54 4c 45 4e 47 45 4f 4d 4e 58 5b 50 48 36 2f 29 1a 0d 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 1a 38 35 3c 3d 3a 40 49 40 44 35 34 40 39 42 41 37 3b 3b 44 37 43 3d 3e 3e 42 44 4e 3a 42 40 42 47 49 47 43 44 41 3f 48 41 41 45 43 4c 42 40 3d 42 4a 42 45 4f 41 46 41 3d 3f 40 4b 3d 44 39 3b 40 3c 3e 45 3c 40 40 46 40 40 3e 3a 4b 4c 50 50 42 47 45 45 44 41 3e 43 3c 40 26 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 45 4a 46 42 49 42 49 4e 55 52 4a 3d 49 3f 47 46 4e 4b 4d 46 4a 45 48 42 4e 49 49 50 4d 50 4a 52 55 4d 52 51 54 5d 51 4e 56 51 51 50 4e 50 51 50 4c 49 4f 46 4c 53 4c 49 44 4c 47 4e 54 4e 4e 4f 5e 51 43 33 29 17 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 17 19 21 2e 35 40 39 43 3f 3c 3d 35 38 33 3a 34 34 3a 3b
 42 39 43 3c 41 44 3b 40 3c 39 43 48 40 40 3e 41 50 3e 4a 44 47 3e 40 47 41 47 48 40 3e 3f 3f 3e 45 3d 42 44 3f 40 3f 3f 40 47 46 40 3e 38 3b 3b 38 37 3d 3d 3e 45 3a 3b 3a 3e 3b 54 51 4c 3f 43 45 48 47 44 49 42 3a 3f 38 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 3e 4b 4e 4e 4c 45 4d 4d 50 47 4e 4a 3d 47 44 49 4c 41 44 40 4b 4d 44 4d 4d 48 44 4a 4e 4e 53 47 46 52 52 52 4d 55 54 55 47 52 4f 49 50 51 4b 4d 54 4a 4b 4d 4d 43 4f 44 4f 4c 47 4e 4f 47 4e 42 4b 47 37 27 22 18 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 11 1a 31 44 42 42 3b 45 42 3d 34 36 3d 39 41 3f 39 37 3e 3a 43 3e 39 3d 40 3c 3a 47 41 3a 44 47 44 44 46 47 4b 44 3e 4b 47 47 49 3f 47 4c 3d 42 4b 42 48 42 45 45 45 41 4c 49 3e 40 45 3c 42 41 3e 45 3c 42 44 3d 43 47 3f 43 45 44 45 4d 4c 4d 50 45 4a 45 43 3e 3f 46 4d 40 35 11 06 05 03 02 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 3f 45 45 3f 4c 48 45 4a 49 4b 4a 4b 4f 42 4a 4a 45 48 45 47 4e 47 4c 4a 50 4a 4b 4e 56 52 4e 46 52 50 4b 55 4f 5a 55 52 54 49 4c 50 4a 4e 52 4e 4e 50 49 4e 53 4c 52 48 42 54 50 4f 49 44 48 58 49 3b 2e 24 1b 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 10 24 36 38 3d 3d 3e 3b 35 39 3a 34 35 36 38 3a 3a 3f 3f 3a 41 3a 42 39 3f 39 45 43 3e 43 45 40 4d 40 40 43 50 3b 3d 4e 45 47 51 3e 4c 45 42 3d 43 4c 41 4e 47 3f 42 40 44 46 43 45 41 3c 3e 3a 45 3d 40 44 39 42 46 40 3d 43 46 47 51 49 59 50 46 44 41 42 3c 41 3e 4d 41 3a 14 06 05 03 04 07 08 03 06 08 0a 05 05 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 3f 44 48 46 46 4f 49 4a 45 46 45 42 47 47 4b 47 44 42 48 41 4d 47 4b 4a 4d 4f 4b 57 56 54 56 4c 4c 54 50 48 44 4e 49 4a 4b 4a 46 55 51 4f 50 4a 46 4f 4e 3d 54 4a 4a 4f 46 47 4d 45 44 47 48 48 3f 35 24 1c 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 25 25 3f 3e 45 3e 34 3a 32 34 31 2e 30 36 3b 3a
 40 37 38 37 43 41 3d 38 3f 3f 40 42 41 47 49 47 46 45 42 45 3a 4e 44 44 42 46 4a 44 44 41 4b 45 3c 45 43 43 4c 43 42 48 43 45 42 47 3f 3a 41 44 44 3a 3f 43 3d 3f 41 42 43 41 46 4a 4b 51 4a 47 45 42 43 45 4f 4b 4d 43 37 20 0a 05 04 0b 0b 0b 03 0a 09 0a 11 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 3a 46 4e 46 45 52 42 43 4c 40 44 4a 46 4e 46 44 46 48 49 3a 44 4b 50 43 51 4c 49 4f 4b 4e 4e 48 49 49 4b 4d 47 4a 51 48 52 4f 4e 49 52 56 52 53 49 4a 4d 47 48 4e 4e 4c 44 49 42 3e 49 46 43 3f 33 32 1c 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 15 29 2f 3b 39 3e 38 36 35 38 38 3b 39 35 32 3a 3f 41 3d 34 37 3b 3b 3e 3d 3d 41 3a 44 41 49 49 44 46 3d 4b 40 4f 43 3f 3e 40 3c 43 40 44 3c 45 45 40 46 44 48 48 48 49 47 38 4c 3c 47 47 44 42 42 41 3c 42 41 39 41 3e 49 48 49 4a 49 4d 4e 46 45 43 53 53 52 4e 4d 46 42 1f 0d 0e 05 11 09 0f 16 18 15 1d 18 10 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 41 45 4d 3d 40 43 44 48 44 44 4f 45 44 3f 44 46 49 3f 48 47 4e 47 4e 49 4e 4c 51 50 50 4d 52 46 45 51 4a 4d 44 4e 47 48 4c 4b 50 4b 4a 51 4f 54 49 49 4d 47 43 47 48 46 41 48 3f 3d 44 41 3e 43 33 22 12 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 16 26 30 33 36 38 35 36 38 3c 36 35 37 3f 3c 3b 39 41 3f 39 38 3c 3e 41 42 3f 43 49 41 44 47 4d 45 47 44 48 45 47 44 41 48 41 48 42 43 45 45 4b 41 43 48 4a 42 44 45 4a 4a 45 42 4a 3e 38 43 42 46 3f 44 45 42 3d 40 4a 46 4c 4f 49 52 4b 47 4a 4d 4a 4b 4b 50 4b 4d 4a 2c 1d 18 10 12 1a 20 21 28 1b 20 20 13 16 06 04 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 3d 3d 4e 40 41 3d 3f 44 48 41 49 42 3f 49 4b 51 44 4e 4f 46 48 48 55 54 53 4f 4a 4b 4c 4e 4e 47 45 50 4a 42 4a 45 4c 50 4e 53 50 4d 57 50 5c 53 4f 44 45 43 48 4c 4a 4a 4b 3e 41 3f 47 41 42 2b 26 15 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 06 18 29 29 32 32 31 34 41 3c 34 3e 34 37 3e
 40 38 3d 40 37 3b 42 3b 45 45 45 44 44 41 41 48 4e 49 42 49 47 49 3f 3c 4f 45 47 43 3d 48 44 43 46 49 41 46 41 45 41 45 4c 3b 3c 3e 3c 3c 3f 44 3b 45 43 3f 4a 3e 48 50 48 4b 47 4a 52 53 50 4c 4c 54 52 53 55 4a 56 51 44 2f 18 0b 11 16 1a 1c 20 22 29 21 22 1a 15 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 2f 3e 44 47 41 4a 45 3d 47 41 4b 40 44 46 48 4d 48 51 48 4d 53 4e 4e 4c 53 4f 46 4f 46 49 47 41 41 3d 44 4b 4f 47 4e 4a 4a 51 52 5b 5d 5a 5b 4c 50 45 43 40 47 3e 45 40 3a 3f 39 3e 3e 3d 2e 23 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 15 1c 23 28 2d 36 3b 37 32 41 2e 2f 3d 2f 3b 39 35 37 3d 34 3e 41 3d 44 41 49 3d 49 49 4b 43 49 4d 45 45 46 4b 44 49 45 3a 44 40 45 44 45 45 43 45 45 43 44 44 43 45 3e 4b 44 41 4b 40 43 3c 3d 39 3f 44 47 47 46 4c 48 50 53 4c 4e 53 4e 57 4e 55 4c 52 52 4f 4e 40 39 25 16 16 22 20 23 1f 25 2b 2b 1f 1e 16 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 2e 37 3b 3e 3f 44 45 41 42 49 44 4a 48 53 49 47 4b 47 4d 52 54 48 47 4a 4b 47 45 47 4f 47 40 46 41 4e 48 48 43 49 4f 4d 51 60 63 60 55 56 4c 44 4d 4a 46 44 42 40 49 3a 3f 3c 3d 3c 3d 30 25 1a 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 13 1f 24 34 32 32 3a 37 3e 3a 3a 35 39 39 3e 3e 3e 3c 3e 3f 40 40 46 49 49 40 50 46 4f 4a 43 50 4c 43 4a 47 45 4d 43 47 4e 3a 44 49 44 49 4b 47 40 42 3c 4a 45 44 43 44 3f 3b 4a 47 42 49 47 3f 48 3b 47 4d 45 4b 54 5a 51 53 5d 5b 5a 5c 5f 60 60 5b 53 58 57 4e 41 28 25 22 1b 29 25 27 32 2a 22 25 27 1e 0b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 32 40 44 38 43 42 41 47 42 54 52 4e 4b 42 44 4f 46 51 51 48 49 41 45 4a 4f 53 4a 4a 48 48 45 48 47 4a 45 48 4a 53 50 5a 55 5a 5e 5a 58 55 49 44 46 46 3c 43 3c 3f 41 3b 3a 3d 42 39 37 29 18 0d 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 13 1d 28 2c 40 31 32 39 34 2e 34 40
 37 3f 30 36 37 3e 34 42 42 3f 46 44 49 4e 4a 43 44 4c 44 46 4c 4a 4c 46 46 43 41 47 47 47 49 4a 40 4b 47 48 3d 44 46 42 44 3c 48 3f 42 48 44 42 48 44 43 47 48 4d 4f 4d 54 50 5a 53 52 5e 5f 62 62 5e 5c 62 5c 58 60 58 51 3b 2a 26 22 20 22 2b 24 29 24 27 20 29 1f 10 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 38 47 40 45 42 44 4d 48 4c 44 4d 4a 46 4f 4d 51 45 42 43 49 46 4d 57 47 51 4e 54 4a 44 4d 45 54 53 4c 4f 54 4a 54 54 58 5b 62 53 4c 47 48 43 46 3c 43 3e 35 3e 3b 44 3f 40 32 31 2e 1b 09 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 18 1b 2a 3a 33 32 37 33 3d 37 30 3b 3c 3c 3d 38 45 38 3e 41 3e 41 43 48 49 42 3f 3f 41 40 49 49 49 4d 3d 48 47 48 46 45 45 43 49 48 45 4b 47 41 45 4a 43 45 4b 50 48 45 44 4b 49 43 45 47 4b 4c 53 56 53 5c 59 5d 62 67 5d 65 64 66 62 62 57 60 56 5a 60 5b 45 2a 24 1a 21 23 22 29 22 24 2a 24 1d 0b 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 30 3b 43 41 48 4a 47 40 4a 53 4c 50 49 45 4c 44 50 43 47 43 44 4e 4f 53 5b 4b 4f 4d 46 41 51 5b 5d 58 54 52 4c 4a 49 50 55 4e 52 4a 42 44 3f 43 41 41 43 3a 39 35 3d 3f 41 3c 33 23 16 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 1d 22 2f 3c 37 3c 34 34 3b 38 44 41 3b 3b 39 43 42 43 3d 3f 3c 42 41 4c 45 40 47 40 49 48 46 4a 4b 48 4c 52 40 4a 4a 42 49 47 44 41 42 48 41 41 42 45 46 47 40 43 53 49 4f 52 54 4d 4d 4d 52 57 5a 55 5d 5b 6f 68 6a 64 66 69 65 69 65 63 5a 5e 61 58 53 45 2a 29 29 20 23 27 23 28 29 25 1d 21 10 0f 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 25 39 40 3f 43 44 3e 46 4a 48 4d 49 4b 52 44 48 48 3f 46 45 45 56 51 5e 5a 52 51 55 54 5e 65 64 5a 5d 57 4c 41 43 44 4c 4e 45 47 47 41 49 40 41 3c 41 3b 3d 35 37 3d 3e 34 35 28 1e 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 14 22 30 35 3b 36 3c 3d 35 45
 3e 45 36 35 35 46 3c 45 40 46 36 3f 3b 47 48 3e 48 49 45 52 4d 45 49 4c 4e 46 4a 49 43 4b 48 51 53 48 4d 4a 42 52 49 49 4c 4b 44 51 55 53 49 4e 55 53 56 57 54 56 5b 54 68 5f 66 6a 6d 71 73 6c 66 6d 68 66 64 5d 5a 56 59 48 26 1f 1e 1c 1c 2d 25 27 25 23 1f 17 0b 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 22 3d 46 3d 49 47 4c 4d 46 4c 50 45 46 42 44 48 4a 48 53 45 52 50 54 52 5d 4d 49 52 52 5f 5b 5c 56 56 4d 45 41 40 46 3c 3f 47 2f 4c 46 3c 44 39 3a 36 40 38 39 39 3a 32 31 2f 21 0d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 17 2e 36 3e 3a 34 35 39 41 38 34 3a 38 3e 39 38 40 3e 3f 46 3f 3c 43 41 4b 4a 45 49 4e 4a 4c 40 4a 49 4d 4c 44 47 49 45 48 46 47 4f 4b 43 41 47 49 4e 4a 4e 55 54 55 60 62 5f 55 60 57 5e 60 59 65 70 70 74 6f 69 70 6e 70 6a 6b 67 65 5b 59 54 52 48 26 1b 1b 12 1e 25 23 20 22 1c 0f 14 0e 09 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 22 40 3a 3b 43 45 3c 44 43 47 49 44 45 45 49 4b 46 48 3f 44 4e 53 54 59 58 55 5b 50 5d 5e 5f 4e 4d 4d 3e 40 49 3b 3e 45 3d 44 46 39 3b 3c 39 32 3a 32 39 3b 36 33 39 34 2b 26 1f 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 1d 26 2d 35 3a 34 3b 3a 35 39 3e 37 37 45 3a 40 3a 43 41 3f 3a 42 3c 44 4a 4e 44 44 48 50 4f 4b 49 4b 4d 44 4a 4c 50 45 48 49 47 4d 49 49 4d 47 48 4e 46 59 5c 58 5a 62 69 64 66 69 6a 69 65 6b 65 6d 6d 6d 6b 73 72 73 6d 68 66 6b 5d 5c 64 61 58 42 29 1c 1c 16 1c 14 21 29 27 1c 1b 0f 06 06 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 3b 42 3e 38 44 3c 48 3f 3b 49 42 46 49 46 48 43 4b 4a 48 53 4e 5c 54 5f 55 5d 60 65 60 5e 5a 4f 4d 43 3b 3f 41 3b 3d 34 3f 3d 36 3e 39 44 3f 34 3d 37 36 3e 33 32 27 19 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 1d 26 36 3d 37 3e 38
 39 3d 3d 39 37 3e 37 39 3c 40 3a 44 43 3e 3d 41 45 43 41 48 42 4a 4e 4b 52 47 4b 47 4a 50 53 51 49 4c 4a 53 47 46 43 4e 49 4b 51 5b 60 67 5e 6b 6f 70 6c 77 75 6b 71 72 6d 6c 7b 6d 75 77 78 70 71 70 64 64 5d 69 5f 60 4a 4b 27 1b 1b 1c 12 1b 20 1f 15 14 0b 14 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 33 45 3d 3a 3f 39 3c 41 3e 43 46 49 41 44 46 47 4b 53 52 56 58 61 62 68 6f 62 6d 72 6a 62 54 4d 45 3b 45 3e 3b 38 35 3b 39 44 3d 41 3d 35 3b 3a 35 34 34 35 2d 26 25 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 20 23 2a 30 32 34 3b 38 41 37 3d 38 32 3e 43 3f 3a 44 38 39 3f 41 3d 40 43 4e 41 46 4c 42 4b 47 4a 42 48 42 44 4c 53 46 44 4c 46 45 4c 48 4e 47 5b 57 5e 68 62 75 78 79 73 72 75 75 72 72 77 72 74 75 76 76 77 81 73 71 66 6a 66 62 62 63 55 46 2c 1e 18 20 11 1c 18 0f 1d 17 13 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 1c 36 39 37 3c 40 40 36 3f 3e 42 45 46 46 44 4e 4d 51 5d 64 66 69 6c 6f 6f 6b 70 6a 68 66 55 54 48 3c 3d 33 36 3f 40 3d 38 37 3c 3c 36 38 36 3f 34 35 2f 2f 29 1c 1a 13 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 15 25 1d 31 33 3a 3b 3e 3e 3c 44 39 3e 33 34 4d 43 44 42 3e 41 42 41 41 48 44 4b 3a 44 46 4c 45 51 53 4f 43 4a 47 49 47 4a 51 3f 49 46 44 47 51 51 61 5c 6a 6b 7b 75 7b 85 7e 78 7e 7b 77 74 6f 79 77 7b 79 76 79 71 6d 72 6e 65 67 6b 5f 5c 53 27 14 12 13 1a 1c 1e 1b 0e 15 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 16 31 3e 39 42 3b 45 3c 42 48 4e 43 4e 42 4c 57 58 66 63 6c 69 6b 78 78 7d 6f 73 71 61 62 5a 48 48 35 41 39 38 41 3f 41 2f 3b 35 3a 3b 41 3a 36 3d 34 37 2c 24 18 16 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 1a 1c 2a 35
 37 37 40 3b 3c 3f 38 40 38 37 41 40 38 45 43 44 41 42 49 4b 43 4a 49 4b 44 4f 49 47 47 42 4c 48 4b 4b 50 4c 4b 4d 49 51 56 56 5c 5c 64 70 66 76 7d 81 7f 85 7d 7c 7e 78 79 78 6d 76 75 78 7d 81 7a 70 72 66 66 68 65 63 57 4f 27 05 1e 18 1a 21 15 13 14 0d 09 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 34 3f 3c 46 39 45 45 43 47 49 46 4e 56 56 66 62 6e 77 71 78 76 73 75 75 68 70 6a 5d 5a 4b 43 3e 3d 42 3d 3b 38 35 36 31 39 36 39 3f 35 36 3c 2d 33 35 27 17 18 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 15 23 28 2e 34 32 3d 3e 36 37 34 3d 3b 3d 39 40 49 48 40 46 49 44 45 4a 3d 4c 4f 55 53 52 55 4b 4c 4d 4a 4b 54 52 49 47 4d 4e 51 53 4e 54 5b 64 69 72 76 77 7a 7e 86 85 80 82 7b 73 7e 6b 78 72 79 79 79 78 73 75 6d 65 65 6d 58 57 49 29 05 1a 16 14 14 0b 14 09 0b 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 3a 3b 2e 45 3f 3c 3b 42 47 4e 47 48 51 5f 69 6e 6d 76 78 78 76 79 6b 6a 6b 61 5c 4e 4e 4e 3c 3c 39 3d 39 3a 31 39 3d 3e 3a 36 35 33 3c 34 30 2e 2f 2a 19 0f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 1a 1d 28 30 2e 37 36 3f 38 44 40 4c 4b 53 48 48 4b 48 4a 4d 55 45 4c 4e 41 53 53 54 52 52 53 56 55 59 52 58 51 53 52 59 50 54 57 50 5a 64 5f 66 71 71 78 76 78 83 80 81 7b 7c 7d 7c 7f 81 72 7e 76 7b 7b 71 6f 70 70 63 66 5d 60 4e 32 1d 10 0f 17 10 12 0f 07 08 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 40 3f 46 40 3c 3b 39 3c 4f 4f 54 56 63 61 68 6e 6f 72 6e 77 73 78 6f 65 65 52 52 4f 4e 43 40 41 39 35 38 3c 43 3f 43 33 34 3a 2d 30 31 3a 29 26 2a 1e 12 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 12 1a
 1f 2b 2d 32 34 34 40 44 47 50 49 53 51 5a 56 54 5c 5b 57 5c 62 58 5a 60 5d 62 6a 61 61 61 5b 58 5e 5d 5e 63 5c 5f 58 56 5f 5e 5e 62 5b 6d 65 71 7f 79 81 89 8a 81 7e 84 7a 82 7b 76 76 78 82 7e 85 77 79 6f 68 66 62 5c 58 4d 30 1a 0d 0d 15 12 15 0c 0d 0a 06 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 3c 49 4a 44 40 3b 46 4c 54 55 5a 60 68 6e 6c 78 6c 73 6b 65 62 66 68 5f 60 52 4c 53 42 3f 46 36 3f 3c 34 3e 35 35 3c 3a 35 3b 32 33 2f 32 2a 29 22 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 11 10 1e 2a 2b 38 36 36 3f 49 50 54 5a 59 65 60 5b 66 63 68 66 61 69 66 6a 67 70 68 6c 70 74 6f 68 68 6f 6b 65 67 69 6b 66 6d 62 66 62 65 6e 64 6b 77 77 79 84 79 84 8c 7f 84 83 82 81 76 80 7e 7e 7d 76 70 75 6b 64 67 62 59 4f 2c 16 10 0f 12 13 0d 10 06 06 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 31 43 3d 3a 42 45 48 50 54 43 5f 61 65 6e 68 70 6a 66 6f 6f 65 71 61 5e 54 4c 4d 46 44 41 3d 39 31 35 3b 3e 3d 31 32 30 39 35 30 2e 32 25 24 1b 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1b 1c 1f 2c 2f 34 3c 52 4e 59 66 63 64 65 68 6f 6b 71 72 6d 6b 74 73 72 6a 6d 71 70 72 71 6d 70 6f 6d 76 70 6f 6f 71 72 70 70 71 72 77 6d 75 73 76 7b 7d 84 86 88 88 8c 81 89 8d 83 82 85 79 76 74 7b 78 71 79 74 69 64 5d 33 17 10 1a 13 14 0d 11 0a 08 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 30 3f 3e 40 39 43 3b 47 4c 5e 5b 5f 67 65 6a 64 60 69 6a 63 62 5e 51 51 50 42 3d 44 3d 32 39 38 3b 34 38 3a 2e 37 3a 36 31 2c 2c 2d 26 20 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 0e 14 16 1f 28 33 37 46 54 61 69 63 6d 68 66 78 70 77 75 71 75 70 6b 77 75 78 73 71 6f 73 7b 7a 78 7c 74 79 73 73 7a 72 74 7c 77 7e 7b 78 7f 8a 8e 8f 93 92 92 91 99 91 99 9a 98 90 95 94 90 87 8a 8d 85 84 83 86 84 78 63 39 1c 15 17 11 13 12 14 10 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 28 38 2f 32 3d 39 41 4d 58 5c 59 5d 5d 63 5f 63 66 64 5e 5d 54 5f 51 44 3c 36 42 35 37 3b 3e 39 36 34 3f 33 38 39 2f 27 2e 2f 27 24 19 0f 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 12 17 26 2e 39 40 4c 51 60 62 6a 69 6e 68 6a 6e 73 6e 6a 7b 6e 75 70 70 6c 6a 76 72 72 77 6c 6e 76 6c 6f 74 73 73 6f 7b 78 7b 7c 82 88 86 90 94 90 9e 9f a5 9d a4 a5 a2 a8 9f a5 9d 98 99 92 92 89 8d 83 90 87 78 61 40 24 19 10 14 1b 1b 17 18 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 2d 39 2e 30 30 32 3d 47 45 51 55 51 54 5d 4a 58 5a 58 59 4c 51 52 4b 4a 43 37 40 38 3a 3c 39 38 39 40 37 27 3b 32 38 2b 22 26 26 12 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 17 1a 21 37 39 4f 53 5a 5e 66 70 69 68 64 6c 71 72 73 6b 6a 67 65 6c 6d 69 6c 69 6c 6e 70 6c 69 65 6e 6f 6c 70 75 74 7d 75 78 79 86 83 85 87 8b 92 9d a3 a4 9e 9f 9e 9e a4 9e a3 97 8f 88 89 86 7e 85 82 73 6d 42 20 1b 1e 1e 1d 1b 1d 11 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 25 35 30 39 2d 2b 37 39 35 45 47 4f 4d 53 51 4f 50 4b 44 44 45 49 4b 44 35 3e 2f 3a 36 34 42 3a 3f 31 35 30 2e 2a 2a 2a 29 21 0c 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 10 13 23 25 32 3e 49 4e 56 59 64 64 69 6a 6a 6c 6f 66 6a 67 65 6b 67 63 6a 65 6b 6a 65 6a 6e 65 67 6b 64 73 63 72 70 6b 6e 6c 76 7e 7f 82 82 86 8e 92 9b 9b 9a 9c 9d 96 a1 97 96 8c 84 8a 86 81 84 86 7d 80 69 3c 2c 24 23 26 23 1d 14 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 36 28 2a 34 32 31 32 37 39 41 3d 3a 44 42 4e 45 44 41 3e 45 3f 40 41 37 3b 39 3b 3a 40 43 41 3b 36 33 30 2d 25 2b 22 21 16 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0e 13 1c 2e 2f 37 44 46 5d 59 5a 64 5f 64 63 6d 6b 64 61 68 66 66 60 64 61 62 69 65 5e 65 67 64 65 67 64 63 69 60 68 6e 6c 6d 6f 72 78 7d 7b 85 84 89 96 9b 8f 90 96 96 89 8d 8e 8a 81 79 7d 7e 7d 81 73 6a 47 28 1e 29 23 1f 23 1c 12 0a 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 23 31 26 25 32 2d 31 38 30 37 2e 36 3a 40 43 43 42 37 3c 3e 3f 3d 36 3c 39 36 38 2f 37 39 40 37 38 35 36 34 2f 20 22 19 0d 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 16 1f 2f 33 45 50 4a 53 54 62 60 63 5e 55 61 63 68 60 56 62 5e 5f 5d 60 60 5c 58 62 5f 58 5f 60 64 62 68 68 5f 65 65 6e 68 6a 6e 6e 75 7e 80 7b 84 8d 91 86 8e 90 84 87 84 82 82 7a 7d 78 79 77 67 51 2e 21 1b 1e 24 23 18 15 07 09 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 29 29 32 2d 2d 22 2e 30 2e 31 31 3a 3b 37 41 3e 43 44 44 45 44 39 39 36 35 30 39 35 37 3a 34 39 33 30 22 19 19 15 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 07 13 1a 22 2d 36 3b 42 47 50 59 55 57 5a 5b 5e 65 5e 5d 59 51 5d 5a 5e 61 5a 5b 5d 5d 5c 5a 64 52 5b 5e 5d 5b 5a 59 60 6a 68 6f 68 70 71 72 7c 78 7a 86 84 84 8a 85 88 85 86 82 7a 81 78 7d 7e 79 73 5a 36 28 21 29 25 21 1a 1e 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 10 34 2d 33 2f 2e 2e 2b 35 2f 35 34 39 42 46 47 45 44 4a 4a 3d 43 3c 38 34 37 33 37 35 36 38 2e 2c 21 1e 1e 16 14 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 08 10 17 21 2a 35 36 4a 44 4d 4e 55 58 59 5b 57 5f 56 5b 5a 5a 5b 58 55 5c 5e 4f 5b 58 52 51 5c 5b 5f 58 64 59 5f 5d 5f 69 68 63 70 67 71 76 75 7b 7f 82 7d 7e 88 7a 85 83 86 7f 84 85 7b 71 74 5b 3a 2d 2f 22 29 1d 23 13 11 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 29 2b 2c 31 29 2c 30 2c 33 31 39 40 44 43 44 45 4d 4b 40 39 36 35 3e 35 31 2f 30 31 3a 2d 25 21 1f 1e 16 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 13 26 23 2a 39 3f 49 49 54 52 4d 5c 5a 5a 54 55 57 4f 58 53 5e 51 54 5c 4e 4e 54 4f 54 57 57 5b 5b 58 5c 5c 5d 5f 5e 66 60 68 67 6a 6a 7a 7c 77 7d 7b 7d 7d 7b 84 84 87 81 82 7f 79 7b 5c 41 2c 1f 22 1d 1c 19 0b 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 2f 2b 30 2b 2c 34 33 2f 31 30 36 36 37 3d 3a 3f 44 3e 40 36 36 37 33 34 2b 2f 30 25 2c 27 1f 17 11 0e 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 11 1e 23 29 33 3e 3d 45 43 49 51 55 50 4d 4d 52 50 55 4b 4d 53 59 4d 51 54 52 59 50 54 52 50 58 55 5a 60 58 62 5e 5a 5f 64 69 67 64 73 78 81 78 79 7b 7a 82 80 84 82 8b 82 8c 83 74 5c 3a 2a 2d 2b 24 1e 12 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 2d 24 2d 33 30 2a 30 2a 30 2f 36 39 3f 35 3f 39 38 41 3f 2e 35 2c 36 2e 30 2c 27 26 27 21 1c 14 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 16 15 1e 27 2b 31 37 41 42 4f 47 4c 45 48 4e 4b 51 53 53 52 4d 51 52 51 49 50 4e 51 52 54 55 51 51 59 5a 55 5a 62 5a 62 5c 67 66 6a 76 77 7c 76 79 7e 7f 7d 84 88 8b 8f 89 80 72 64 36 2d 23 23 1e 23 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 2d 28 27 28 2b 2d 29 38 34 27 2f 3a 34 38 3d 3d 44 41 34 34 36 33 2e 30 25 29 2e 1a 1a 13 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 12 22 29 2a 35 39 3d 47 3a 41 44 3f 42 48 48 49 48 4a 4f 4e 47 50 4c 46 43 4f 4b 50 54 55 52 50 4e 57 5a 63 5a 59 65 5f 62 64 71 74 77 7a 7b 7a 7d 87 89 81 8d 84 7e 7e 63 35 28 1e 1c 1c 0d 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 2d 27 2c 29 29 2c 30 32 34 2d 2a 32 39 3b 3f 37 40 3b 35 2f 30 31 30 25 1f 1c 20 19 13 0a 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 14 10 1d 24 24 2b 36 34 31 32 33 3f 46 43 43 42 42 47 4f 51 47 44 49 49 49 53 4e 4f 40 4c 54 54 59 60 54 5e 58 59 61 63 5e 62 68 6e 75 7a 7c 7e 82 8f 81 85 91 83 7c 74 62 36 22 19 16 1a 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 32 30 2f 36 2f 2f 29 30 29 35 35 36 37 41 3a 35 38 3e 3b 2d 2c 25 2d 24 1b 19 1b 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0a 15 15 23 28 26 29 2e 38 39 3a 39 39 45 42 47 41 4d 49 48 52 4b 4e 49 4a 53 52 4c 57 4f 50 55 54 54 5a 58 59 61 68 6c 6c 70 73 6c 7a 7b 83 85 8a 87 93 93 82 84 6e 37 22 15 10 12 0b 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 2e 2e 2e 34 36 2b 3a 30 36 36 34 39 40 3e 41 41 39 34 2f 30 2c 21 1d 19 1b 11 0c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0b 0b 17 26 23 2a 26 2b 2c 33 32 3a 3c 35 2d 46 3c 45 44 42 48 49 4f 4a 50 47 4d 4e 50 58 51 58 5a 4f 58 56 58 64 67 68 63 68 75 79 87 84 8b 82 8e 90 7f 82 71 34 15 14 0a 0a 0e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 30 24 3e 39 2c 30 2f 31 3d 43 3d 3c 3f 3f 3c 37 37 37 2a 25 28 1a 1b 19 09 0b 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 0d 15 1f 20 26 25 2b 2c 34 39 3c 37 31 36 3d 40 4b 40 3d 43 41 4d 4c 4b 49 50 4c 52 55 55 4d 57 5d 64 69 62 62 6b 6a 6f 77 7c 7d 7c 86 89 84 85 76 66 3d 1f 1a 08 09 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 32 2f 27 30 2a 2c 34 30 36 43 36 36 3c 30 38 35 28 24 18 1a 0d 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0c 11 0f 10 19 1c 2a 29 2a 30 32 33 32 39 38 3d 35 41 41 41 48 4a 45 46 46 4a 4b 50 53 53 48 56 59 63 64 5e 65 62 6b 6d 73 75 79 80 86 88 7f 81 79 72 3b 23 14 11 0c 0b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 21 2a 2f 2c 28 2c 2e 2f 33 35 31 39 34 33 1f 2a 23 1f 1f 1b 0f 14 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0a 11 17 21 24 2c 29 22 2a 2d 34 3b 35 34 3e 3c 37 3e 41 47 4a 46 48 4c 4e 55 51 53 53 5e 5b 58 67 61 60 6c 68 6b 74 6d 7d 7b 82 7b 85 73 3d 1e 10 10 09 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 22 27 29 1e 25 2c 25 2b 2a 29 25 27 27 21 1e 19 0c 0f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 14 11 15 19 24 25 26 23 26 2e 2e 2b 34 36 3e 32 3c 36 3d 3b 3a 44 49 49 4c 52 53 50 57 5b 62 5a 66 5d 60 68 6b 73 70 6d 7a 6f 73 67 3d 13 19 0d 0f 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 18 22 1f 11 20 21 1b 27 22 19 1b 19 19 10 12 17 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 06 13 14 12 13 1f 25 24 25 2b 29 26 30 2f 39 36 32 31 35 3d 41 44 42 4d 44 53 51 4b 56 56 60 58 5e 5d 64 67 61 6b 67 67 61 5b 3e 1c 1a 09 0a 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 19 1b 1b 1c 18 15 1d 1e 23 15 1c 0b 0d 0d 0b 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 07 0b 11 13 0e 16 14 1d 20 22 22 1b 21 2c 29 24 2d 2e 3a 39 3d 44 45 37 44 44 49 4f 48 4c 4c 55 53 4e 5a 4d 53 53 50 4e 33 18 0e 12 0d 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0f 0e 09 05 0b 0a 16 0b 07 0a 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0b 0d 10 0a 0f 09 16 12 12 16 1e 27 2e 32 2c 30 29 2c 32 29 37 3b 3e 39 35 38 3d 38 3a 40 3c 3c 34 37 27 0e 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 03 06 05 03 00 06 06 09 09 09 15 21 1d 24 25 1c 24 1e 21 22 28 2f 2a 24 23 23 22 28 29 28 2d 2c 22 25 1a 0f 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 12 16 15 0e 0f 0f 0d 09 16 10 0e 19 14 15 14 19 13 19 1e 15 11 0f 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 09 00 0f 05 07 09 10 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
