 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 04 04 04 03 03 03 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 04 04 04 05 05 05 06 06 06 09 09 09 07 07 07 05 05 05 06 06 06 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 06 06 06 0b 0b 0b 0a 0a 0a 11 11 11 13 13 13 1b 1b 1b 15 15 15 0e 0e 0e 0c 0c 0c 06 06 06 05 05 05 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 02 02 02 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 05 05 05 07 07 07 09 09 09 0e 0e 0e 17 17 17 1a 1a 1a 21 21 21 25 25 25 24 24 24 27 27 27 21 21 21 14 14 14 0d 0d 0d 0e 0e 0e 0d 0d 0d 07 07 07 06 06 06 06 06 06 04 04 04 04 04 04 03 03 03 04 04 04 03 03 03 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 09 09 09 0b 0b 0b 0e 0e 0e 1c 1c 1c 21 21 21 42 42 42 4c 4c 4c 60 60 60 68 68 68 b1 b1 b1 ba ba ba 59 59 59 47 47 47 35 35 35 2f 2f 2f 2b 2b 2b 1e 1e 1e 11 11 11 0f 0f 0f 14 14 14 08 08 08 09 09 09 09 09 09 05 05 05 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 03 03 03 04 04 04 06 06 06 07 07 07 0c 0c 0c 18 18 18 20 20 20 2a 2a 2a 4b 4b 4b 56 56 56 8f 8f 8f cd cd cd e7 e7 e7 e5 e5 e5 f8 f8 f8 f0 f0 f0 d6 d6 d6 b7 b7 b7 94 94 94 6f 6f 6f 6d 6d 6d 62 62 62 40 40 40 29 29 29 25 25 25 17 17 17 13 13 13 11 11 11 10 10 10 09 09 09 09 09 09 04 04 04 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 08 08 08 0f 0f 0f 14 14 14 1f 1f 1f 37 37 37 5d 5d 5d bd bd bd c9 c9 c9 e3 e3 e3 fa fa fa fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 d5 d5 d5 c0 c0 c0 ba ba ba af af af 8f 8f 8f 6b 6b 6b 5b 5b 5b 49 49 49 37 37 37 26 26 26 18 18 18 0f 0f 0f 08 08 08 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 09 09 09 13 13 13 24 24 24 41 41 41 5d 5d 5d 82 82 82 a2 a2 a2 cd cd cd f6 f6 f6 ff ff ff ff ff ff fe fe fe fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f9 f9 df df df d8 d8 d8 d5 d5 d5 e8 e8 e8 ed ed ed db db db c3 c3 c3 a6 a6 a6 93 93 93 84 84 84 65 65 65 48 48 48 2f 2f 2f 13 13 13 0a 0a 0a 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 0a 0a 0a 17 17 17 37 37 37 63 63 63 96 96 96 c4 c4 c4 d2 d2 d2 e6 e6 e6 f7 f7 f7 fa fa fa fe fe fe ff ff ff ff ff ff fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f5 f5 f5 ea ea ea e4 e4 e4 f5 f5 f5 f6 f6 f6 db db db c9 c9 c9 c2 c2 c2 b3 b3 b3 a7 a7 a7 9c 9c 9c a9 a9 a9 94 94 94 47 47 47 2e 2e 2e 17 17 17 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 08 08 08 1f 1f 1f 48 48 48 79 79 79 8a 8a 8a c3 c3 c3 c7 c7 c7 e8 e8 e8 fc fc fc fe fe fe fa fa fa fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe fe fe fe ff ff ff fe fe fe fd fd fd fa fa fa f9 f9 f9 df df df bf bf bf 96 96 96 95 95 95 9f 9f 9f 70 70 70 5c 5c 5c 42 42 42 23 23 23 0a 0a 0a 05 05 05 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 09 09 09 2b 2b 2b 82 82 82 f3 f3 f3 f6 f6 f6 e4 e4 e4 d9 d9 d9 ec ec ec fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd e7 e7 e7 b8 b8 b8 9a 9a 9a 8b 8b 8b 9a 9a 9a 9a 9a 9a 78 78 78 66 66 66 44 44 44 16 16 16 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0a 0a 0a 39 39 39 75 75 75 b4 b4 b4 d9 d9 d9 cb cb cb d3 d3 d3 dd dd dd f6 f6 f6 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 d3 d3 d3 b9 b9 b9 c0 c0 c0 dc dc dc d7 d7 d7 a2 a2 a2 86 86 86 88 88 88 49 49 49 14 14 14 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 08 08 08 2e 2e 2e 6e 6e 6e 90 90 90 b9 b9 b9 c0 c0 c0 cd cd cd d9 d9 d9 f6 f6 f6 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 da da da d0 d0 d0 ee ee ee fe fe fe f5 f5 f5 b3 b3 b3 87 87 87 8b 8b 8b 8f 8f 8f 4b 4b 4b 0b 0b 0b 03 03 03 02 02 02 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 1c 1c 1c 50 50 50 6e 6e 6e 9f 9f 9f ba ba ba cf cf cf e4 e4 e4 e7 e7 e7 f7 f7 f7 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f0 f0 f0 e0 e0 e0 ea ea ea fd fd fd ff ff ff e8 e8 e8 ae ae ae 8b 8b 8b 83 83 83 9b 9b 9b 9f 9f 9f 2a 2a 2a 04 04 04 03 03 03 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 09 09 09 3d 3d 3d 64 64 64 64 64 64 b0 b0 b0 c7 c7 c7 e6 e6 e6 f3 f3 f3 f1 f1 f1 f3 f3 f3 f9 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f0 f0 f0 e4 e4 e4 f6 f6 f6 ff ff ff fe fe fe e3 e3 e3 ae ae ae 9d 9d 9d 94 94 94 93 93 93 c1 c1 c1 47 47 47 04 04 04 03 03 03 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 18 18 18 5e 5e 5e 63 63 63 6f 6f 6f be be be e2 e2 e2 ed ed ed fb fb fb f6 f6 f6 ed ed ed fa fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f3 f3 f3 e7 e7 e7 ee ee ee fe fe fe fc fc fc d3 d3 d3 b2 b2 b2 ac ac ac a2 a2 a2 99 99 99 b6 b6 b6 72 72 72 0a 0a 0a 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 46 46 46 7b 7b 7b 73 73 73 8a 8a 8a d6 d6 d6 eb eb eb f1 f1 f1 fe fe fe fb fb fb f3 f3 f3 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fa fa fa ee ee ee e5 e5 e5 e5 e5 e5 e4 e4 e4 df df df be be be b1 b1 b1 a6 a6 a6 99 99 99 94 94 94 98 98 98 90 90 90 0c 0c 0c 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0d 0d 0d 6a 6a 6a a2 a2 a2 8a 8a 8a b4 b4 b4 f3 f3 f3 f2 f2 f2 fa fa fa fb fb fb fd fd fd fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fb fb fb ee ee ee e4 e4 e4 df df df dd dd dd d6 d6 d6 df df df c1 c1 c1 aa aa aa a3 a3 a3 99 99 99 8f 8f 8f 92 92 92 83 83 83 0a 0a 0a 03 03 03 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 79 79 79 b3 b3 b3 ac ac ac da da da f6 f6 f6 e4 e4 e4 f1 f1 f1 f7 f7 f7 fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f5 f5 f5 e6 e6 e6 d8 d8 d8 d0 d0 d0 d4 d4 d4 d2 d2 d2 cc cc cc c5 c5 c5 b6 b6 b6 9f 9f 9f 99 99 99 90 90 90 82 82 82 7f 7f 7f 69 69 69 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0e 0e 0e 6a 6a 6a c0 c0 c0 be be be d7 d7 d7 d7 d7 d7 d3 d3 d3 df df df eb eb eb f7 f7 f7 fd fd fd fb fb fb fc fc fc fc fc fc fe fe fe fe fe fe fe fe fe fe fe fe fe fe fe fa fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd eb eb eb d9 d9 d9 cb cb cb c3 c3 c3 c2 c2 c2 c2 c2 c2 c3 c3 c3 bb bb bb b4 b4 b4 ab ab ab 9b 9b 9b 98 98 98 8b 8b 8b 80 80 80 78 78 78 47 47 47 04 04 04 03 03 03 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0d 0d 0d 5e 5e 5e b6 b6 b6 b8 b8 b8 d2 d2 d2 dd dd dd c9 c9 c9 cf cf cf d8 d8 d8 e1 e1 e1 e3 e3 e3 e7 e7 e7 f2 f2 f2 f7 f7 f7 fa fa fa f6 f6 f6 f4 f4 f4 f3 f3 f3 e2 e2 e2 d8 d8 d8 fe fe fe fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f0 f0 f0 db db db ce ce ce c2 c2 c2 bc bc bc bf bf bf be be be b8 b8 b8 b3 b3 b3 b7 b7 b7 a6 a6 a6 9e 9e 9e 8e 8e 8e 89 89 89 7c 7c 7c 6e 6e 6e 35 35 35 06 06 06 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 65 65 65 b5 b5 b5 ae ae ae be be be b0 b0 b0 b6 b6 b6 bf bf bf c8 c8 c8 cb cb cb d1 d1 d1 db db db e6 e6 e6 eb eb eb e8 e8 e8 e6 e6 e6 e5 e5 e5 e0 e0 e0 c9 c9 c9 bd bd bd df df df b3 b3 b3 d3 d3 d3 e7 e7 e7 f4 f4 f4 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fa fa ee ee ee de de de ce ce ce c5 c5 c5 bd bd bd b9 b9 b9 b5 b5 b5 b4 b4 b4 ab ab ab a6 a6 a6 a0 a0 a0 98 98 98 8d 8d 8d 87 87 87 80 80 80 77 77 77 71 71 71 49 49 49 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 20 20 20 77 77 77 b7 b7 b7 a4 a4 a4 a8 a8 a8 86 86 86 96 96 96 a6 a6 a6 b1 b1 b1 bc bc bc c7 c7 c7 d3 d3 d3 da da da d7 d7 d7 dc dc dc dc dc dc df df df d9 d9 d9 bd bd bd ac ac ac 93 93 93 48 48 48 46 46 46 52 52 52 66 66 66 87 87 87 c2 c2 c2 fd fd fd ea ea ea f0 f0 f0 ef ef ef df df df cc cc cc c1 c1 c1 bc bc bc b6 b6 b6 b5 b5 b5 b1 b1 b1 a6 a6 a6 a2 a2 a2 99 99 99 99 99 99 8e 8e 8e 85 85 85 80 80 80 7c 7c 7c 78 78 78 74 74 74 77 77 77 5d 5d 5d 16 16 16 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 07 07 07 2f 2f 2f 83 83 83 a9 a9 a9 8e 8e 8e 81 81 81 7a 7a 7a 88 88 88 93 93 93 9d 9d 9d b1 b1 b1 c5 c5 c5 ce ce ce d2 d2 d2 cf cf cf d6 d6 d6 d6 d6 d6 da da da d1 d1 d1 b5 b5 b5 a6 a6 a6 72 72 72 23 23 23 1f 1f 1f 21 21 21 2a 2a 2a 37 37 37 5a 5a 5a cb cb cb c3 c3 c3 cc cc cc cd cd cd c4 c4 c4 b4 b4 b4 a8 a8 a8 a8 a8 a8 aa aa aa a9 a9 a9 a9 a9 a9 9e 9e 9e 90 90 90 8b 8b 8b 8a 8a 8a 7f 7f 7f 7c 7c 7c 7b 7b 7b 7a 7a 7a 76 76 76 75 75 75 68 68 68 6a 6a 6a 2a 2a 2a 05 05 05 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0a 0a 0a 3c 3c 3c 91 91 91 83 83 83 70 70 70 76 76 76 78 78 78 87 87 87 98 98 98 a4 a4 a4 b0 b0 b0 c1 c1 c1 cb cb cb c8 c8 c8 cf cf cf d1 d1 d1 d1 d1 d1 d3 d3 d3 ca ca ca b2 b2 b2 9e 9e 9e 5e 5e 5e 10 10 10 0f 0f 0f 11 11 11 14 14 14 1d 1d 1d 3f 3f 3f 9e 9e 9e aa aa aa b3 b3 b3 b3 b3 b3 aa aa aa a2 a2 a2 96 96 96 92 92 92 a1 a1 a1 9e 9e 9e 9d 9d 9d 95 95 95 8d 8d 8d 84 84 84 7f 7f 7f 7f 7f 7f 7e 7e 7e 7c 7c 7c 7a 7a 7a 74 74 74 68 68 68 5c 5c 5c 69 69 69 3d 3d 3d 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0b 0b 0b 45 45 45 92 92 92 7d 7d 7d 76 76 76 74 74 74 78 78 78 8b 8b 8b 9c 9c 9c a6 a6 a6 ae ae ae b8 b8 b8 b5 b5 b5 be be be c6 c6 c6 cb cb cb ca ca ca cb cb cb c6 c6 c6 ae ae ae 98 98 98 5d 5d 5d 09 09 09 08 08 08 07 07 07 08 08 08 13 13 13 2e 2e 2e 90 90 90 9c 9c 9c 9e 9e 9e 9b 9b 9b 93 93 93 91 91 91 8c 8c 8c 8b 8b 8b 96 96 96 92 92 92 8f 8f 8f 8a 8a 8a 85 85 85 7f 7f 7f 7a 7a 7a 7d 7d 7d 7a 7a 7a 76 76 76 73 73 73 69 69 69 5d 5d 5d 54 54 54 60 60 60 4b 4b 4b 09 09 09 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0f 0f 0f 4c 4c 4c 95 95 95 7a 7a 7a 73 73 73 78 78 78 7d 7d 7d 8c 8c 8c 95 95 95 9d 9d 9d a1 a1 a1 a1 a1 a1 a8 a8 a8 b2 b2 b2 b9 b9 b9 bd bd bd bd bd bd c3 c3 c3 bc bc bc ab ab ab 96 96 96 64 64 64 06 06 06 06 06 06 05 05 05 05 05 05 0b 0b 0b 1c 1c 1c 85 85 85 91 91 91 94 94 94 8f 8f 8f 8c 8c 8c 8d 8d 8d 8b 8b 8b 90 90 90 93 93 93 98 98 98 8e 8e 8e 84 84 84 7f 7f 7f 78 78 78 72 72 72 75 75 75 76 76 76 6c 6c 6c 67 67 67 62 62 62 5c 5c 5c 56 56 56 5a 5a 5a 53 53 53 0d 0d 0d 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 10 10 10 51 51 51 91 91 91 80 80 80 69 69 69 74 74 74 78 78 78 81 81 81 8c 8c 8c 96 96 96 94 94 94 96 96 96 9c 9c 9c a6 a6 a6 a9 a9 a9 ab ab ab ab ab ab b1 b1 b1 ad ad ad a3 a3 a3 93 93 93 6a 6a 6a 05 05 05 04 04 04 04 04 04 03 03 03 06 06 06 13 13 13 7c 7c 7c 8e 8e 8e 92 92 92 8e 8e 8e 91 91 91 95 95 95 92 92 92 93 93 93 9d 9d 9d 95 95 95 87 87 87 7b 7b 7b 73 73 73 6f 6f 6f 6a 6a 6a 6a 6a 6a 69 69 69 61 61 61 5f 5f 5f 5b 5b 5b 59 59 59 56 56 56 58 58 58 54 54 54 0d 0d 0d 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 10 10 10 50 50 50 88 88 88 74 74 74 60 60 60 68 68 68 72 72 72 7e 7e 7e 8a 8a 8a 93 93 93 8e 8e 8e 8f 8f 8f 98 98 98 9d 9d 9d 9f 9f 9f 9e 9e 9e 9a 9a 9a 9c 9c 9c 9c 9c 9c 95 95 95 8b 8b 8b 6a 6a 6a 05 05 05 04 04 04 03 03 03 03 03 03 05 05 05 0d 0d 0d 6e 6e 6e 88 88 88 90 90 90 90 90 90 8c 8c 8c 8f 8f 8f 91 91 91 98 98 98 98 98 98 84 84 84 75 75 75 6d 6d 6d 69 69 69 67 67 67 64 64 64 61 61 61 60 60 60 5d 5d 5d 5a 5a 5a 58 58 58 59 59 59 53 53 53 53 53 53 57 57 57 12 12 12 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0c 0c 0c 4f 4f 4f 81 81 81 64 64 64 5e 5e 5e 61 61 61 6a 6a 6a 7d 7d 7d 86 86 86 83 83 83 83 83 83 8b 8b 8b 94 94 94 97 97 97 98 98 98 93 93 93 8f 8f 8f 8c 8c 8c 8a 8a 8a 88 88 88 83 83 83 6a 6a 6a 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 63 63 63 85 85 85 8c 8c 8c 90 90 90 90 90 90 94 94 94 90 90 90 94 94 94 8e 8e 8e 79 79 79 6c 6c 6c 65 65 65 5e 5e 5e 60 60 60 5f 5f 5f 5f 5f 5f 5d 5d 5d 5b 5b 5b 57 57 57 55 55 55 59 59 59 56 56 56 52 52 52 54 54 54 10 10 10 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 07 07 07 45 45 45 7a 7a 7a 57 57 57 5d 5d 5d 5c 5c 5c 60 60 60 6b 6b 6b 75 75 75 76 76 76 77 77 77 82 82 82 8c 8c 8c 92 92 92 92 92 92 8d 8d 8d 86 86 86 82 82 82 7e 7e 7e 7b 7b 7b 75 75 75 66 66 66 09 09 09 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 59 59 59 86 86 86 88 88 88 8b 8b 8b 8e 8e 8e 8e 8e 8e 87 87 87 86 86 86 7a 7a 7a 6b 6b 6b 63 63 63 5d 5d 5d 5a 5a 5a 5a 5a 5a 59 59 59 58 58 58 5a 5a 5a 56 56 56 53 53 53 57 57 57 58 58 58 52 52 52 50 50 50 4c 4c 4c 0a 0a 0a 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 2e 2e 2e 78 78 78 58 58 58 5c 5c 5c 56 56 56 56 56 56 5e 5e 5e 65 65 65 65 65 65 6b 6b 6b 75 75 75 7d 7d 7d 85 85 85 88 88 88 8a 8a 8a 84 84 84 7e 7e 7e 78 78 78 71 71 71 6d 6d 6d 63 63 63 0b 0b 0b 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 4c 4c 4c 86 86 86 82 82 82 85 85 85 8c 8c 8c 8a 8a 8a 7d 7d 7d 73 73 73 6b 6b 6b 66 66 66 60 60 60 5a 5a 5a 58 58 58 55 55 55 54 54 54 55 55 55 54 54 54 54 54 54 51 51 51 57 57 57 52 52 52 52 52 52 4d 4d 4d 32 32 32 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 15 15 15 6a 6a 6a 61 61 61 5a 5a 5a 53 53 53 54 54 54 55 55 55 59 59 59 58 58 58 5d 5d 5d 69 69 69 71 71 71 75 75 75 76 76 76 7f 7f 7f 85 85 85 81 81 81 76 76 76 6f 6f 6f 6e 6e 6e 67 67 67 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 43 43 43 82 82 82 7d 7d 7d 7e 7e 7e 86 86 86 88 88 88 75 75 75 6c 6c 6c 68 68 68 64 64 64 60 60 60 5d 5d 5d 5a 5a 5a 54 54 54 50 50 50 50 50 50 51 51 51 51 51 51 51 51 51 54 54 54 54 54 54 57 57 57 4c 4c 4c 18 18 18 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 41 41 41 5e 5e 5e 54 54 54 50 50 50 4d 4d 4d 50 50 50 52 52 52 52 52 52 52 52 52 5a 5a 5a 64 64 64 6a 6a 6a 6c 6c 6c 74 74 74 81 81 81 82 82 82 73 73 73 6a 6a 6a 6a 6a 6a 68 68 68 10 10 10 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 3c 3c 3c 82 82 82 7c 7c 7c 81 81 81 7a 7a 7a 7d 7d 7d 6d 6d 6d 61 61 61 5f 5f 5f 5d 5d 5d 5d 5d 5d 5b 5b 5b 58 58 58 53 53 53 4f 4f 4f 4e 4e 4e 4f 4f 4f 50 50 50 54 54 54 54 54 54 56 56 56 57 57 57 46 46 46 0c 0c 0c 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 26 26 26 47 47 47 4a 4a 4a 47 47 47 45 45 45 44 44 44 45 45 45 4d 4d 4d 50 50 50 51 51 51 58 58 58 60 60 60 65 65 65 68 68 68 70 70 70 75 75 75 70 70 70 68 68 68 68 68 68 68 68 68 17 17 17 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 31 31 31 80 80 80 78 78 78 7d 7d 7d 78 78 78 72 72 72 69 69 69 60 60 60 5a 5a 5a 5a 5a 5a 56 56 56 52 52 52 4f 4f 4f 51 51 51 50 50 50 52 52 52 53 53 53 52 52 52 55 55 55 55 55 55 59 59 59 57 57 57 3a 3a 3a 06 06 06 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 1f 1f 1f 41 41 41 43 43 43 42 42 42 3f 3f 3f 43 43 43 42 42 42 43 43 43 49 49 49 4e 4e 4e 4e 4e 4e 55 55 55 5b 5b 5b 5a 5a 5a 5d 5d 5d 62 62 62 65 65 65 69 69 69 61 61 61 64 64 64 1b 1b 1b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 26 26 26 77 77 77 71 71 71 6e 6e 6e 72 72 72 67 67 67 63 63 63 5c 5c 5c 57 57 57 53 53 53 50 50 50 50 50 50 52 52 52 53 53 53 4f 4f 4f 4f 4f 4f 51 51 51 4f 4f 4f 50 50 50 56 56 56 59 59 59 56 56 56 29 29 29 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 19 19 19 3d 3d 3d 44 44 44 42 42 42 3e 3e 3e 41 41 41 41 41 41 42 42 42 45 45 45 48 48 48 4b 4b 4b 4b 4b 4b 4f 4f 4f 54 54 54 53 53 53 54 54 54 54 54 54 5c 5c 5c 61 61 61 5a 5a 5a 1c 1c 1c 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 1e 1e 1e 72 72 72 6a 6a 6a 65 65 65 64 64 64 5b 5b 5b 57 57 57 57 57 57 56 56 56 50 50 50 4e 4e 4e 4e 4e 4e 52 52 52 4f 4f 4f 4d 4d 4d 57 57 57 53 53 53 53 53 53 52 52 52 54 54 54 58 58 58 55 55 55 19 19 19 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 36 36 36 44 44 44 45 45 45 42 42 42 43 43 43 42 42 42 43 43 43 43 43 43 46 46 46 47 47 47 4a 4a 4a 4a 4a 4a 4c 4c 4c 4e 4e 4e 4c 4c 4c 4b 4b 4b 50 50 50 54 54 54 57 57 57 1f 1f 1f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 15 15 15 68 68 68 65 65 65 65 65 65 5e 5e 5e 57 57 57 53 53 53 52 52 52 54 54 54 4e 4e 4e 4d 4d 4d 4d 4d 4d 4b 4b 4b 4c 4c 4c 4d 4d 4d 51 51 51 50 50 50 52 52 52 54 54 54 5c 5c 5c 64 64 64 45 45 45 08 08 08 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 2e 2e 2e 41 41 41 41 41 41 44 44 44 42 42 42 40 40 40 40 40 40 43 43 43 46 46 46 48 48 48 48 48 48 48 48 48 48 48 48 47 47 47 4a 4a 4a 47 47 47 47 47 47 4a 4a 4a 4b 4b 4b 1e 1e 1e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 10 10 10 63 63 63 5e 5e 5e 61 61 61 61 61 61 58 58 58 50 50 50 50 50 50 4d 4d 4d 4b 4b 4b 4e 4e 4e 4a 4a 4a 49 49 49 4e 4e 4e 4d 4d 4d 4b 4b 4b 4d 4d 4d 50 50 50 58 58 58 58 58 58 5b 5b 5b 27 27 27 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 20 20 20 41 41 41 3e 3e 3e 3d 3d 3d 41 41 41 41 41 41 3f 3f 3f 40 40 40 44 44 44 46 46 46 49 49 49 49 49 49 46 46 46 46 46 46 47 47 47 49 49 49 46 46 46 48 48 48 45 45 45 1e 1e 1e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 0a 0a 0a 62 62 62 5b 5b 5b 5a 5a 5a 5d 5d 5d 5a 5a 5a 54 54 54 52 52 52 4c 4c 4c 4d 4d 4d 4d 4d 4d 4f 4f 4f 4d 4d 4d 53 53 53 4e 4e 4e 4d 4d 4d 4e 4e 4e 57 57 57 60 60 60 4e 4e 4e 3c 3c 3c 0b 0b 0b 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 14 14 14 38 38 38 3e 3e 3e 3b 3b 3b 42 42 42 42 42 42 3f 3f 3f 40 40 40 43 43 43 45 45 45 46 46 46 48 48 48 46 46 46 42 42 42 42 42 42 46 46 46 46 46 46 48 48 48 47 47 47 23 23 23 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 08 08 08 59 59 59 58 58 58 55 55 55 58 58 58 5a 5a 5a 57 57 57 53 53 53 4c 4c 4c 50 50 50 59 59 59 55 55 55 47 47 47 46 46 46 49 49 49 4a 4a 4a 4a 4a 4a 5a 5a 5a 52 52 52 48 48 48 20 20 20 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 31 31 31 44 44 44 3a 3a 3a 3c 3c 3c 3b 3b 3b 3e 3e 3e 41 41 41 42 42 42 41 41 41 42 42 42 46 46 46 4a 4a 4a 42 42 42 40 40 40 40 40 40 43 43 43 42 42 42 43 43 43 24 24 24 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 06 06 06 4d 4d 4d 54 54 54 54 54 54 59 59 59 58 58 58 53 53 53 4e 4e 4e 4d 4d 4d 52 52 52 4f 4f 4f 44 44 44 44 44 44 48 48 48 47 47 47 48 48 48 49 49 49 4f 4f 4f 48 48 48 3d 3d 3d 0b 0b 0b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 25 25 25 3e 3e 3e 3c 3c 3c 3b 3b 3b 38 38 38 3a 3a 3a 3c 3c 3c 3e 3e 3e 41 41 41 3f 3f 3f 40 40 40 47 47 47 42 42 42 3f 3f 3f 3d 3d 3d 3e 3e 3e 3c 3c 3c 3b 3b 3b 23 23 23 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 41 41 41 4e 4e 4e 50 50 50 57 57 57 52 52 52 4e 4e 4e 4b 4b 4b 4e 4e 4e 51 51 51 43 43 43 45 45 45 46 46 46 45 45 45 44 44 44 45 45 45 47 47 47 49 49 49 45 45 45 26 26 26 04 04 04 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 18 18 18 36 36 36 3b 3b 3b 3b 3b 3b 37 37 37 38 38 38 37 37 37 3a 3a 3a 3c 3c 3c 40 40 40 3e 3e 3e 40 40 40 43 43 43 46 46 46 3d 3d 3d 3c 3c 3c 37 37 37 36 36 36 23 23 23 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 3d 3d 3d 4d 4d 4d 4d 4d 4d 51 51 51 52 52 52 55 55 55 4b 4b 4b 4e 4e 4e 48 48 48 43 43 43 43 43 43 45 45 45 44 44 44 42 42 42 40 40 40 44 44 44 44 44 44 39 39 39 0d 0d 0d 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 35 35 35 3d 3d 3d 3d 3d 3d 38 38 38 37 37 37 38 38 38 3a 3a 3a 39 39 39 38 38 38 37 37 37 3a 3a 3a 3d 3d 3d 48 48 48 39 39 39 35 35 35 35 35 35 35 35 35 24 24 24 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 35 35 35 4a 4a 4a 4a 4a 4a 4f 4f 4f 54 54 54 58 58 58 50 50 50 4d 4d 4d 4a 4a 4a 47 47 47 41 41 41 41 41 41 44 44 44 47 47 47 4c 4c 4c 4f 4f 4f 41 41 41 22 22 22 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 25 25 25 46 46 46 39 39 39 36 36 36 37 37 37 39 39 39 3a 3a 3a 37 37 37 35 35 35 33 33 33 35 35 35 35 35 35 37 37 37 35 35 35 33 33 33 33 33 33 34 34 34 26 26 26 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 2b 2b 2b 42 42 42 45 45 45 4a 4a 4a 49 49 49 4a 4a 4a 4f 4f 4f 53 53 53 4d 4d 4d 4b 4b 4b 4c 4c 4c 57 57 57 65 65 65 6d 6d 6d 6d 6d 6d 66 66 66 3c 3c 3c 0c 0c 0c 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 3b 3b 3b 36 36 36 35 35 35 36 36 36 35 35 35 37 37 37 35 35 35 37 37 37 32 32 32 32 32 32 31 31 31 31 31 31 31 31 31 31 31 31 33 33 33 36 36 36 2d 2d 2d 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 24 24 24 39 39 39 39 39 39 3a 3a 3a 3e 3e 3e 3d 3d 3d 41 41 41 51 51 51 65 65 65 70 70 70 76 76 76 75 75 75 73 73 73 6c 6c 6c 67 67 67 5e 5e 5e 23 23 23 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 35 35 35 35 35 35 37 37 37 33 33 33 33 33 33 33 33 33 32 32 32 2f 2f 2f 2f 2f 2f 2e 2e 2e 2e 2e 2e 2d 2d 2d 2e 2e 2e 2d 2d 2d 2d 2d 2d 29 29 29 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 1b 1b 1b 33 33 33 34 34 34 36 36 36 3a 3a 3a 4b 4b 4b 69 69 69 7b 7b 7b 7e 7e 7e 79 79 79 72 72 72 6a 6a 6a 62 62 62 5d 5d 5d 5c 5c 5c 39 39 39 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 22 22 22 34 34 34 3a 3a 3a 36 36 36 34 34 34 33 33 33 31 31 31 2e 2e 2e 2f 2f 2f 2b 2b 2b 29 29 29 26 26 26 27 27 27 27 27 27 26 26 26 20 20 20 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 13 13 13 2c 2c 2c 30 30 30 42 42 42 59 59 59 6c 6c 6c 6f 6f 6f 6e 6e 6e 69 69 69 63 63 63 5d 5d 5d 54 54 54 51 51 51 4e 4e 4e 35 35 35 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 25 25 25 34 34 34 34 34 34 31 31 31 33 33 33 2d 2d 2d 27 27 27 25 25 25 22 22 22 19 19 19 0b 0b 0b 18 18 18 18 18 18 14 14 14 0e 0e 0e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 06 06 06 11 11 11 1d 1d 1d 23 23 23 27 27 27 28 28 28 23 23 23 23 23 23 21 21 21 22 22 22 1f 1f 1f 1e 1e 1e 1d 1d 1d 12 12 12 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 1b 1b 1b 27 27 27 20 20 20 17 17 17 12 12 12 09 09 09 0a 0a 0a 07 07 07 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
