((X"#!/", X"bin", X"/ba", X"sh "),
(X"SAV", X"EIF", X"S=$", X"IFS", X" IF", X"S=$", X"(ec", X"ho ", X"-en", X" "\", X"n\b", X"") "),
(X" fo", X"r a", X"rq ", X"in ", X"*.b", X"mp "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"txt", X" ] "),
(X"  t", X"hen", X"   ", X"  e", X"cho", X" "$", X"{ar", X"q::", X"-4}", X""  ", X"   ", X"od ", X"-j ", X"107", X"8 -", X"w29", X"6 -", X"A n", X" -v", X" -t", X" x1", X" $a", X"rq ", X"> "", X"${a", X"rq:", X":-4", X"}".", X"txt", X"   ", X"fi "),
(X"don", X"e "),
(X" fo", X"r a", X"rq ", X"in ", X"*.t", X"xt "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"vhd", X" ] "),
(X"  t", X"hen", X"   ", X"  s", X"aid", X"a="", X"${a", X"rq:", X":-4", X"}".", X"vhd", X"   ", X"  e", X"cho", X" $s", X"aid", X"a  ", X"   ", X"ech", X"o -", X"n "", X"(("", X" >>", X" $s", X"aid", X"a  ", X"   ", X"cat", X" $a", X"rq ", X"| w", X"hil", X"e I", X"FS=", X" re", X"ad ", X"-r ", X"-N ", X"3 i", X"; d", X"o  ", X"   ", X"  i", X"f [", X"[ "", X"$i"", X" ==", X" *$", X"'\n", X"' ]", X"]; ", X"the", X"n  ", X"   ", X"   ", X" ec", X"ho ", X" "X", X"\""", X"$i"", X"\")", X"," ", X">> ", X"$sa", X"ida", X"   ", X"   ", X"   ", X"ech", X"o  ", X"-n ", X""("", X" >>", X" $s", X"aid", X"a  ", X"   ", X"  e", X"lse", X"   ", X"   ", X"   ", X"ech", X"o -", X"n "", X"X\"", X""$i", X""\"", X", "", X" >>", X" $s", X"aid", X"a  ", X"   ", X"  f", X"i  ", X"   ", X"don", X"e  ", X"   ", X"ech", X"o "", X"));", X"" >", X"> $", X"sai", X"da "),
(X"  f", X"i d", X"one", X" "),
(X"# f", X"or ", X"arq", X" in", X" Im", X"g30", X"*.v", X"hd "),
(X"# d", X"o  "),
(X"#  ", X" if", X" [ ", X"$ar", X"q -", X"nt ", X""${", X"arq", X"::-", X"4}"", X".tx", X"t ]", X" # ", X"   ", X" ec", X"ho ", X""${", X"arq", X"::-", X"4}"", X" # ", X"   ", X" # ", X"tou", X"ch ", X""${", X"arq", X"::-", X"4}"", X".tx", X"t #", X"   ", X"  #", X"  #", X"   ", X"  c", X"at ", X"Img", X"301", X"1.v", X"hd ", X"| w", X"hil", X"e r", X"ead", X" -n", X" 3 ", X"i; ", X"do ", X" # ", X"   ", X"   ", X"# i", X"f [", X"$i ", X"== ", X"*$'", X"\n'", X"*] "),
(X"#  ", X"   ", X"   ", X" # ", X"cat", X" "X", X"" $", X"i "", X"),"", X" >>", X" "$", X"{ar", X"q::", X"-4}", X"".t", X"xt;", X"   "),
(X"#  ", X"   ", X"  #", X" el", X"se "),
(X"#  ", X"   ", X"   ", X" # ", X"cat", X" "X", X"\""", X" $i", X" "\", X"","", X" >>", X" "$", X"{ar", X"q::", X"-4}", X"".t", X"xt;", X"  #", X"   ", X"   ", X"   ", X"ech", X"o "", X"leg", X"a" "),
(X"#  ", X"   ", X"  #", X" fi", X" # ", X"   ", X" do", X"ne "),
(X" #", X"   ", X"fi "),
(X"# d", X"one", X" I", X"FS=", X"$SA", X"VEI", X"FS "),
());
((X"#!/", X"bin", X"/ba", X"sh "),
(X"SAV", X"EIF", X"S=$", X"IFS", X" IF", X"S=$", X"(ec", X"ho ", X"-en", X" "\", X"n\b", X"") "),
(X" fo", X"r a", X"rq ", X"in ", X"*.b", X"mp "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"txt", X" ] "),
(X"  t", X"hen", X"   ", X"  e", X"cho", X" "$", X"{ar", X"q::", X"-4}", X""  ", X"   ", X"od ", X"-j ", X"107", X"8 -", X"w29", X"6 -", X"A n", X" -v", X" -t", X" x1", X" $a", X"rq ", X"> "", X"${a", X"rq:", X":-4", X"}".", X"txt", X"   ", X"fi "),
(X"don", X"e "),
(X" fo", X"r a", X"rq ", X"in ", X"*.t", X"xt "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"vhd", X" ] "),
(X"  t", X"hen", X"   ", X"  s", X"aid", X"a="", X"${a", X"rq:", X":-4", X"}".", X"vhd", X"   ", X"  e", X"cho", X" $s", X"aid", X"a  ", X"   ", X"ech", X"o -", X"n "", X"(("", X" >>", X" $s", X"aid", X"a  ", X"   ", X"cat", X" $a", X"rq ", X"| w", X"hil", X"e I", X"FS=", X" re", X"ad ", X"-r ", X"-N ", X"3 i", X"; d", X"o  ", X"   ", X"  i", X"f [", X"[ "", X"$i"", X" ==", X" *$", X"'\n", X"' ]", X"]; ", X"the", X"n  ", X"   ", X"   ", X" ec", X"ho ", X" "X", X"\""", X""${", X"i::", X"2}"", X""\"", X"),"", X"   ", X"   ", X"   ", X"ech", X"o  ", X""X\", X"""$", X"i"\", X""),", X"" >", X"> $", X"sai", X"da "),
(X"   ", X"   ", X"  e", X"cho", X"  -", X"n "", X"(" ", X">> ", X"$sa", X"ida", X"   ", X"   ", X" el", X"se "),
(X"   ", X"   ", X"  e", X"cho", X" -n", X" "X", X"\""", X"$i"", X"\",", X" " ", X">> ", X"$sa", X"ida", X"   ", X"   ", X" fi", X"   ", X"  d", X"one", X"   ", X"  e", X"cho", X" ")", X");"", X" >>", X" $s", X"aid", X"a  ", X" fi", X" do", X"ne "),
(X" #", X" fo", X"r a", X"rq ", X"in ", X"Img", X"30*", X".vh", X"d #", X" do", X"  #", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"txt", X" ] "),
(X"#  ", X"   ", X"ech", X"o "", X"${a", X"rq:", X":-4", X"}" "),
(X"#  ", X"   ", X"# t", X"ouc", X"h "", X"${a", X"rq:", X":-4", X"}".", X"txt", X" # ", X"   ", X" # ", X" # ", X"   ", X" ca", X"t I", X"mg3", X"011", X".vh", X"d |", X" wh", X"ile", X" re", X"ad ", X"-n ", X"3 i", X"; d", X"o  "),
(X"#  ", X"   ", X"  #", X" if", X" [$", X"i =", X"= *", X"$'\", X"n'*", X"] #", X"   ", X"   ", X"   ", X"# c", X"at ", X""X"", X" $i", X" ")", X"," ", X">> ", X""${", X"arq", X"::-", X"4}"", X".tx", X"t; ", X"  #", X"   ", X"   ", X" # ", X"els", X"e #", X"   ", X"   ", X"   ", X"# c", X"at ", X""X\", X""" ", X"$i ", X""\"", X"," ", X">> ", X""${", X"arq", X"::-", X"4}"", X".tx", X"t; ", X" # ", X"   ", X"   ", X"  e", X"cho", X" "l", X"ega", X"" #", X"   ", X"   ", X" # ", X"fi "),
(X"#  ", X"   ", X"don", X"e "),
(X" # ", X"  f", X"i #", X" do", X"ne "),
(X" IF", X"S=$", X"SAV", X"EIF", X"S "),
());
((X"#!/", X"bin", X"/ba", X"sh "),
(X"SAV", X"EIF", X"S=$", X"IFS", X" IF", X"S=$", X"(ec", X"ho ", X"-en", X" "\", X"n\b", X"") "),
(X" fo", X"r a", X"rq ", X"in ", X"*.b", X"mp "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"txt", X" ] "),
(X"  t", X"hen", X"   ", X"  e", X"cho", X" "$", X"{ar", X"q::", X"-4}", X""  ", X"   ", X"od ", X"-j ", X"107", X"8 -", X"w29", X"6 -", X"A n", X" -v", X" -t", X" x1", X" $a", X"rq ", X"> "", X"${a", X"rq:", X":-4", X"}".", X"txt", X"   ", X"fi "),
(X"don", X"e "),
(X" fo", X"r a", X"rq ", X"in ", X"*.t", X"xt "),
(X"do ", X"   ", X"if ", X"[ $", X"arq", X" -n", X"t "", X"${a", X"rq:", X":-4", X"}".", X"vhd", X" ] "),
(X"  t", X"hen", X"   ", X"  s", X"aid", X"a="", X"${a", X"rq:", X":-4", X"}".", X"vhd", X"   ", X"  e", X"cho", X" $s", X"aid", X"a  ", X"   ", X"ech", X"o -", X"n "", X"(("", X" >>", X" $s", X"aid", X"a  ", X"   ", X"cat", X" $a", X"rq ", X"| w", X"hil", X"e I", X"FS=", X" re", X"ad ", X"-r ", X"-N ", X"3 i", X"; d", X"o  ", X"   ", X"  i", X"f [", X"[ "", X"$i"", X" ==", X" *$", X"'\n", X"' ]", X"]; ", X"the", X"n  ", X"   ", X"   ", X" ec", X"ho ", X" "X", X"\"$", X"{i:", X":2}", X"\")", X"," "),
(X"   ", X"   ", X"  e", X"cho", X"  "", X"X\"", X""$i", X""\"", X"),"", X" >>", X" $s", X"aid", X"a  ", X"   ", X"   ", X" ec", X"ho ", X" -n", X" "(", X"" >", X"> $", X"sai", X"da "),
(X"   ", X"   ", X"els", X"e  ", X"   ", X"   ", X" ec", X"ho ", X"-n ", X""X\", X"""$", X"i"\", X"", ", X"" >", X"> $", X"sai", X"da "),
(X"   ", X"   ", X"fi "),
(X"   ", X" do", X"ne "),
(X"   ", X" ec", X"ho ", X""))", X";" ", X">> ", X"$sa", X"ida", X"   ", X"fi "),
(X"don", X"e "),
(X" # ", X"for", X" ar", X"q i", X"n I", X"mg3", X"0*.", X"vhd", X" # ", X"do ", X" # ", X"  i", X"f [", X" $a", X"rq ", X"-nt", X" "$", X"{ar", X"q::", X"-4}", X"".t", X"xt ", X"] #", X"   ", X"  e", X"cho", X" "$", X"{ar", X"q::", X"-4}", X"" #", X"   ", X"  #", X" to", X"uch", X" "$", X"{ar", X"q::", X"-4}", X"".t", X"xt "),
(X"#  ", X"   ", X"#  "),
(X"#  ", X"   ", X"cat", X" Im", X"g30", X"11.", X"vhd", X" | ", X"whi", X"le ", X"rea", X"d -", X"n 3", X" i;", X" do", X"  #", X"   ", X"   ", X" # ", X"if ", X"[$i", X" ==", X" *$", X"'\n", X"'*]", X" # ", X"   ", X"   ", X"  #", X" ca", X"t "", X"X" ", X"$i ", X""),", X"" >", X"> "", X"${a", X"rq:", X":-4", X"}".", X"txt", X";  ", X" # ", X"   ", X"   ", X"# e", X"lse", X" # ", X"   ", X"   ", X"  #", X" ca", X"t "", X"X\"", X"" $", X"i "", X"\",", X"" >", X"> "", X"${a", X"rq:", X":-4", X"}".", X"txt", X";  "),
(X"#  ", X"   ", X"   ", X" ec", X"ho ", X""le", X"ga"", X" # ", X"   ", X"   ", X"# f", X"i #", X"   ", X"  d", X"one", X" "),
(X"#  ", X" fi", X" # ", X"don", X"e "),
(X"IFS", X"=$S", X"AVE", X"IFS", ));
((X"#!", X"bi", X"/b", X"sh"),
(X"SA", X"EI", X"S=", X"IF", X"
I", X"S=", X"(e", X"ho", X"-e", X" "", X"n\", X"")"),
(X"
f", X"r ", X"rq", X"in", X"*.", X"mp"),
(X"do", X"
 ", X"if", X"[ ", X"ar", X" -", X"t ", X"${", X"rq", X":-", X"}"", X"tx", X" ]"),
(X"  ", X"he", X"
 ", X"  ", X"ch", X" "", X"{a", X"q:", X"-4", X""
", X"  ", X"od", X"-j", X"10", X"8 ", X"w2", X"6 ", X"A ", X" -", X" -", X" x", X" $", X"rq", X"> ", X"${", X"rq", X":-", X"}"", X"tx", X"
 ", X"fi"),
(X"do", X"e
"),
(X"
f", X"r ", X"rq", X"in", X"*.", X"xt"),
(X"do", X"
 ", X"if", X"[ ", X"ar", X" -", X"t ", X"${", X"rq", X":-", X"}"", X"vh", X" ]"),
(X"  ", X"he", X"
 ", X"  ", X"ai", X"a=", X"${", X"rq", X":-", X"}"", X"vh", X"
 ", X"  ", X"ch", X" $", X"ai", X"a
", X"  ", X"ec", X"o ", X"n ", X"((", X" >", X" $", X"ai", X"a
", X"  ", X"ca", X" $", X"rq", X"| ", X"hi", X"e ", X"FS", X" r", X"ad", X"-r", X"-N", X"3 ", X"; ", X"o
", X"  ", X"  ", X"f ", X"[ ", X"$i", X" =", X" *", X"'\", X"' ", X"];", X"th", X"n
", X"  ", X"  ", X" e", X"ho", X" "", X"\"", X"{i", X":2", X"\"", X","", X">>", X"$s", X"id", X"
 ", X"  ", X"  ", X"ec", X"o ", X"-n", X""(", X" >", X" $", X"ai", X"a
", X"  ", X"  ", X"ls", X"
 ", X"  ", X"  ", X"ec", X"o ", X"n ", X"X\", X"${", X"::", X"}\", X", ", X" >", X" $", X"ai", X"a
", X"  ", X"  ", X"i
", X"  ", X"do", X"e
", X"  ", X"ec", X"o ", X"))", X"" ", X"> ", X"sa", X"da"),
(X"  ", X"i
", X"on", X"

"),
(X"# ", X"or", X"ar", X" i", X" I", X"g3", X"*.", X"hd"),
(X"# ", X"o "),
(X"# ", X" i", X" [", X"$a", X"q ", X"nt", X""$", X"ar", X"::", X"4}", X".t", X"t ", X"
#", X"  ", X" e", X"ho", X""$", X"ar", X"::", X"4}", X"
#", X"  ", X" #", X"to", X"ch", X""$", X"ar", X"::", X"4}", X".t", X"t
", X"  ", X"  ", X" 
", X"  ", X"  ", X"at", X"Im", X"30", X"1.", X"hd", X"| ", X"hi", X"e ", X"ea", X" -", X" 3", X"i;", X"do", X"
#", X"  ", X"  ", X"# ", X"f ", X"$i", X"==", X"*$", X"\n", X"*]"),
(X"# ", X"  ", X"  ", X" #", X"ca", X" "", X"" ", X"i ", X"),", X" >", X" "", X"{a", X"q:", X"-4", X"".", X"xt", X"  "),
(X"# ", X"  ", X"  ", X" e", X"se"),
(X"# ", X"  ", X"  ", X" #", X"ca", X" "", X"\"", X" $", X" "", X"",", X" >", X" "", X"{a", X"q:", X"-4", X"".", X"xt", X" 
", X"  ", X"  ", X"  ", X"ec", X"o ", X"le", X"a""),
(X"# ", X"  ", X"  ", X" f", X"
#", X"  ", X" d", X"ne"),
(X"

", X"  ", X"fi"),
(X"# ", X"on", X"

", X"FS", X"$S", X"VE", X"FS"),
());
((X"#!",X"bi",X"/b",X"sh"),
(X"SA",X"EI",X"S=",X"IF",X"
I",X"S=",X"(e",X"ho",X"-e",X" "",X"n\",X"")"),
(X"
f",X"r ",X"rq",X"in",X"*.",X"mp"),
(X"do",X"
 ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]"),
(X"  ",X"he",X"
 ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
",X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx",X"
 ",X"fi"),
(X"do",X"e
"),
(X"
f",X"r ",X"rq",X"in",X"*.",X"xt"),
(X"do",X"
 ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"vh",X" ]"),
(X"  ",X"he",X"
 ",X"  ",X"ai",X"a=",X"${",X"rq",X":-",X"}"",X"vh",X"
 ",X"  ",X"ch",X" $",X"ai",X"a
",X"  ",X"ec",X"o ",X"n ",X"((",X" >",X" $",X"ai",X"a
",X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X" r",X"ad",X"-r",X"-N",X"3 ",X"; ",X"o
",X"  ",X"  ",X"f ",X"[ ",X"$i",X" =",X" *",X"'\",X"' ",X"];",X"th",X"n
",X"  ",X"  ",X" e",X"ho",X" "",X"\"",X"{i",X":2",X"\"",X","",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"ec",X"o ",X"-n",X""(",X" >",X" $",X"ai",X"a
",X"  ",X"  ",X"ls",X"
 ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X"::",X"}\",X","",X">>",X"$s",X"id",X"
 ",X"  ",X" f",X"
 ",X"  ",X"on",X"
 ",X"  ",X"ch",X" "",X");",X" >",X" $",X"ai",X"a
",X" f",X"
d",X"ne"),
(X"

",X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
",X" d",X" 
",X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]"),
(X"# ",X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}""),
(X"# ",X"  ",X"# ",X"ou",X"h ",X"${",X"rq",X":-",X"}"",X"tx",X"
#",X"  ",X" #",X"
#",X"  ",X" c",X"t ",X"mg",X"01",X".v",X"d ",X" w",X"il",X" r",X"ad",X"-n",X"3 ",X"; ",X"o "),
(X"# ",X"  ",X"  ",X" i",X" [",X"i ",X"= ",X"$'",X"n'",X"]
",X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
",X"  ",X"  ",X" #",X"el",X"e
",X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X"
#",X"  ",X"  ",X"  ",X"ch",X" "",X"eg",X""
",X"  ",X"  ",X" #",X"fi"),
(X"# ",X"  ",X"do",X"e
"),
(X"
#",X"  ",X"i
",X" d",X"ne"),
(X"
I",X"S=",X"SA",X"EI",X"S
"),
());
((X"#!/",X"bin",X"/ba",X"sh
"),
(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"",X"-en",X""\",X"n\b",X"")
"),
(X"
fo",X"a",X"",X"",X"*.b",X"mp
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"]
"),
(X"t",X"hen",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X"",X"",X"",X"",X"107",X"-",X"w29",X"-",X"n",X"-v",X"-t",X"x1",X"$a",X"",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"fi
"),
(X"don",X"e

"),
(X"
fo",X"a",X"",X"",X"*.t",X"xt
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"]
"),
(X"t",X"hen",X"",X"s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"",X"e",X"cho",X"$s",X"aid",X"",X"",X"ech",X"-",X""",X"(("",X">>",X"$s",X"aid",X"",X"",X"cat",X"$a",X"",X"w",X"hil",X"I",X"FS=",X"re",X"",X"",X"",X"i",X"d",X"",X"",X"i",X"[",X""",X"$i"",X"==",X"*$",X"'\n",X"]",X"",X"the",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"}\"",X"),"",X">>",X"$s",X"aid",X"",X"",X"",X"ec",X"",X"-n",X""(",X">",X"$",X"sai",X"da
"),
(X"",X"",X"els",X"",X"",X"",X"ec",X"",X"",X""X\",X""${",X"i##",X"}",X"\",",X">",X"$",X"sai",X"da
"),
(X"",X"",X"fi
"),
(X"",X"do",X"ne
"),
(X"",X"ec",X"",X""))",X"",X"",X"$sa",X"ida",X"",X"fi
"),
(X"don",X"e

"),
(X"",X"for",X"ar",X"i",X"I",X"mg3",X"0*.",X"vhd",X"",X"",X"",X"i",X"[",X"$a",X"",X"-nt",X""$",X"{ar",X"q::",X"-4}",X"".t",X"",X"]
#",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X""
#",X"",X"#",X"to",X"uch",X""$",X"{ar",X"q::",X"-4}",X"".t",X"xt
"),
(X"",X"",X"
"),
(X"",X"",X"cat",X"Im",X"g30",X"11.",X"vhd",X"",X"whi",X"",X"rea",X"-",X"3",X"i;",X"do",X"
#",X"",X"",X"",X"",X"[$i",X"==",X"*$",X"'\n",X"'*]",X"",X"",X"",X"#",X"ca",X""",X"",X"",X""),",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"",X"",X"",X"e",X"lse",X"",X"",X"",X"#",X"ca",X""",X"X\"",X"$",X""",X"\",",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"
"),
(X"",X"",X"",X"ec",X"",X""le",X"ga"",X"",X"",X"",X"f",X"i
#",X"",X"d",X"one",X"


"),
(X"",X"fi",X"",X"don",X"e

"),
(X"IFS",X"=$S",X"AVE",X"IFS",));
((X"#!/",X"bin",X"/ba",X"sh
"),(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"",X"-en",X""\",X"n\b",X"")
"),(X"
fo",X"a",X"",X"",X"*.b",X"mp
"),(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"]
"),(X"t",X"hen",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X"",X"",X"",X"",X"107",X"-",X"w29",X"-",X"n",X"-v",X"-t",X"x1",X"$a",X"",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"fi
"),(X"don",X"e

"),(X"
fo",X"a",X"",X"",X"*.t",X"xt
"),(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"]
"),(X"t",X"hen",X"",X"s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"",X"e",X"cho",X"$s",X"aid",X"",X"",X"ech",X"-",X""",X"(("",X">>",X"$s",X"aid",X"",X"",X"cat",X"$a",X"",X"w",X"hil",X"I",X"FS=",X"re",X"",X"",X"",X"i",X"d",X"",X"",X"i",X"[",X""",X"$i"",X"==",X"*$",X"'\n",X"]",X"",X"the",X"",X"",X"",X"ec",X"",X"-n",X""X",X"\"$",X"{i#",X"",X"}\"",X"),"",X">>",X"$s",X"aid",X"",X"",X"",X"ec",X"",X"-n",X""(",X">",X"$",X"sai",X"da
"),(X"",X"",X"els",X"",X"",X"",X"ec",X"",X"",X""X\",X""${",X"i##",X"}",X"\",",X">",X"$",X"sai",X"da
"),(X"",X"",X"fi
"),(X"",X"do",X"ne
"),(X"",X"ec",X"",X""))",X"",X"",X"$sa",X"ida",X"",X"fi
"),(X"don",X"e

"),(X"",X"for",X"ar",X"i",X"I",X"mg3",X"0*.",X"vhd",X"",X"",X"",X"i",X"[",X"$a",X"",X"-nt",X""$",X"{ar",X"q::",X"-4}",X"".t",X"",X"]
#",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X""
#",X"",X"#",X"to",X"uch",X""$",X"{ar",X"q::",X"-4}",X"".t",X"xt
"),(X"",X"",X"
"),(X"",X"",X"cat",X"Im",X"g30",X"11.",X"vhd",X"",X"whi",X"",X"rea",X"-",X"3",X"i;",X"do",X"
#",X"",X"",X"",X"",X"[$i",X"==",X"*$",X"'\n",X"'*]",X"",X"",X"",X"#",X"ca",X""",X"",X"",X""),",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"",X"",X"",X"e",X"lse",X"",X"",X"",X"#",X"ca",X""",X"X\"",X"$",X""",X"\",",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"
"),(X"",X"",X"",X"ec",X"",X""le",X"ga"",X"",X"",X"",X"f",X"i
#",X"",X"d",X"one",X"


"),(X"",X"fi",X"",X"don",X"e

"),(X"IFS",X"=$S",X"AVE",X"IFS",));
((X"#!/",X"bin",X"/ba",X"sh
"),
(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"",X"-en",X""\",X"n\b",X"")
"),
(X"
fo",X"a",X"",X"",X"*.b",X"mp
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"]
"),
(X"t",X"hen",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X"",X"",X"",X"",X"107",X"-",X"w29",X"-",X"n",X"-v",X"-t",X"x1",X"$a",X"",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"fi
"),
(X"don",X"e

"),
(X"
fo",X"a",X"",X"",X"*.t",X"xt
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"]
"),
(X"t",X"hen",X"",X"s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"",X"e",X"cho",X"$s",X"aid",X"",X"",X"ech",X"-",X""",X"(("",X">>",X"$s",X"aid",X"",X"",X"cat",X"$a",X"",X"w",X"hil",X"I",X"FS=",X"re",X"",X"",X"",X"i",X"d",X"",X"",X"i",X"[",X""",X"$i"",X"==",X"*$",X"'\n",X"]",X"",X"the",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"}\"",X"),"",X"",X"",X"",X"ech",X"",X""X\",X""${",X"i##",X"}",X"\")",X"",X"",X"$sa",X"ida",X"",X"",X"",X"ech",X"",X"",X""("",X">>",X"$s",X"aid",X"",X"",X"e",X"lse",X"",X"",X"",X"ech",X"-",X""",X"X\"",X"${i",X"##*",X"}\",X"","",X">>",X"$s",X"aid",X"",X"",X"f",X"",X"",X"don",X"",X"",X"ech",X""",X"));",X">",X"$",X"sai",X"da
"),
(X"f",X"i
d",X"one",X"


"),
(X"f",X"",X"arq",X"in",X"Im",X"g30",X"*.v",X"hd
"),
(X"d",X"
"),
(X"",X"if",X"",X"$ar",X"-",X"",X""${",X"arq",X"::-",X"4}"",X".tx",X"]",X"",X"",X"ec",X"",X""${",X"arq",X"::-",X"4}"",X"",X"",X"",X"tou",X"",X""${",X"arq",X"::-",X"4}"",X".tx",X"t
#",X"",X"#",X"
#",X"",X"c",X"",X"Img",X"301",X"1.v",X"",X"w",X"hil",X"r",X"ead",X"-n",X"",X"",X"",X"",X"",X"",X"i",X"[",X"",X"",X"*$'",X"\n'",X"*]
"),
(X"",X"",X"",X"",X"cat",X""X",X"$",X""",X"),"",X">>",X""$",X"{ar",X"q::",X"-4}",X"".t",X"xt;",X"
"),
(X"",X"",X"#",X"el",X"se
"),
(X"",X"",X"",X"",X"cat",X""X",X"\""",X"$i",X""\",X"","",X">>",X""$",X"{ar",X"q::",X"-4}",X"".t",X"xt;",X"
#",X"",X"",X"",X"ech",X""",X"leg",X"a"
"),
(X"",X"",X"#",X"fi",X"",X"",X"do",X"ne
"),
(X"

#",X"",X"fi
"),
(X"d",X"one",X"

I",X"FS=",X"$SA",X"VEI",X"FS
"),
());
((X"#!/",X"bin",X"/ba",X"sh
"),
(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"",X"-en",X""\",X"n\b",X"")
"),
(X"
fo",X"a",X"",X"",X"*.b",X"mp
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"]
"),
(X"t",X"hen",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X"",X"",X"",X"",X"107",X"-",X"w29",X"-",X"n",X"-v",X"-t",X"x1",X"$a",X"",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"fi
"),
(X"don",X"e

"),
(X"
fo",X"a",X"",X"",X"*.t",X"xt
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"]
"),
(X"t",X"hen",X"",X"s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"",X"e",X"cho",X"$s",X"aid",X"",X"",X"ech",X"-",X""",X"(("",X">>",X"$s",X"aid",X"",X"",X"cat",X"$a",X"",X"w",X"hil",X"I",X"FS=",X"re",X"",X"",X"",X"i",X"d",X"",X"",X"i",X"[",X""",X"$i"",X"==",X"*$",X"'\n",X"]",X"",X"the",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"::-",X"1}\",X""),",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"}\"",X"),"",X">>",X"$s",X"aid",X"",X"",X"",X"ec",X"",X"-n",X""(",X">",X"$",X"sai",X"da
"),
(X"",X"",X"els",X"",X"",X"",X"ec",X"",X"",X""X\",X""${",X"i##",X"}",X"\",",X">",X"$",X"sai",X"da
"),
(X"",X"",X"fi
"),
(X"",X"do",X"ne
"),
(X"",X"ec",X"",X""))",X"",X"",X"$sa",X"ida",X"",X"fi
"),
(X"don",X"e

"),
(X"",X"for",X"ar",X"i",X"I",X"mg3",X"0*.",X"vhd",X"",X"",X"",X"i",X"[",X"$a",X"",X"-nt",X""$",X"{ar",X"q::",X"-4}",X"".t",X"",X"]
#",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X""
#",X"",X"#",X"to",X"uch",X""$",X"{ar",X"q::",X"-4}",X"".t",X"xt
"),
(X"",X"",X"
"),
(X"",X"",X"cat",X"Im",X"g30",X"11.",X"vhd",X"",X"whi",X"",X"rea",X"-",X"3",X"i;",X"do",X"
#",X"",X"",X"",X"",X"[$i",X"==",X"*$",X"'\n",X"'*]",X"",X"",X"",X"#",X"ca",X""",X"",X"",X""),",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"",X"",X"",X"e",X"lse",X"",X"",X"",X"#",X"ca",X""",X"X\"",X"$",X""",X"\",",X">",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"
"),
(X"",X"",X"",X"ec",X"",X""le",X"ga"",X"",X"",X"",X"f",X"i
#",X"",X"d",X"one",X"


"),
(X"",X"fi",X"",X"don",X"e

"),
(X"IFS",X"=$S",X"AVE",X"IFS",));
((X"#!/",X"bin",X"/ba",X"sh
"),
(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"",X"-en",X""\",X"n\b",X"")
"),
(X"
fo",X"a",X"",X"",X"*.b",X"mp
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X" ]
"),
(X"t",X"hen",X"",X"e",X"cho",X""$",X"{ar",X"q::",X"-4}",X"",X"",X"",X"",X"107",X"-",X"w29",X"-",X"n",X"-v",X"-t",X"x1",X"$a",X"",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"fi
"),
(X"don",X"e

"),
(X"
fo",X"a",X"",X"",X"*.t",X"xt
"),
(X"",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"vhd",X" ]
"),
(X"t",X"hen",X"",X"s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"",X"e",X"cho",X"$s",X"aid",X"",X"",X"ech",X"-",X""",X"(("",X">>",X"$s",X"aid",X"",X"",X"cat",X"$a",X"",X"w",X"hil",X"I",X"FS=",X"re",X"",X"",X"",X"i",X"d",X"",X"",X"i",X"[",X""",X"$i"",X"==",X"*$",X"'\n",X"]",X"",X"the",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"::-",X"1}\",X""),",X"",X"",X"",X"ec",X"",X""X",X"\"$",X"{i#",X"",X"::-",X"1}\",X""),",X">",X"$",X"sai",X"da
"),
(X"",X"",X"e",X"cho",X"-",X""",X"",X"",X"$sa",X"ida",X"",X"",X"el",X"se
"),
(X"",X"",X"e",X"cho",X"-n",X""X",X"\"$",X"{i#",X"",X"}\"",X"",X"",X"$sa",X"ida",X"",X"",X"fi",X"",X"d",X"one",X"",X"e",X"cho",X"")",X");"",X">>",X"$s",X"aid",X"",X"fi",X"
do",X"ne
"),
(X"

#",X"fo",X"a",X"",X"",X"Img",X"30*",X".vh",X"d
#",X"do",X"
#",X"",X"",X"$",X"arq",X"-n",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X" ]
"),
(X"",X"",X"ech",X""",X"${a",X"rq:",X":-4",X"}"
"),
(X"",X"",X"t",X"ouc",X""",X"${a",X"rq:",X":-4",X"}".",X"txt",X"",X"",X"",X"",X"",X"ca",X"I",X"mg3",X"011",X".vh",X"|",X"wh",X"ile",X"re",X"",X"",X"i",X"d",X"o 
"),
(X"",X"",X"#",X"if",X"[$",X"=",X"*",X"$'\",X"n'*",X"]
#",X"",X"",X"",X"c",X"",X""X"",X"$i",X"")",X"",X"",X""${",X"arq",X"::-",X"4}"",X".tx",X"",X"
#",X"",X"",X"",X"els",X"e
#",X"",X"",X"",X"c",X"",X""X\",X"",X"",X""\"",X"",X"",X""${",X"arq",X"::-",X"4}"",X".tx",X"",X"",X"",X"",X"e",X"cho",X""l",X"ega",X""
#",X"",X"",X"",X"fi
"),
(X"",X"",X"don",X"e

"),
(X"",X"f",X"i
#",X"do",X"ne
"),
(X"
IF",X"S=$",X"SAV",X"EIF",X"S

"),
());
((X"#!/",X"bin",X"/ba",X"sh
"),
(X"SAV",X"EIF",X"S=$",X"IFS",X"
IF",X"S=$",X"(ec",X"ho ",X"-en",X" "\",X"n\b",X"")
"),
(X"
fo",X"r a",X"rq ",X"in ",X"*.b",X"mp
"),
(X"do ",X"
  ",X"if ",X"[ $",X"arq",X" -n",X"t "",X"${a",X"rq:",X":-4",X"}".",X"txt",X" ]
"),
(X"  t",X"hen",X"
  ",X"  e",X"cho",X" "$",X"{ar",X"q::",X"-4}",X""
 ",X"   ",X"od ",X"-j ",X"107",X"8 -",X"w29",X"6 -",X"A n",X" -v",X" -t",X" x1",X" $a",X"rq ",X"> "",X"${a",X"rq:",X":-4",X"}".",X"txt",X"
  ",X"fi
"),
(X"don",X"e

"),
(X"
fo",X"r a",X"rq ",X"in ",X"*.t",X"xt
"),
(X"do ",X"
  ",X"if ",X"[ $",X"arq",X" -n",X"t "",X"${a",X"rq:",X":-4",X"}".",X"vhd",X" ]
"),
(X"  t",X"hen",X"
  ",X"  s",X"aid",X"a="",X"${a",X"rq:",X":-4",X"}".",X"vhd",X"
  ",X"  e",X"cho",X" $s",X"aid",X"a
 ",X"   ",X"ech",X"o -",X"n "",X"(("",X" >>",X" $s",X"aid",X"a
 ",X"   ",X"cat",X" $a",X"rq ",X"| w",X"hil",X"e I",X"FS=",X" re",X"ad ",X"-r ",X"-N ",X"3 i",X"; d",X"o
 ",X"   ",X"  i",X"f [",X"[ "",X"$i"",X" ==",X" *$",X"'\n",X"' ]",X"]; ",X"the",X"n
 ",X"   ",X"   ",X" ec",X"ho ",X" "X",X"\"$",X"{i:",X"-2}",X"\")",X","
"),
(X"   ",X"   ",X"  e",X"cho",X"  "",X"X\"",X"${i",X":-2",X"}\"",X"),"",X" >>",X" $s",X"aid",X"a
 ",X"   ",X"   ",X" ec",X"ho ",X" -n",X" "(",X"" >",X"> $",X"sai",X"da
"),
(X"   ",X"   ",X"els",X"e
 ",X"   ",X"   ",X" ec",X"ho ",X"-n ",X""X\",X""${",X"i:-",X"2}\",X"","",X" >>",X" $s",X"aid",X"a
 ",X"   ",X"  f",X"i
 ",X"   ",X"don",X"e
 ",X"   ",X"ech",X"o "",X"));",X"" >",X"> $",X"sai",X"da
"),
(X"  f",X"i
d",X"one",X"


"),
(X"# f",X"or ",X"arq",X" in",X" Im",X"g30",X"*.v",X"hd
"),
(X"# d",X"o 
"),
(X"#  ",X" if",X" [ ",X"$ar",X"q -",X"nt ",X""${",X"arq",X"::-",X"4}"",X".tx",X"t ]",X"
# ",X"   ",X" ec",X"ho ",X""${",X"arq",X"::-",X"4}"",X"
# ",X"   ",X" # ",X"tou",X"ch ",X""${",X"arq",X"::-",X"4}"",X".tx",X"t
#",X"   ",X"  #",X" 
#",X"   ",X"  c",X"at ",X"Img",X"301",X"1.v",X"hd ",X"| w",X"hil",X"e r",X"ead",X" -n",X" 3 ",X"i; ",X"do ",X"
# ",X"   ",X"   ",X"# i",X"f [",X"$i ",X"== ",X"*$'",X"\n'",X"*]
"),
(X"#  ",X"   ",X"   ",X" # ",X"cat",X" "X",X"" $",X"i "",X"),"",X" >>",X" "$",X"{ar",X"q::",X"-4}",X"".t",X"xt;",X"  
"),
(X"#  ",X"   ",X"  #",X" el",X"se
"),
(X"#  ",X"   ",X"   ",X" # ",X"cat",X" "X",X"\""",X" $i",X" "\",X"","",X" >>",X" "$",X"{ar",X"q::",X"-4}",X"".t",X"xt;",X" 
#",X"   ",X"   ",X"   ",X"ech",X"o "",X"leg",X"a"
"),
(X"#  ",X"   ",X"  #",X" fi",X"
# ",X"   ",X" do",X"ne
"),
(X"

#",X"   ",X"fi
"),
(X"# d",X"one",X"

I",X"FS=",X"$SA",X"VEI",X"FS
"),
());
((X"!/",X"in",X"ba",X"h
"),
(X"AV",X"IF",X"=$",X"FS",X"IF",X"=$",X"ec",X"o ",X"en",X""\",X"\b",X")
"),
(X"fo",X" a",X"q ",X"n ",X".b",X"p
"),
(X"o ",X"  ",X"f ",X" $",X"rq",X"-n",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"]
"),
(X" t",X"en",X"  ",X" e",X"ho",X""$",X"ar",X"::",X"4}",X"
 ",X"  ",X"d ",X"j ",X"07",X" -",X"29",X" -",X" n",X"-v",X"-t",X"x1",X"$a",X"q ",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"  ",X"i
"),
(X"on",X"

"),
(X"fo",X" a",X"q ",X"n ",X".t",X"t
"),
(X"o ",X"  ",X"f ",X" $",X"rq",X"-n",X" "",X"{a",X"q:",X"-4",X"".",X"hd",X"]
"),
(X" t",X"en",X"  ",X" s",X"id",X"="",X"{a",X"q:",X"-4",X"".",X"hd",X"  ",X" e",X"ho",X"$s",X"id",X"
 ",X"  ",X"ch",X" -",X" "",X"("",X">>",X"$s",X"id",X"
 ",X"  ",X"at",X"$a",X"q ",X" w",X"il",X" I",X"S=",X"re",X"d ",X"r ",X"N ",X" i",X" d",X"
 ",X"  ",X" i",X" [",X" "",X"i"",X"==",X"*$",X"\n",X" ]",X"; ",X"he",X"
 ",X"  ",X"  ",X"ec",X"o ",X""X",X""$",X"i:",X"-2",X"\"",X","",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"ec",X"o ",X"-n",X""(",X" >",X" $",X"ai",X"a
"),
(X"  ",X"  ",X"ls",X"
 ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
"),
(X"  ",X"  ",X"i
"),
(X"  ",X"do",X"e
"),
(X"  ",X"ec",X"o ",X"))",X"" ",X"> ",X"sa",X"da",X"  ",X"i
"),
(X"on",X"

"),
(X"# ",X"or",X"ar",X" i",X" I",X"g3",X"*.",X"hd",X"# ",X"o ",X"# ",X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",X"
#",X"  ",X" e",X"ho",X""$",X"ar",X"::",X"4}",X"
#",X"  ",X" #",X"to",X"ch",X""$",X"ar",X"::",X"4}",X".t",X"t
"),
(X"  ",X"  ",X" 
"),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do",X"
#",X"  ",X"  ",X"# ",X"f ",X"$i",X"==",X"*$",X"\n",X"*]",X"# ",X"  ",X"  ",X" #",X"ca",X" "",X"" ",X"i ",X"),",X" >",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"  ",X"# ",X"  ",X"  ",X" e",X"se",X"# ",X"  ",X"  ",X" #",X"ca",X" "",X"\"",X" $",X" "",X"",",X" >",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X" 
"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a"",X"# ",X"  ",X"  ",X" f",X"
#",X"  ",X" d",X"ne",X"

"),
(X"  ",X"fi",X"# ",X"on",X"

"),
(X"FS",X"$S",X"VE",X"FS",));
((X"!/",X"in",X"ba",X"sh
"),
(X"AV",X"IF",X"=$",X"FS",X"IF",X"=$",X"ec",X"o ",X"en",X""\",X"\b",X"")
"),
(X"fo",X" a",X"q ",X"n ",X".b",X"mp
"),
(X"o ",X"  ",X"f ",X" $",X"rq",X"-n",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X" ]
"),
(X" t",X"en",X"  ",X" e",X"ho",X""$",X"ar",X"::",X"4}",X"
 ",X"  ",X"d ",X"j ",X"07",X" -",X"29",X" -",X" n",X"-v",X"-t",X"x1",X"$a",X"q ",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"  ",X"fi
"),
(X"on",X"e

"),
(X"fo",X" a",X"q ",X"n ",X".t",X"xt
"),
(X"o ",X"  ",X"f ",X" $",X"rq",X"-n",X" "",X"{a",X"q:",X"-4",X"".",X"hd",X" ]
"),
(X" t",X"en",X"  ",X" s",X"id",X"="",X"{a",X"q:",X"-4",X"".",X"hd",X"  ",X" e",X"ho",X"$s",X"id",X"
 ",X"  ",X"ch",X" -",X" "",X"("",X">>",X"$s",X"id",X"
 ",X"  ",X"at",X"$a",X"q ",X" w",X"il",X" I",X"S=",X"re",X"d ",X"r ",X"N ",X" i",X" d",X"
 ",X"  ",X" i",X" [",X" "",X"i"",X"==",X"*$",X"\n",X" ]",X"; ",X"he",X"
 ",X"  ",X"  ",X"ec",X"o ",X""X",X""$",X"\"",X","",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"ec",X"o ",X"-n",X""(",X" >",X" $",X"ai",X"da
"),
(X"  ",X"  ",X"ls",X"
 ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"da
"),
(X"  ",X"  ",X"fi
"),
(X"  ",X"do",X"ne
"),
(X"  ",X"ec",X"o ",X"))",X"" ",X"> ",X"sa",X"da",X"  ",X"fi
"),
(X"on",X"e

"),
(X"# ",X"or",X"ar",X" i",X" I",X"g3",X"*.",X"hd",X"# ",X"o ",X"# ",X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",X"
#",X"  ",X" e",X"ho",X""$",X"ar",X"::",X"4}",X"
#",X"  ",X" #",X"to",X"ch",X""$",X"ar",X"::",X"4}",X".t",X"xt
"),
(X"  ",X"  ",X"# 
"),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do",X"
#",X"  ",X"  ",X"# ",X"f ",X"$i",X"==",X"*$",X"\n",X"*]",X"# ",X"  ",X"  ",X" #",X"ca",X" "",X"" ",X"i ",X"),",X" >",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"  ",X"# ",X"  ",X"  ",X" e",X"se",X"# ",X"  ",X"  ",X" #",X"ca",X" "",X"\"",X" $",X" "",X"",",X" >",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"; 
"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a"",X"# ",X"  ",X"  ",X" f",X"
#",X"  ",X" d",X"ne",X"


"),
(X"  ",X"fi",X"# ",X"on",X"e

"),
(X"FS",X"$S",X"VE",X"FS",));
((X"!/",X"in",X"ba",(
));
((X"!/",X"in",X"ba",(
X""),X"VE",X"FS",X"$I",(
X""),X"S=",X"(e",X"ho",X"-e",X" "",X"n\",X"")",X"
f",X"r ",X"rq",X"in",X"*.",X"mp",X"do",X"
 ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]",X"  ",X"he",X"
 ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",(
X""),X"  ",X"d ",X"j ",X"07",X" -",X"29",X" -",X" n",X"-v",X"-t",X"x1",X"$a",X"q ",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"  ",(
X""),X"ne",(
X""),X"r ",X"rq",X"in",X"*.",X"xt",X"do",X"
 ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"vh",X" ]",X"  ",X"he",X"
 ",X"  ",X"ai",X"a=",X"${",X"rq",X":-",X"}"",X"vh",X"
 ",X"  ",X"ch",X" $",X"ai",(
X""),X"  ",X"ch",X" -",X" "",X"("",X">>",X"$s",X"id",X"
 ",X"  ",X"at",X"$a",X"q ",X" w",X"il",X" I",X"S=",X"re",X"d ",X"r ",X"N ",X" i",X" d",X"
 ",X"  ",X" i",X" [",X" "",X"i"",X"==",X"*$",X"\n",X" ]",X"; ",X"he",X"
 ",X"  ",X"  ",X"re",X"d ",X"r ",X"N ",X" i",X"  ",X"  ",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"ec",X"o ",X"-n",X""X",X""$",X"i:",X"-2",X"\"",X","",X">>",X"$s",X"id",X"
 ",X"  ",X" e",X"se",X"  ",X"  ",X"  ",X"ch",X" -",X" "",X"\"",X"{i",X" -",X"}\",X","",X">>",X"$s",X"id",X"
 ",X"  ",X" f",X"
 ",X"  ",X"on",X"
 ",X"  ",X"ch",X" "",X");",X" >",X" $",X"ai",(
X""),X"fi",X"do",(
X""),X"# ",X"or",X"ar",X" i",X" I",X"g3",X"*.",X"hd",X"# ",X"o ",X"# ",X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",X"
#",X"  ",X" e",X"ho",X""$",X"ar",X"::",X"4}",X"
#",X"  ",X" #",X"to",X"ch",X""$",X"ar",X"::",X"4}",X".t",(
X""),X"  ",X" #",X"
#",X"  ",X" c",X"t ",X"mg",X"01",X".v",X"d ",X" w",X"il",X" r",X"ad",X"-n",X"3 ",X"; ",X"o ",X"# ",X"  ",X"  ",X" i",X" [",X"i ",X"= ",X"$'",X"n'",(
X""),X"  ",X"  ",X"  ",X" c",X"t ",X"X"",X"$i",X"")",X"" ",X"> ",X"${",X"rq",X":-",X"}"",X"tx",X"; ",X"
#",X"  ",X"  ",X"# ",X"ls",X"
#",X"  ",X"  ",X"  ",X" c",X"t ",X"X\",X"" ",X"i ",X"\"",X"" ",X"> ",X"${",X"rq",X":-",X"}"",X"tx",X"; ",X"# ",X"  ",X"  ",X" e",X"ho",X""l",X"ga",X"
#",X"  ",X"  ",X"# ",(
X""),X"  ",X" d",X"ne",(
X""),X"  ",(
X""),X"do",(
X""),X"FS",X"$S",X"VE",X"FS",));
(((
),
(
),
(
),
(
X"or",X"ar",X" i",X" *",X"bm",X"
d",X" 
",X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",X"
 ",X"th",X"n
",X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}"",X"  ",X" o",X" -",X" 1",X"78",X"-w",X"96",X"-A",X"n ",X"v ",X"t ",X"1 ",X"ar",X" >",X""$",X"ar",X"::",X"4}",X".t",X"t
",X" f",X"
d",X"ne",X"

",X"or",X"ar",X" i",X" *",X"tx",X"
d",X" 
",X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d ",X"
 ",X"th",X"n
",X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
",X"  ",X"ec",X"o ",X"sa",X"da",X"  ",X" e",X"ho",X"-n",X""(",X"" ",X"> ",X"sa",X"da",X"  ",X" c",X"t ",X"ar",X" |",X"wh",X"le",X"IF",X"='",X" r",X"ad",X"-r",X"li",X"e ",X"| ",X"[ ",X"n ",X"$l",X"ne",X" ]",X"; ",X"o
",X"  ",X"  ",X"ch",X" "",X"" ",X"> ",X"sa",X"da",X"  ",X"  ",X"ca",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do",X"  ",X"  ",X"  ",X" i",X" [",X" "",X"i"",X"==",X"*$",X"\n",X" ]",X"; ",X"he",X"
 ",X"  ",X"  ",X"# ",X" e",X"ho",X" "",X"" ",X"> ",X"sa",X"da",X"  ",X"  ",X"  ",X"  ",X"ec",X"o ",X"-n",X""X",X""$",X"i:",X"-2",X"\"",X","",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"# ",X"ls",X"
 ",X"  ",X"  ",X"  ",X"ch",X" -",X" "",X"\"",X"{i",X" -",X"}\",X","",X">>",X"$s",X"id",X"
 ",X"  ",X"  ",X"# ",X"i
",X"  ",X"  ",X"on",X"
 ",X"  ",X" e",X"ho",X"")",X"" ",X"> ",X"sa",X"da",X"  ",X" d",X"ne",X"  ",X" e",X"ho",X"")",X";"",X">>",X"$s",X"id",X"
 ",X"fi",X"do",X"e
",X"
#",X"fo",X" a",X"q ",X"n ",X"mg",X"0*",X"vh",X"
#",X"do",X"
#",X"  ",X"f ",X" $",X"rq",X"-n",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"]
",X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
",X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt",X"# ",X"  ",X"# ",X"# ",X"  ",X"ca",X" I",X"g3",X"11",X"vh",X" |",X"wh",X"le",X"re",X"d ",X"n ",X" i",X" d",X" 
",X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*",X"
#",X"  ",X"  ",X"  ",X" c",X"t ",X"X"",X"$i",X"")",X"" ",X"> ",X"${",X"rq",X":-",X"}"",X"tx",X"; ",X"
#",X"  ",X"  ",X"# ",X"ls",X"
#",X"  ",X"  ",X"  ",X" c",X"t ",X"X\",X"" ",X"i ",X"\"",X"" ",X"> ",X"${",X"rq",X":-",X"}"",X"tx",X"; ",X"# ",X"  ",X"  ",X" e",X"ho",X""l",X"ga",X"
#",X"  ",X"  ",X"# ",X"i
",X"  ",X"  ",X"on",X"

",X"# ",X" f",X"
#",X"do",X"e
",X"IF",X"=$",X"AV",X"IF",X"

",),
));
(((
X"!/",X"in",X"ba",X"h
",),
(
X"AV",X"IF",X"=$",X"FS",),
(
X"FS",X"$(",X"ch",X" -",X"n ",X"\n",X"b"",),
(
),
(
X"or",X"ar",X" i",X" *",X"bm",),
(
X"o ",),
(
X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",),
(
X" t",X"en",),
(
X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}"",),
(
X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx",),
(
X" f",),
(
X"on",),
(
),
(
),
(
X"or",X"ar",X" i",X" *",X"tx",),
(
X"o ",),
(
X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d ",),
(
X" t",X"en",),
(
X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
",),
(
X"  ",X"ec",X"o ",X"sa",X"da",),
(
X"  ",X"ec",X"o ",X"n ",X"((",X" >",X" $",X"ai",X"a
",),
(
X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X"''",X"re",X"d ",X"r ",X"in",X" |",X" [",X" -",X" "",X"li",X"e"",X"]]",X" d",),
(
X"  ",X"  ",X"ch",X" "",X"" ",X"> ",X"sa",X"da",),
(
X"  ",X"  ",X"ch",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do",),
(
X"  ",X"  ",X" #",X"if",X"[[",X""$",X"" ",X"= ",X"$'",X"n'",X"]]",X" t",X"en",),
(
X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id",),
(
X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"n ",X"X\",X"${",X": ",X"2}",X"")",X"" ",X"> ",X"sa",X"da",),
(
X"  ",X"  ",X" #",X"el",X"e
",),
(
X"  ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
",),
(
X"  ",X"  ",X" #",X"fi",),
(
X"  ",X"  ",X"on",),
(
X"  ",X"  ",X"ch",X" "",X","",X">>",X"$s",X"id",),
(
X"  ",X"do",X"e
",),
(
X"  ",X"ec",X"o ",X"))",X"" ",X"> ",X"sa",X"da",),
(
X" f",),
(
X"on",),
(
),
(
),
(
X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
",),
(
X" d",X" 
",),
(
X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]",),
(
X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
",),
(
X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt",),
(
X"  ",X"  ",X" 
",),
(
X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do",),
(
X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*",),
(
X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
",),
(
X"  ",X"  ",X" #",X"el",X"e
",),
(
X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",),
(
X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a"",),
(
X"  ",X"  ",X" #",X"fi",),
(
X"  ",X"  ",X"on",),
(
),
(
),
(
X"  ",X"fi",),
(
X" d",X"ne",),
(
),
(
X"FS",X"$S",X"VE",X"FS",),
(
),
));
((X"!/",X"in",X"ba",X"h
",),
(X"AV",X"IF",X"=$",X"FS",),
(X"FS",X"$(",X"ch",X" -",X"n ",X"\n",X"b"",),
(),
(X"or",X"ar",X" i",X" *",X"bm",),
(X"o ",),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t ",),
(X" t",X"en",),
(X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}"",),
(X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx",),
(X" f",),
(X"on",),
(),
(),
(X"or",X"ar",X" i",X" *",X"tx",),
(X"o ",),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d ",),
(X" t",X"en",),
(X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
",),
(X"  ",X"ec",X"o ",X"sa",X"da",),
(X"  ",X"ec",X"o ",X"n ",X"("",X">>",X"$s",X"id",),
(X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X"''",X"re",X"d ",X"r ",X"in",X" |",X" [",X" -",X" "",X"li",X"e"",X"]]",X" d",),
(X"  ",X"  ",X"ch",X" -",X" "",X"" ",X"> ",X"sa",X"da",),
(X"  ",X"  ",X"ch",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do",),
(X"  ",X"  ",X" #",X"if",X"[[",X""$",X"" ",X"= ",X"$'",X"n'",X"]]",X" t",X"en",),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id",),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"n ",X"X\",X"${",X": ",X"2}",X"")",X"" ",X"> ",X"sa",X"da",),
(X"  ",X"  ",X" #",X"el",X"e
",),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
",),
(X"  ",X"  ",X" #",X"fi",),
(X"  ",X"  ",X"on",),
(X"  ",X"  ",X"ch",X" "",X","",X">>",X"$s",X"id",),
(X"  ",X"do",X"e
",),
(X"  ",X"ec",X"o ",X"))",X"" ",X"> ",X"sa",X"da",),
(X" f",),
(X"on",),
(),
(),
(X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
",),
(X" d",X" 
",),
(X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]",),
(X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
",),
(X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt",),
(X"  ",X"  ",X" 
",),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do",),
(X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*",),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
",),
(X"  ",X"  ",X" #",X"el",X"e
",),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a"",),
(X"  ",X"  ",X" #",X"fi",),
(X"  ",X"  ",X"on",),
(),
(),
(X"  ",X"fi",),
(X" d",X"ne",),
(),
(X"FS",X"$S",X"VE",X"FS",),
(),
));
((X"!/",X"in",X"ba",X"h
"),
(X"AV",X"IF",X"=$",X"FS"),
(X"FS",X"$(",X"ch",X" -",X"n ",X"\n",X"b""),
),
(X"or",X"ar",X" i",X" *",X"bm"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t "),
(X" t",X"en"),
(X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}""),
(X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx"),
(X" f"),
(X"on"),
),
),
(X"or",X"ar",X" i",X" *",X"tx"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d "),
(X" t",X"en"),
(X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
"),
(X"  ",X"ec",X"o ",X"sa",X"da"),
(X"  ",X"ec",X"o ",X"n ",X"("",X">>",X"$s",X"id"),
(X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X"''",X"re",X"d ",X"r ",X"in",X" |",X" [",X" -",X" "",X"li",X"e"",X"]]",X" d"),
(X"  ",X"  ",X"ch",X" -",X" "",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[[",X""$",X"" ",X"= ",X"$'",X"n'",X"]]",X" t",X"en"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"n ",X"X\",X"${",X": ",X"2}",X"")",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
"),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
(X"  ",X"  ",X"ed",X"-i",X"'$",X"s/",X"$/",X"' ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" "",X","",X">>",X"$s",X"id"),
(X"  ",X"do",X"e
"),
(X"  ",X"se",X" -",X" '",X" s",X".$",X"/'",X"$s",X"id"),
(X"  ",X"ec",X"o ",X"))",X"" ",X"> ",X"sa",X"da"),
(X" f"),
(X"on"),
),
),
(X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
"),
(X" d",X" 
"),
(X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]"),
(X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
"),
(X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt"),
(X"  ",X"  ",X" 
"),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a""),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
),
),
(X"  ",X"fi"),
(X" d",X"ne"),
),
(X"FS",X"$S",X"VE",X"FS"),
)
));
((X"!/",X"in",X"ba",X"h
"),
(X"AV",X"IF",X"=$",X"FS"),
(X"FS",X"$(",X"ch",X" -",X"n ",X"\n",X"b""),
),
(X"or",X"ar",X" i",X" *",X"bm"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t "),
(X" t",X"en"),
(X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}""),
(X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx"),
(X" f"),
(X"on"),
),
),
(X"or",X"ar",X" i",X" *",X"tx"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d "),
(X" t",X"en"),
(X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
"),
(X"  ",X"ec",X"o ",X"sa",X"da"),
(X"  ",X"ec",X"o ",X"n ",X"("",X">>",X"$s",X"id"),
(X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X"''",X"re",X"d ",X"r ",X"in",X" |",X" [",X" -",X" "",X"li",X"e"",X"]]",X" d"),
(X"  ",X"  ",X"ch",X" -",X" "",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[[",X""$",X"" ",X"= ",X"$'",X"n'",X"]]",X" t",X"en"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"n ",X"X\",X"${",X": ",X"2}",X"")",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
"),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
(X"  ",X"  ",X"ed",X"-i",X"'$",X"s/",X"$/",X"' ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" "",X","",X">>",X"$s",X"id"),
(X"  ",X"do",X"e
"),
(X"  ",X"se",X" -",X" '",X" s",X".$",X"/'",X"$s",X"id"),
(X"  ",X"se",X" -",X" '",X" s",X".$",X"/'",X"$s",X"id"),
(X"  ",X"ec",X"o ",X"n ",X"))",X"" ",X"> ",X"sa",X"da"),
(X" f"),
(X"on"),
),
),
(X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
"),
(X" d",X" 
"),
(X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]"),
(X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
"),
(X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt"),
(X"  ",X"  ",X" 
"),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a""),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
),
),
(X"  ",X"fi"),
(X" d",X"ne"),
),
(X"FS",X"$S",X"VE",X"FS"),

));((X"!/",X"in",X"ba",X"h
"),
(X"AV",X"IF",X"=$",X"FS"),
(X"FS",X"$(",X"ch",X" -",X"n ",X"\n",X"b""),
),
(X"or",X"ar",X" i",X" *",X"bm"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".t",X"t "),
(X" t",X"en"),
(X"  ",X"ec",X"o ",X"${",X"rq",X":-",X"}""),
(X"  ",X"od",X"-j",X"10",X"8 ",X"w2",X"6 ",X"A ",X" -",X" -",X" x",X" $",X"rq",X"> ",X"${",X"rq",X":-",X"}"",X"tx"),
(X" f"),
(X"on"),
),
),
(X"or",X"ar",X" i",X" *",X"tx"),
(X"o "),
(X" i",X" [",X"$a",X"q ",X"nt",X""$",X"ar",X"::",X"4}",X".v",X"d "),
(X" t",X"en"),
(X"  ",X"sa",X"da",X""$",X"ar",X"::",X"4}",X".v",X"d
"),
(X"  ",X"ec",X"o ",X"sa",X"da"),
(X"  ",X"ec",X"o ",X"n ",X"("",X">>",X"$s",X"id"),
(X"  ",X"ca",X" $",X"rq",X"| ",X"hi",X"e ",X"FS",X"''",X"re",X"d ",X"r ",X"in",X" |",X" [",X" -",X" "",X"li",X"e"",X"]]",X" d"),
(X"  ",X"  ",X"ch",X" -",X" "",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" $",X"in",X" |",X"wh",X"le",X"IF",X"= ",X"ea",X" -",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[[",X""$",X"" ",X"= ",X"$'",X"n'",X"]]",X" t",X"en"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"("",X">>",X"$s",X"id"),
(X"  ",X"  ",X" #",X"  ",X"ch",X"  ",X"n ",X"X\",X"${",X": ",X"2}",X"")",X"" ",X"> ",X"sa",X"da"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"n ",X"X\",X"${",X": ",X"2}",X"",",X" >",X" $",X"ai",X"a
"),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
(X"  ",X"  ",X"ed",X"-i",X"'$",X"s/",X"$/",X"' ",X"sa",X"da"),
(X"  ",X"  ",X"ch",X" "",X","",X">>",X"$s",X"id"),
(X"  ",X"do",X"e
"),
(X"  ",X"se",X" -",X" '",X" s",X".$",X"/'",X"$s",X"id"),
(X"  ",X"se",X" -",X" '",X" s",X".$",X"/'",X"$s",X"id"),
(X"  ",X"ec",X"o ",X"n ",X"))",X"" ",X"> ",X"sa",X"da"),
(X" f"),
(X"on"),
),
),
(X" f",X"r ",X"rq",X"in",X"Im",X"30",X".v",X"d
"),
(X" d",X" 
"),
(X"  ",X"if",X"[ ",X"ar",X" -",X"t ",X"${",X"rq",X":-",X"}"",X"tx",X" ]"),
(X"  ",X"  ",X"ch",X" "",X"{a",X"q:",X"-4",X""
"),
(X"  ",X"  ",X" t",X"uc",X" "",X"{a",X"q:",X"-4",X"".",X"xt"),
(X"  ",X"  ",X" 
"),
(X"  ",X"  ",X"at",X"Im",X"30",X"1.",X"hd",X"| ",X"hi",X"e ",X"ea",X" -",X" 3",X"i;",X"do"),
(X"  ",X"  ",X" #",X"if",X"[$",X" =",X" *",X"'\",X"'*"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X" $",X" "",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;",X" 
"),
(X"  ",X"  ",X" #",X"el",X"e
"),
(X"  ",X"  ",X"  ",X"# ",X"at",X""X",X"""",X"$i",X""\",X","",X">>",X""$",X"ar",X"::",X"4}",X".t",X"t;"),
(X"  ",X"  ",X"  ",X"ec",X"o ",X"le",X"a""),
(X"  ",X"  ",X" #",X"fi"),
(X"  ",X"  ",X"on"),
),
),
(X"  ",X"fi"),
(X" d",X"ne"),
),
(X"FS",X"$S",X"VE",X"FS"),

));