 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 04 00 08 05 05 0a 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 06 05 03 00 06 05 03 00 0b 05 03 05 06 05 04 05 06 06 03 04 09 05 0b 00 06 05 03 00 06 05 03 07 06 05 04 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0a 06 05 0b 07 06 05 04 03 06 09 0c 00 06 05 04 02 06 05 03 05 06 06 03 09 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 00 06 05 06 04 06 05 03 06 06 05 03 05 06 05 03 01 07 05 0a 00 06 05 03 00 06 05 03 0a 06 05 03 03 06 05 03 00 06 05 03 01 06 05 03 05 06 05 03 00 06 05 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 08 08 05 04 00 08 05 03 04 06 05 03 04 08 05 03 04 06 05 03 06 06 05 03 07 06 07 03 06 06 05 03 06 06 05 03 06 06 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 0a 06 08 06 09 06 05 0c 01 07 05 05 0b 0e 07 04 0a 06 06 07 0d 06 0c 0a 0c 0b 07 05 05 06 05 06 0d 06 05 03 00 06 09 08 00 0b 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 0a 03 00 06 05 03 09 06 05 03 00 08 06 08 09 09 05 0a 06 08 09 07 06 06 0f 08 0f 08 05 03 09 0c 08 03 06 06 05 03 08 06 05 0a 08 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 01 06 05 03 05 06 05 03 00 06 05 03 02 06 05 08 06 07 0d 0d 08 06 0b 0f 0f 06 0b 0f 07 0d 0e 11 10 06 09 09 0b 10 0d 12 14 0b 12 0e 15 19 08 0a 04 06 09 03 0d 09 05 0f 04 06 07 07 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 09 06 05 03 00 06 08 09 05 0a 05 07 08 06 0a 0a 10 09 0c 18 0c 0a 05 08 0e 0d 0f 0a 0f 06 0e 14 10 0c 14 0f 1e 19 17 12 1d 1a 0a 0a 0d 06 07 0a 07 06 0c 12 10 0c 06 0b 00 06 05 03 06 07 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 01 06 05 0d 0a 06 05 0b 10 07 0c 11 0e 07 0c 0d 0e 0b 0c 0d 18 19 12 14 10 0d 10 0c 0e 07 0b 0a 15 16 1d 14 1a 0b 15 0e 11 15 0f 10 0a 09 0e 15 07 06 0a 03 00 0a 05 03 0b 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 11 07 0e 08 05 0c 0e 0e 09 0b 11 12 0b 11 07 14 08 12 12 0f 10 11 19 14 0e 16 12 18 11 1e 1b 17 17 1e 1a 16 13 0c 18 19 18 0b 10 11 11 0b 0f 06 0d 09 03 06 0d 03 08 06 06 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 01 08 05 03 05 06 0c 04 0d 0a 05 12 0c 0a 06 0e 0e 11 10 11 14 10 18 18 14 16 09 0b 0c 1b 16 1e 16 16 1b 1a 1a 1f 17 25 16 1b 24 12 17 15 19 16 20 16 11 11 1c 06 13 0a 10 15 05 04 09 09 05 05 05 06 05 03 01 0a 05 07 02 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 04 08 07 03 0b 0b 08 11 13 0f 0f 20 12 15 18 12 13 1b 19 1b 1f 20 1c 1a 18 15 1b 1a 15 21 27 1e 22 17 1d 1b 1f 22 28 1c 1e 17 17 15 0f 16 0c 11 14 0d 16 03 09 06 05 09 09 07 05 07 08 06 05 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 03 06 05 03 00 06 05 03 00 06 05 0b 0b 06 05 08 0b 10 05 0a 14 15 0f 12 0a 09 17 10 11 18 21 1e 15 18 14 26 24 34 24 15 1a 25 29 29 29 26 3d 29 26 24 29 26 21 23 25 26 26 19 24 1f 19 15 16 14 18 10 1b 03 0e 0b 07 11 0b 06 05 08 0b 06 05 0f 07 06 05 03 00 06 05 03 01 06 05 03 04 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 05 03 00 06 0f 03 0c 06 0d 0a 03 09 05 10 0c 0e 0f 0a 0c 0d 09 18 09 1a 0c 11 1c 16 1f 22 1c 20 1a 21 20 19 1e 24 23 2c 32 2f 28 28 2c 30 26 2a 3b 36 28 2f 2b 2b 35 2e 30 28 35 2f 2a 2a 20 1c 1e 20 11 14 15 0d 15 0e 13 0f 0d 08 17 0d 0d 0b 0b 04 06 09 05 05 00 06 05 09 00 06 05 05 00 08 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 04 02 06 06 03 01 06 09 10 0f 06 05 0f 09 09 0d 0c 11 0e 12 0b 1c 10 1b 16 0f 1d 1a 2e 26 28 2c 2a 22 23 30 25 2e 36 34 27 36 39 35 3d 38 30 3d 3d 36 3a 3f 37 41 48 36 3e 45 3a 3e 30 2f 23 25 1b 16 15 14 12 12 14 14 10 0f 0c 14 12 0f 0b 0d 05 08 07 05 03 09 07 0a 04 01 06 05 03 01 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 12 05 03 03 08 07 0a 0d 0d 0e 0c 0a 07 0f 0e 0b 14 1b 1a 1f 1d 23 22 1c 22 25 2f 34 34 34 39 32 2b 30 31 36 39 46 47 45 3e 39 48 45 45 43 4c 5a 61 6b 64 6a 65 72 66 62 52 47 37 34 30 25 29 24 20 19 1b 11 1d 19 18 16 1c 14 10 11 0d 15 06 15 08 13 0e 04 0c 05 08 0a 06 05 03 07 0a 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 04 01 06 07 08 10 0d 05 0d 06 14 18 10 0f 0f 10 10 15 1b 2a 1c 21 25 26 2e 27 1f 2b 2e 3c 41 39 46 43 49 59 56 4f 58 60 6e 65 5f 63 59 5a 65 6b 87 a0 b8 b2 ab ae a9 b5 a0 81 81 74 69 4e 42 42 30 31 2c 26 2a 29 25 29 23 28 1b 27 17 13 0f 18 1e 16 14 18 15 10 0a 10 0f 0e 08 08 0a 08 0a 10 06 09 06 05 05 06 06 05 05 00 06 05 03 04 06 06 03 06 06 06 03 00 06 05 03 02 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 06 05 03 00 06 0b 12 0b 0c 18 14 11 0f 12 10 11 15 16 19 1a 1b 19 30 27 1e 27 27 28 36 35 34 41 47 4f 54 4e 68 6f 70 7c 89 9d a8 a7 a8 a1 92 9a 9c a4 dc fa ff ff ff f6 ff fd b9 94 85 86 81 70 66 55 41 41 39 3e 32 30 32 27 21 26 22 2f 2c 1b 1d 1b 1e 20 14 14 1a 16 14 0d 15 10 0a 05 03 0b 06 0e 03 05 06 0c 0a 00 06 05 04 02 06 05 03 02 0c 06 03 00 06 0d 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 02 06 05 03 00 06 0a 0c 0f 11 1a 09 0d 0d 2a 26 15 10 1d 16 15 12 13 1a 1b 2c 2b 2c 31 31 2b 31 46 4e 45 5d 6d 6a 60 63 70 74 7b a5 b7 c4 eb fe ff ff f3 f6 f9 f1 e5 f5 ff ff ff ff ff ff ff e2 bd a0 8d 7f 6f 6a 64 58 4c 45 4c 3f 41 39 34 25 25 22 25 21 24 23 1f 2a 22 1d 13 12 0d 17 19 22 19 10 12 10 0d 09 08 0c 09 0d 0f 14 0b 06 05 03 02 06 05 05 02 06 07 04 08 06 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 09 0b 0a 05 09 0c 06 08 0b 0a 15 12 05 0e 13 22 1f 19 24 14 1f 19 21 13 23 29 37 3e 33 42 39 4c 4b 55 61 5f 80 8e 9d a0 9a 90 ab c7 eb f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa cf bc a2 9b 8c 7e 76 63 55 48 48 63 5a 52 3c 2b 1e 23 22 2f 2c 2b 1c 2b 30 2a 20 1b 22 1d 1c 1e 12 11 14 12 16 0b 0d 12 0a 20 25 0d 09 05 03 08 06 05 03 04 06 06 06 0a 06 05 03 0a 06 05 03 07 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 04 06 05 06 05 06 05 03 08 0e 05 12 11 16 0f 11 13 15 1a 12 1b 1e 1c 22 1e 1d 25 23 33 44 4d 53 76 68 68 7f 7b 85 a4 c3 d1 e2 fb f5 eb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc db d1 d4 e4 d7 c9 bb 91 61 58 5f 7e 84 65 43 27 20 2b 2b 34 2e 33 34 38 3b 44 34 31 25 1c 19 20 21 18 13 19 17 16 13 11 07 0c 10 16 15 0c 10 00 08 07 05 00 0b 05 0c 05 06 08 08 0d 06 05 03 05 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 06 06 05 0a 0f 06 0b 12 0f 0a 12 17 15 19 1a 23 28 24 29 28 2e 26 22 27 32 58 78 81 94 9a a3 bd c1 c5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 db d9 e7 ed dc d0 ed cb a1 7e 70 96 9b 8b 52 49 34 3a 37 43 48 40 4d 51 45 45 4f 45 37 3b 31 2e 20 1d 23 21 25 23 15 16 0f 08 15 12 15 09 05 0a 09 08 06 0d 0d 09 16 11 06 09 07 09 0a 05 03 02 06 05 03 01 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 04 06 05 07 01 06 07 03 0b 0f 0b 0a 0c 08 0e 10 0b 0e 13 17 12 15 1f 17 11 09 16 22 38 3d 39 39 34 2b 2a 36 6e 98 b2 bd bc bb b8 b2 ba cc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc d4 a5 7b 96 b1 9b 77 6b 5f 5f 60 60 6a 57 5e 5b 55 52 52 5f 50 4a 4a 4d 49 44 41 3e 3f 39 28 25 19 23 23 1c 21 1e 12 18 10 0c 0b 0f 0d 11 0a 0d 07 0d 09 09 09 0a 0a 0c 06 05 08 0d 06 05 07 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 12 05 0e 0e 06 1c 0f 14 0a 0b 13 12 19 17 1f 18 22 21 1b 21 2a 3e 4c 46 43 46 47 3c 45 5b 7f 81 8c 8a 9c cc cb d9 e3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ce a6 a1 a7 9b 9e 93 8f 93 81 7d 75 70 6a 69 6d 67 67 62 59 5f 62 5f 62 57 54 4d 54 4f 36 2b 23 27 2c 30 2b 25 22 26 25 18 13 21 11 11 1b 0e 15 0d 09 04 09 07 0f 11 08 09 0b 01 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 04 06 06 05 03 00 06 05 03 00 09 0b 0d 09 15 12 0e 0a 13 0f 12 0f 13 14 16 18 1c 1b 18 2c 30 44 52 50 55 4b 4d 52 4e 5b 5e 69 75 7a 73 80 a6 cc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c7 b0 a4 a9 a8 9f a2 92 95 83 8f 89 7e 79 7d 77 76 6f 70 72 76 73 6f 70 65 63 65 5f 62 52 4f 47 44 42 43 44 39 33 33 2f 31 21 25 2b 1c 23 1f 1b 1c 12 10 07 0e 05 07 06 05 03 01 06 0d 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 05 03 00 06 06 12 0e 08 17 0e 15 10 11 12 11 12 16 15 21 1d 1c 26 22 25 29 32 6b 92 70 58 47 4a 57 61 5e 69 7c 81 8e 8f 94 94 9e b7 d7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 c0 b0 a0 a3 a6 9e 9a 93 96 91 94 90 91 8f 8f 8c 87 7f 81 84 82 7e 80 7d 78 73 6f 69 6d 6a 6c 63 5e 58 55 58 50 52 52 4f 44 3e 37 3a 3b 2e 2f 31 2c 24 1e 1a 11 15 11 0a 0a 0b 09 09 05 09 07 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 08 03 02 06 05 0b 09 0d 05 0a 09 11 0d 14 19 18 08 1b 18 19 25 22 20 2b 43 3e 35 39 39 62 bc f1 b0 50 4a 4e 70 8c 8a 89 99 99 9c a0 a6 a7 af d3 de f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e5 c5 a8 af a5 aa 9f a4 9e 96 9b 9d 97 94 94 9d 91 96 97 8e 8a 92 92 89 85 82 7c 7d 6a 74 6b 70 73 71 6b 6c 66 60 60 5f 5e 51 52 54 4f 4e 4b 55 50 50 35 2d 22 24 1a 1c 18 0f 0a 09 07 14 09 04 06 05 04 00 07 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 07 06 05
 03 00 06 05 03 00 06 05 03 03 09 05 0a 0e 07 0c 04 17 12 14 1b 0c 15 11 18 1c 1d 1c 24 24 2a 44 63 6a 5c 74 84 b8 d3 9f 73 6e 72 8a ab a7 b2 bc bd b0 b6 bc bb c7 d6 e4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed cd c2 b1 b8 ab b5 a5 a5 a0 a3 9d 9f 9f 96 9a 9b 98 9a 93 97 8b 8f 92 8a 8e 8b 83 86 7f 7d 75 6c 6c 6a 64 69 5b 6b 6b 69 71 62 5f 64 66 6e 6c 5f 6a 5e 50 45 48 39 36 29 18 18 10 19 0e 16 0c 0a 06 05 03 00 06 06 04 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 07 07 03 09 12 05 11 01 07 09 1f 23 24 13 1d 1f 23 20 25 26 1e 2a 24 27 30 49 86 92 98 ae c0 ba 9f 8c 8b 89 99 9b a1 ab b2 c0 c2 b5 bb c2 c9 d5 df ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 df c5 c5 c2 b9 b0 ae ad ac ae a4 a7 a9 9b 99 9f 9e a1 a1 98 9e 99 9b 9f 8c 91 8d 8a 8a 80 85 78 6a 72 71 6a 6c 69 6d 6e 70 72 67 6a 72 62 72 73 73 73 63 64 62 5b 4c 37 32 26 23 2f 1f 16 18 0a 0b 14 0b 0d 06 06 0c 05 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0c 1a 09 09 0f 0b 06 0d 1a 15 20 1d 1e 18 1a 26 24 28 27 24 29 2c 32 33 44 4c 65 89 94 a6 b5 bf b9 99 9a a0 9f a8 a6 b4 b9 be ba ca cc cd d0 d3 d8 e0 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef e6 d5 ce d4 ca c8 c4 bf bc c4 b8 bd af af ac b1 aa a7 a5 a2 a1 a5 a2 9d 9a 9e 9a 99 8c 8f 7d 80 7d 79 77 75 77 72 6e 76 77 6e 69 65 6c 73 74 6b 6d 6e 69 6d 71 7f 67 5a 48 42 34 2b 29 24 17 17 18 14 0b 0e 0f 05 09 0e 06 05 03 04 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 05 00 06 08 08 09 09 05 06 0c 06 12 1c 15 23 1b 19 20 25 1f 24 25 2c 36 3b 38 4e 4c 62 6a 76 7b 9f b3 bf c1 be b9 a1 aa a3 ab b4 bc b9 c2 c2 c9 d2 cd d5 d4 d5 e0 ed fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f0 e9 e3 e0 d6 db db d4 c6 d1 ca c4 c2 c1 b9 bc b3 ae af b0 aa aa ad a0 9b a2 a2 9a 95 8c 88 88 87 83 7e 78 82 76 6d 74 79 75 73 75 69 72 6d 69 68 6b 67 63 75 81 86 81 66 55 42 39 2c 31 27 20 1e 1d 15 14 18 0f 15 12 0d 05 09 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 06 05 08 0a 0a 08 07 0f 07 18 25 26 1b 19 24 24 20 2f 2f 3c 46 48 58 5f 64 76 84 99 ac af b2 b5 b9 bc b8 ad aa a9 b9 b1 b7 cc cd c7 ce d2 d2 ca d5 db dc ee f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 ee f0 ed ee e3 e3 e3 e0 de d8 d0 c8 c9 be be c4 c8 bb b3 bd af b0 b2 aa a5 9d 9e 98 96 8d 89 8c 92 87 85 84 7c 77 7b 7b 7d 72 6e 75 76 6a 6a 6c 67 5f 66 6d 87 8a 81 74 64 55 50 4a 3d 34 34 30 28 25 20 20 1c 18 10 05 07 06 06 10 08 0a 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 04 06 05 03 08 06 05 0f 11 08 08 0d 06 0b 11 0e 16 1b 25 37 2e 2a 2d 2d 31 41 4b 51 50 64 65 79 89 a3 b3 bf bc bc b3 ae ad b2 b5 b2 b3 b0 b8 bb bb c0 d0 d2 d1 d5 d9 dc dc df e4 e8 ed fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff f7 ef f2 f3 e8 e7 e6 e0 db e0 dc d1 d4 c7 c3 c5 c7 cb be b9 b6 ab ab a5 a8 a5 a3 99 94 a0 93 8d 8c 8d 8d 88 7b 80 7a 7c 7b 77 76 71 6d 61 63 65 63 69 78 82 82 7a 6e 67 5c 56 4d 4a 45 37 39 2b 2c 20 1c 19 15 0d 15 08 10 04 0b 0e 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 05
 0e 06 0a 0a 08 05 10 13 17 24 2e 38 37 46 3f 4d 4d 4d 54 5c 66 74 8d 9d b9 ba bd b9 b9 ac b3 b0 af ab b4 b6 b7 bc b6 c0 c2 c2 c9 da ce da db dc e6 e0 e3 eb ea f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f1 f6 ed ea f0 e2 e0 e4 e4 df d9 d4 d3 d4 d3 c9 c3 bd b7 b6 b2 ae ad ab a3 a6 9d a0 9e 9c 99 94 8e 8c 87 84 85 80 7d 7a 79 78 6d 6f 6e 67 6e 66 6e 6e 76 6c 6b 67 67 60 60 58 52 4f 41 34 2d 27 25 23 0f 16 0a 10 05 09 0c 12 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 0c 09 0b 0d 13 0a 0c 0d 11 19 2c 36 35 3a 37 38 48 49 56 5d 6b 82 9b ae c1 bc bb af b1 af b4 b9 b7 b5 b2 b2 af b7 ba c0 c0 c0 c6 cd ca cc bf c1 e2 e2 e2 ee ea ed f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f9 f4 f6 ea f2 eb dd de d5 e0 da d4 dc d8 cf ce cb c6 b8 bb b5 b1 b6 a7 ab a0 a1 a1 a0 9e 94 9d 8c 90 8c 8f 95 81 86 87 7a 7f 81 7a 73 71 71 75 73 73 6e 74 6b 6d 72 68 5d 5e 48 41 37 32 39 33 2e 20 12 0a 10 0e 06 0d 08 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 02 06 05 03 04 06 0a 07 05 06 05 03 00 0b 13 0d 10 14 11 18 26 2d 34 32 38 32 37 43 50 51 66 71 86 a2 b4 c2 c3 b6 ad a2 a7 ab b5 b0 b1 bd bd c4 be c1 c5 c1 c3 ce ca cf d6 d5 dd de e2 e3 ec f3 f4 f9 ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fa f2 f2 e5 e9 e2 e9 e4 df e6 e1 d4 db d5 d2 cc c7 bb bb b9 b2 b3 b9 aa a7 ac a3 a4 a7 a3 9d 9d 9d 9a a0 95 8f 95 98 90 7c 7d 7d 7f 75 6b 73 6f 7c 6a 6c 6e 71 69 67 65 5d 50 3f 35 40 3b 3a 37 28 20 17 0d 0f 0d 0c 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 03 03 06 05 09 00 06 0f 03 06 07 05
 17 17 19 1a 2f 38 3e 3a 37 3b 41 4d 5c 6a 7f 9a ad b2 c1 c2 a7 af a4 a2 aa aa ad b9 b9 be c3 be c7 c9 c9 c9 c9 d1 d3 d1 d7 d2 de e7 e2 e6 ed ea fa fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f9 f8 ee eb ef e9 e9 e8 dd df dc d6 d1 ce c3 c7 c2 c5 bb b8 bd ba b2 b5 b2 b4 ab b0 b1 b5 b7 a3 b2 ad a7 a3 a0 95 8b 81 7a 7f 7a 79 74 7f 77 74 75 73 69 6a 6d 69 66 61 50 47 4f 3f 3d 37 2c 21 15 18 11 15 08 05 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 07 12 0c 10 17 26 2f 3c 46 33 36 3a 42 49 5e 6d 8e a2 ac b6 b7 a8 9e a8 aa 9f a9 ab ab b2 b4 b6 c2 c6 c2 c5 cc cc c9 d1 ce db d6 d3 e0 d4 e5 e9 f1 ef f2 ff f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb f3 f6 f3 ea e9 ea e9 dd e0 d6 d4 cd d8 d0 cf c5 c9 c8 bf c2 c0 c2 be c2 c3 c3 b9 c1 bc ba b9 b5 a9 ac a3 96 92 87 85 84 7f 7e 7c 72 77 74 6f 6f 6b 68 63 65 6d 7a 75 65 5a 4f 47 3b 32 33 29 16 17 1c 07 0a 0b 09 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 08 0a 0e 09 08 16 0d 12 1b 11 25 3b 3e 38 36 41 40 4f 67 6e 92 a9 bd c0 b3 9e 9a 9c a1 9e a3 a9 ad b0 af b1 b7 c3 bb c4 cb ce cf d7 d4 d4 d5 dd db de e2 e4 ea ec ec f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f5 f8 f3 f4 ec ec f2 e9 ed e2 e5 dc d6 d2 d8 da d2 d5 d0 d4 d2 cd ca c9 ce c9 cb c7 c2 cb c7 c1 b9 b3 ae ab a7 9e 8b 86 81 86 7d 80 7e 73 73 75 73 6d 6d 68 68 65 71 7d 7d 6e 68 4d 4f 44 49 39 3b 20 1b 15 13 13 0f 0b 0c 08 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 06 09 0b 07 05 09 0e 0f 1c 18 12 27 30
 30 36 35 3a 44 4a 58 68 94 b1 bb bf ac ad 8a 93 9c 9d a4 a6 ac b1 b0 bb c5 bc bf cc cd d1 cd db db d8 e0 e1 e4 eb ed e4 f1 ef f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f8 fe f5 f8 f5 ee ec ed e5 e2 e8 e7 d9 dd d9 de de dd d9 db d8 db d0 d3 d7 cd cf cc c5 c0 b7 ba af a7 ab 9e 93 91 8f 8b 84 81 80 7a 7a 71 70 6e 6b 6a 6b 67 6a 72 71 77 7b 7f 70 5b 46 49 42 41 2e 28 13 1c 10 10 08 08 06 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 06 06 05 10 0d 0a 05 0b 0a 14 23 1d 25 2a 2f 34 3b 3e 49 5d 60 8d a6 bd c1 b3 94 94 91 96 92 9b 9e 99 a0 ab b8 bc bf c1 c9 cc ce ce d0 d2 e2 e2 dd ea e9 f4 f0 f0 f9 ff f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fa f1 f8 f7 f4 f3 ef f2 ec e6 eb e9 f1 e6 e6 e4 e5 e2 e1 d4 d1 cd d4 d5 d4 c4 c9 b9 b5 a9 b2 9e 9f 97 8d 8e 80 79 7c 7d 7c 75 80 6f 71 6e 6b 71 71 6f 72 6c 6f 77 87 7a 71 59 50 50 47 46 3b 3a 25 11 0c 0d 09 00 08 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 0a 0e 10 11 15 16 18 1f 30 33 2f 3a 34 41 51 55 61 73 9c c2 d1 c8 bd 97 8b 8b 8d 92 96 9b 9c a6 a6 ac b3 c1 bf cb c8 ce ce dc d8 e2 ea f6 f3 f6 ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff fa ff ff fc fe f5 f2 fd fa f8 f2 f5 ef f0 ea f0 e8 de eb df d7 de d9 d8 c6 cb bb b2 ab ad 9d 9d 98 96 94 8e 87 83 84 7a 76 73 78 70 76 70 6b 72 70 6b 75 70 78 79 78 70 64 62 61 4e 49 49 48 3f 31 15 1e 14 0b 08 08 09 00 07 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 06 06 0f 08 0e 06 0f 1b 1b 1e 25 28 39 3e 3f 46 51
 5b 61 74 93 b4 d4 ee e9 ce ad 87 90 90 8f 9e 96 9e a2 a7 ae b6 bb b8 c5 cc cd d3 d7 e4 df ee f6 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe ff ff ff ff fd ff ff ff f5 f0 f0 f1 e9 ec e4 e4 e2 e4 d0 cc c8 bb b8 b4 ae ae 95 9b a0 95 95 91 86 86 82 7c 79 7c 79 73 7c 71 77 6d 68 6e 7d 71 74 73 6f 6b 67 53 5d 4b 4b 4f 46 3a 21 16 0f 0d 12 0d 09 08 05 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 07 06 05 03 02 0a 0a 08 12 25 1f 25 30 36 43 45 54 55 60 80 93 a8 c8 de f7 ff f7 ce ad 91 8d 8e 93 94 a0 ac a3 a9 b0 b3 be ba c0 cd d5 db dc de e7 ee fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fe f4 eb eb ec e5 dc de d4 cf cb bd bc b9 b0 b2 9d 9e 92 92 9a 95 90 89 82 84 78 71 7c 76 77 70 72 76 77 70 6f 7b 74 6b 6d 63 63 64 5f 5c 52 4c 47 4c 37 22 19 18 10 0f 0a 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 01 09 05 03 00 06 05 05 0e 11 0d 1a 26 2c 31 26 41 4a 5c 67 6a 7a 8f a4 b6 d5 f2 ff ff ff e2 ba ab a0 96 a3 a9 ad b3 b7 b1 b5 b1 b8 be c2 c6 d5 d2 e1 e4 ec e8 f6 fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa f8 f8 ee e8 e4 e2 e2 d5 cb cf b3 bb b8 b5 b0 ad 9f a0 a1 a2 96 96 90 80 84 80 75 7d 7e 79 74 74 77 7c 72 76 70 6e 75 6b 6f 66 6d 6c 6b 6e 55 4a 45 3e 2d 28 19 1e 1d 18 10 11 05 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0a 06 10 08 0e 15 16 23 31 32 3d 3f 55 54 7d 8e 8c 9e ad
 b6 d8 f6 fe ff ef da b9 b7 c3 b8 b6 c0 bd c6 c8 cc d0 c1 c5 ba be d5 d4 d2 d5 dd e7 ef f0 fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f2 ed ed e7 de d9 dc d2 c7 c5 c5 be b8 b5 af ae aa a4 aa a2 9f 9d 8c 8c 8e 84 7f 81 81 76 81 79 7b 75 75 76 76 73 73 70 68 6e 6a 64 6d 71 61 51 40 36 2c 30 30 2b 21 1b 0e 10 16 0e 0f 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 0a 0d 07 14 14 1c 2b 29 35 32 45 4b 5f 66 79 80 92 a4 ac cf de e4 e2 d6 cc c1 be c6 c1 c3 cf d1 d6 d9 d8 dd d8 d9 cd ca d6 cd d5 e1 df e5 e9 f0 ef fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f2 ed eb de d9 cf dc cf c8 c4 bd bc bd b4 b3 ac ad a7 a2 a3 a6 9b 96 92 90 8d 81 7e 82 84 80 7f 84 79 74 6f 71 75 72 70 70 65 6d 66 6e 6e 75 75 5e 34 2c 2f 34 39 30 1d 16 16 15 0c 0a 0f 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 09 05 03 11 0a 0f 14 1d 24 28 32 2f 45 58 68 71 75 85 88 92 a8 b4 c9 c7 cf c1 be c9 ca c8 ca e4 d7 db e1 d9 da e5 ea e5 e9 df dc e0 e4 dd e1 e0 de e6 f3 f2 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f1 ed dc dc df d6 dc d8 cf c6 c0 ba bc bb b2 ac ad a4 ac 9f 9d a1 9d 9e 91 9a 94 80 89 80 8b 89 7c 7c 7f 74 6f 75 75 74 71 6c 69 68 66 60 71 85 a1 8a 58 38 35 3d 3b 40 23 1b 1a 13 1c 16 12 08 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 0a 08 13 17 1c 19 2a 2e 32 39 3e 53 65 73 87 89 85 8a 92 97 a9
 bb b6 bc c5 c5 d1 d5 d4 e1 dd e2 e3 df e7 e5 e5 f2 e5 e5 ef eb eb ee f2 ea ef f1 f9 fe f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f2 e5 e0 d7 d6 d8 cc cb c7 bf bc be b5 b3 b3 b5 af a4 a9 9e a4 a5 a9 a1 96 91 97 91 92 8f 86 85 7e 85 84 80 88 72 76 71 73 6d 70 6c 65 6f 7d a4 b2 9f 76 65 63 53 4c 43 39 25 22 23 19 14 15 15 08 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 06 09 05 06 09 11 1d 21 22 28 2b 31 32 40 50 60 75 84 83 83 8a 91 9a a0 af b5 b9 bb c5 d1 cb d1 d7 de e0 dc da d3 d0 d1 da e1 e0 e5 ee ec f5 ee f0 f4 f6 ff fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f4 ec e7 e4 d4 d6 d0 c8 ca c4 bf ba bb b1 b2 af ad ac ab 9d a3 9f 9f 9e 95 96 97 90 8f 8b 8b 87 87 83 84 83 79 7c 6b 79 6a 72 6d 76 71 6c 6a 80 a5 b3 a7 93 87 75 70 64 52 4b 35 32 23 1f 18 1e 1c 0d 0b 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 08 06 03 07 08 0d 14 22 21 26 2d 32 3d 40 4f 60 76 7f 89 8a 89 8c 8d 9c a6 aa b5 b3 b3 ba bc bd c6 ce cf cf c5 c9 c0 c5 c7 ce d3 dc e1 e4 e8 f2 f5 f8 fe ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f4 e9 e9 de df e4 d0 d3 cb c5 be c1 bb b5 b1 af af a1 a5 a6 9e 9b a0 9c 9f 9c 92 92 90 94 8f 8e 89 81 8e 85 7c 79 75 75 79 73 79 6e 67 78 6a 77 7f af ae a5 98 92 8b 84 70 63 50 3f 3b 21 1d 24 1b 1e 16 16 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 00 0c 0f 13 0f 10 12 24 25 2e 2a 35 3f 47 4f 63 6d 7d 82 81 90 91 8f 97 9b a4 9c
 a3 ac ae b0 b8 c4 c3 c9 cc cd bd be bd c1 c6 c4 ca c7 d4 df e2 ea f1 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f3 f0 ed e3 da e2 dc da d1 cf c6 c6 bd b9 b4 af af ad a7 a6 a3 9f 9c 98 98 98 90 95 9a 8c 90 8d 91 82 89 89 7c 7c 79 7c 78 71 76 68 6f 70 71 70 81 9f a5 ab a3 a7 9b 8e 80 79 6c 63 4f 42 32 25 24 1e 18 0b 0b 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 06 0b 07 0d 12 15 17 1d 25 2a 2c 38 38 49 5b 6d 6a 78 7d 87 8d 8b 8d 8f 94 93 98 9a 9f a8 a9 b3 b9 bc bd bc b8 b8 ac a7 b4 b7 bd b9 b9 c5 cf d8 e5 eb f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f0 f0 f1 ea f0 e2 de d6 d7 dd d5 ce c1 c4 c1 b8 b7 b1 b4 b0 a9 a9 a1 9d 9c 9f 9c 9c 9b 95 8d 94 8c 8e 8f 88 86 7c 7e 80 87 84 7b 76 72 7d 74 6e 74 75 8f a2 ab ab b0 a7 9c 93 8c 81 6d 5a 4e 3c 2e 30 2b 24 1f 11 05 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 04 08 05 12 12 22 2f 2a 2c 36 44 51 70 73 6b 80 80 7e 82 7c 88 82 86 8b 81 8f 92 a3 9d ad ac b0 a9 a7 a0 a8 a6 a4 a9 ab b1 b5 bc be c2 d0 cf e0 ef fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc f3 f2 ee ef eb e6 e0 e0 dd db d7 d1 c7 c3 b8 c0 b6 b3 b1 a6 aa a5 9d a1 99 a1 9c 9d 9b 9c 97 8f 97 99 8a 8f 8d 81 7c 80 86 7c 71 7a 78 74 6c 6e 68 6e 7e 96 9f a7 a3 a1 a5 9b 99 8f 75 74 55 53 45 3c 33 28 26 17 13 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 08 06 0e 18 27 30 36 43 41 50 60 71 78 82 77 73 78 7c 7c 79 7b 77 7c 7a 84 89 8c
 9b 9f 95 9c 9f 9d 96 9b 9f a6 a4 a9 b4 af bc b8 c3 bf d1 dd e4 ed fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 f1 eb ef e9 e8 e7 e0 e1 e4 e4 d5 d1 c9 bf c4 c4 ba b9 a9 ac a4 a6 a2 a5 a9 a8 a1 9b 9f 92 8e 95 98 98 97 8d 84 7f 86 83 79 81 7b 78 79 71 6d 6c 65 73 84 86 94 9d 8f 94 98 9a 9b 96 83 77 66 59 46 3b 30 2f 2f 15 0f 0c 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 0a 0e 06 08 16 20 30 32 3b 43 56 68 77 81 85 7d 79 6f 6b 73 6e 73 74 77 77 7e 84 83 88 89 8f 85 86 8e 94 94 98 9a a3 aa ac b2 bd b4 c7 c8 c8 d6 e2 e6 f4 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f3 f1 f0 f3 e4 e7 e4 f0 e4 e3 d2 d4 d2 cc c7 bf bc b9 b1 a8 ac b1 a5 ad ab a5 a7 9c 9f 97 9f 99 93 96 91 92 94 88 88 8a 7c 7a 80 73 7c 6d 6e 77 6f 74 70 7d 89 83 88 84 87 96 a0 a2 9d 88 7d 63 59 4d 39 34 2e 2c 1f 0b 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 08 0a 0c 0d 1d 23 2d 31 3b 4b 61 79 7e 81 7c 73 6e 69 6c 67 6b 6d 6f 70 7b 80 77 72 81 80 82 85 83 89 93 8d 9c a0 9c ab a7 ad b8 b8 c1 cc cd df df e9 f1 fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff fb f4 f3 ed ed ed e4 ea e3 e5 ed dd dd d2 d0 cd c5 c7 ba b8 b0 b1 ac af a4 ae a3 a7 9e 99 9c 9d 9c 97 98 9a 97 92 8e 87 81 7e 79 7f 75 76 6e 71 67 76 73 7b 77 7f 7c 76 72 76 8b a0 ab aa 91 7f 75 6b 5a 50 3f 31 2c 26 1e 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 06 0b 09 05 16 13 24 37 2c 39 44 49 64 6b 7c 82 6f 74 61 53 62 6a 6e 6d 6e 74 75 77 79 78 7f
 80 83 83 84 97 8e 95 9c 9a a7 aa ac b9 c1 c2 d3 d2 d8 e2 e3 f1 fb fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fa fc f6 fb ef f3 eb f0 ef ef f3 f5 e1 e8 dd d2 d1 d6 d1 c4 c3 c1 bd b5 b0 b5 b9 a6 ad aa a7 a2 a4 a6 98 9a 99 98 92 8a 8e 81 84 76 78 6c 71 73 6f 71 70 74 73 78 79 6f 6c 79 6f 7f 9d b9 b3 9b 99 89 77 6c 56 45 31 2c 2a 1e 09 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 06 0c 0e 12 16 21 28 2b 2d 2d 42 4f 70 74 84 75 6e 68 58 5e 62 6a 69 6a 6e 72 76 73 7b 70 86 86 84 83 84 91 8d 97 92 a2 a5 b0 ad c0 c2 ca d3 da dd e7 ec f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa ff fa f3 f5 f6 f5 f7 f9 f2 ef fb e9 ea e9 dd d8 d7 d1 cf cf ba ba bd b3 b6 af b9 ad a9 ab a9 a3 a0 a8 9f 90 97 91 8c 8e 81 78 79 7d 7d 7c 74 7b 76 75 76 75 6f 74 70 6d 69 72 7b a0 b9 bb aa 91 8a 85 6f 5f 51 3c 36 2a 22 0c 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 0f 09 0c 14 21 25 26 33 45 4c 5f 65 7d 80 7d 7a 5f 5d 5a 61 6e 66 70 6e 6c 75 71 7d 7a 7a 83 83 80 8a 92 95 90 9c a1 a3 a3 b1 b9 bd c8 cc e0 dd de e4 ee fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fd fe f9 ff fb f0 fd fa f1 ee ea ee d9 e5 db d2 cc cb cb c5 bf c2 bb b8 b7 b0 b6 ae a4 a0 a2 9f a9 97 93 8f 85 8b 85 84 7f 81 7e 78 7e 7d 7d 78 7b 6d 6d 72 6c 6d 67 77 7f 96 ab b9 aa 9f 90 81 76 67 53 47 3a 35 1b 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0f 0f 0e 10 0f 22 2d 2d 44 41 62 72 78 8c 96 87 75 63 67 66 64 6a 64 73 71 71 6f 6b 7c 79 84 89
 8e 8e 8d 90 9c 9c a3 9f ac b0 b1 cb cb c5 d8 df e2 e7 f0 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f6 ff f5 f8 f0 f2 ed e2 e4 dd d4 ca ce c1 cc c2 c0 bc c0 c2 bb b5 b6 ab aa a2 9a a1 91 96 86 80 8a 87 86 7e 8a 81 8a 82 7e 79 80 73 6c 71 68 5f 64 6d 6e 7d 7b 96 a9 b3 ab 98 96 7f 6a 5c 4d 3f 31 1e 14 05 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 06 06 05 06 09 0f 18 16 2b 2d 2b 39 3d 52 72 7a 8c 98 95 78 68 66 6a 6f 70 6d 77 76 71 7c 7e 7f 7d 89 7e 87 90 89 8b a0 9b a3 b1 b7 ab c2 c6 ce cd d9 d8 e2 ed ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fd f8 f5 e9 f2 e8 e1 e7 dc dd da c9 cf c3 c5 c1 c6 c5 b4 bb b3 b2 ab a0 a7 a8 a2 9e 95 94 85 8d 88 92 97 85 89 8b 7e 7d 78 78 72 6f 6c 74 60 65 6e 6d 70 7e 7e a5 a4 a0 a3 90 82 79 62 54 46 3b 2d 1c 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0d 0d 14 0f 1e 25 2b 27 37 40 51 69 7c 7d 90 8b 7c 72 69 62 6d 78 75 75 75 76 77 7e 7c 8b 88 86 8e 8c 91 94 a3 a6 a9 b5 b7 b4 bd c8 d0 d9 db e2 e1 f5 f2 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff f6 ff fd f0 f7 eb e2 e5 dd df d7 ce ce c6 c8 cb c6 bc bd c0 b9 ae aa a5 a5 9e 9d 9e 96 9a 93 94 8d 93 8b 8f 89 81 78 72 6e 74 69 6f 63 64 61 66 76 79 73 70 72 87 98 9f a6 8b 85 72 6b 50 38 36 26 1a 09 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 09 14 1e 17 24 32 2e 31 32 42 53 69 74 82 81 7c 74 70 73 6d 6a 72 74 7d 7d 81 82 84 84 86 8e 89
 94 90 96 a1 a1 a8 aa b4 b2 bf c8 d1 dc de e9 e3 f5 f5 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f4 f4 f6 ee e8 e5 e4 e0 d6 d1 d6 ce ca ca c2 bc bc bf b3 b6 b0 a9 a7 aa a6 a0 a0 9c 92 98 93 8e 92 89 80 84 7e 74 6f 71 64 69 68 6a 6d 72 75 75 70 62 68 73 8a 9c 99 98 85 7f 67 57 4d 38 2e 25 10 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 09 09 06 0b 0d 12 18 24 2d 2f 2a 39 46 48 55 6f 73 7e 7b 75 6c 76 75 6d 6c 79 7a 7e 7b 7f 7e 7d 83 8d 94 95 93 94 9a a9 ae aa b1 bb c4 c5 c6 ce d7 e0 ee e8 f4 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff fc ff f6 eb ee e7 e8 e4 e8 d3 d9 d6 c9 c4 c8 bc c1 b7 b2 ae af b5 ab af a5 a5 a3 a1 9a 9d 98 91 94 90 90 80 83 79 78 70 70 69 6b 6b 6a 6a 79 7a 75 6a 6c 64 71 75 92 90 9b 96 77 71 56 4f 4a 38 2e 1e 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0e 0a 0a 18 17 1e 2e 36 39 35 40 45 51 59 62 6e 72 76 70 6e 77 73 77 76 70 73 80 78 80 88 89 8c 8b 8b 8d a0 97 a3 a5 b4 a9 b9 bf c5 d2 d6 d9 df df e6 f6 f3 f9 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fc fc ff fc f9 fc f5 f0 ed e1 e6 df da d5 d1 cf ce c5 ca ba c4 b8 b2 b9 b6 ad ad ad a9 a4 a4 a4 a5 a1 9b 95 8e 8a 89 85 7f 75 77 6e 6d 6f 67 71 75 76 75 65 69 6c 66 63 67 61 72 7f 99 8d 82 76 66 5d 50 38 30 1e 11 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 09 03 06 08 03 07 0a 11 12 1d 28 3a 4b 59 5e 5c 52 59 68 71 73 6d 71 6f 6e 6f 6f 70 7c 78 85 83 86 85 8f 8e 8a 94 97 92
 98 9f a5 ab a8 be b4 c2 ca d0 d1 de db e5 ea ee f0 f3 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 ff fa f7 f2 f9 f4 ee ed e7 e0 da d8 d7 d0 d0 c8 c5 bc c1 ba b8 b9 ba b6 b1 ab b2 a5 a9 9f 98 98 92 98 8d 8c 85 89 83 7b 6c 6f 6d 70 75 76 7b 7b 78 76 76 6a 6c 64 63 5b 64 65 75 88 8d 7f 7f 68 5c 4f 3f 35 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 08 05 0f 06 06 19 1e 2a 39 43 54 65 79 7f 7b 76 7d 78 73 6b 68 69 6c 74 75 78 72 7a 7c 87 89 8a 8f 92 94 99 9e 9b 9f 9f ad a7 ba b5 be c5 d2 d0 da e0 e8 e2 e5 f2 f3 fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fc f3 f6 f9 ed fc ee e7 ed e6 e0 de dc d2 d4 d2 c3 cb bd b7 bd bb b8 bb ac b3 ad b2 a4 a8 a0 a3 9c 9a 94 92 84 80 84 73 7c 76 79 71 67 7a 7c 83 7d 79 79 73 6c 6f 60 5c 65 62 5e 6b 7b 87 85 7f 6f 59 58 41 31 21 0d 09 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 02 09 1c 23 41 53 5c 6b 6f 80 84 92 9b 8b 75 69 6d 69 67 69 65 6b 78 75 7a 87 84 89 85 8e 95 8e 95 a0 a5 a9 a6 ae ba c0 bd cc c9 d0 de d5 e3 ec f0 f5 f7 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd ff fc fe ff ff ff fc f5 ed ea f0 f8 e3 e9 e6 df df e0 d7 d3 d5 c9 cd c6 c2 bf bd c1 b5 bb b2 ac a6 a1 a0 a4 99 97 97 87 92 84 82 84 80 7d 80 6f 7f 82 7a 80 7b 7d 7c 78 7b 73 74 62 6e 62 5f 62 64 61 64 7c 89 85 70 66 59 4b 3d 1a 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 0f 12 1f 37 43 5b 62 70 80 86 8f 99 9d 92 75 62 5d 69 71 67 71 76 6d 7d 74 87 86 88 90 8b 9a 9d 9f 9d a9
 a9 aa b5 b6 bf c5 c5 cb d2 d0 db e4 ea f3 f8 fb fe f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fc f8 f5 fb f3 fc f9 ff ff fe fb f4 f3 e4 f2 e2 e3 e7 d8 e0 db d3 d5 d2 c9 cd c5 c5 be ba bb af ac ae ab a4 a4 a4 a0 96 8e 8c 88 8a 8d 81 85 81 7a 77 80 7c 7b 7a 7e 79 75 7a 79 6f 73 73 6a 63 61 62 63 5f 59 5c 6a 87 82 72 61 5b 3f 36 23 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 07 08 0e 18 2d 44 54 66 74 74 80 8c 98 9e a6 8d 67 68 66 65 6c 74 77 7b 81 83 82 8c 81 8d 93 9b 9d a3 a0 a9 ab b2 b8 b5 be c6 c2 ca cf d0 d6 de df e9 ea f1 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff fc fb f9 fb fe f9 f6 fe ff ff f5 ef ec e8 e4 eb e6 e4 de de d5 d4 de d9 ce d1 c8 c3 bb b7 ba af b1 ae aa a3 a5 98 9e 95 95 95 8c 90 82 84 7c 84 82 84 85 82 82 80 7d 7f 7c 80 7d 74 74 74 6f 68 61 62 5f 5f 61 69 63 85 88 79 67 5f 4d 35 1a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 04 06 05 07 16 19 43 49 58 74 79 7e 8c 96 9a ac a1 7c 68 62 64 64 6b 70 73 80 7c 85 89 85 8a 96 9a 9b a8 a1 a6 a9 ac b9 bb be c1 c3 c8 c9 c4 cc d8 d7 e1 e5 f0 f1 fb fb f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb fe f9 fb f8 f0 f5 f1 f8 fb f9 fc ff ff fe f2 eb e9 f0 e6 e2 e3 dd dd df d5 dd d0 ce cc c4 c0 be ba b8 ae ae b1 a1 9d 9e 9c 9c 90 91 8f 8d 8e 8f 89 88 84 85 84 85 84 87 87 7b 84 87 85 85 81 6f 72 73 6d 64 65 62 60 59 56 65 78 85 75 70 5b 43 34 18 06 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 12 14 28 3a 59 62 6b 77 85 95 97 a3 a6 91 72 60 68 65 72 6f 6d 7a 82 81 8e 8b 8b 97 9a 99 9d a5 aa ab ae b0
 be b8 c2 bd bc c9 c5 cf d6 d8 df e5 ed e9 f2 f7 f7 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 fb fb f8 f9 f4 f5 f3 f5 f0 f2 ef fe ff fd f0 f1 e9 e7 df e0 db d1 d6 d3 cf e0 d6 c9 ca c2 be b6 b5 b7 ab a8 a5 9c 9e 96 98 a0 9a 96 91 85 89 8f 88 8f 8a 88 8c 83 8b 7e 84 89 8a 86 78 83 80 77 6e 73 6b 64 5d 5d 5f 5f 64 6a 75 8a 80 63 54 46 2d 1b 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 0c 09 0e 1a 2e 44 62 70 79 89 92 9a 9f a6 a2 83 70 63 68 6d 6b 73 72 75 80 7e 8c 90 8f 96 a1 9e a5 b1 a9 b4 ba b6 ba ba c0 c3 c3 c4 cd d0 d3 d4 e1 e5 e4 eb eb f4 ff f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f7 f8 f6 f6 ed f8 f8 f1 f1 f0 ea ec f6 f4 f9 e9 dc e7 e8 dc e3 d6 d3 cc d0 d4 cc d1 cc c2 c0 bd b9 b2 b3 9f a4 a6 9a 9e 9e 94 9b 91 97 95 8e 92 8d 8e 8f 8c 88 8c 86 83 89 84 89 81 7b 88 79 7a 76 79 78 67 6a 64 62 64 67 60 6e 73 85 7c 66 57 44 2b 1b 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 04 02 0a 05 10 1a 2c 4d 61 75 88 8c 99 a2 a7 a7 a0 7f 6b 62 6b 6f 72 75 79 7e 83 8e 92 99 8f 97 97 9e a6 ae b2 b3 b4 b8 c2 bc c1 c0 c6 c5 ca d0 d5 da dd e4 e7 f1 f1 f1 f5 f0 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef fa ec e3 e8 eb ea f0 eb ef eb ed ea ea e6 df e3 da d6 d4 d3 cf ce c6 c5 c6 c6 c7 c0 b7 ba ae b1 b1 ac b2 a2 9b 9b a2 97 a2 99 98 97 9b 95 98 8f 92 8f 93 88 8b 8b 7d 80 85 79 7f 85 7a 77 75 71 68 66 68 65 6a 65 64 64 76 8b 7a 66 59 41 2a 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 07 01 06 06 10 1f 2b 4d 65 72 8d 90 a0 a6 aa ac 92 73 67 67 67 6f 78 76 7f 89 84 8c 91 98 9b 9a 9d a5 aa ac ac a9 b4 a9
 bc bb b5 c1 c5 c7 d0 cf cf d9 d9 d7 e0 e6 ea ee f9 f8 f7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 fa fa f6 f7 f6 f1 f0 e7 e7 eb e6 e8 e9 e7 e1 e3 e0 e0 e9 dd e0 d3 d2 d1 cd cb cd c0 bf bd bd c1 be b8 ba b4 ad b0 a4 a4 a2 a0 a5 91 98 96 9f 9d 98 9b 98 8e 90 95 95 91 8f 85 88 82 81 83 83 7b 73 73 77 6e 71 6b 6a 68 61 5e 66 5a 67 78 85 7b 64 57 3a 2f 14 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 0f 06 08 11 22 3a 58 67 71 87 a0 ab b6 b5 a1 80 6f 6a 6d 6e 7a 79 7d 79 89 85 8e 8b 97 9c 9f a3 a4 a8 aa aa b2 c0 bb bc b8 bc bb c4 c4 c3 ca d0 d0 d4 e0 e2 e1 ea f1 f5 fb f3 fe f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f3 f5 f1 ea e9 f6 ef ed e4 e3 e2 df e7 e6 e1 e6 de da d5 d2 dc d0 cb ca c9 c4 c0 bb c3 bc b8 bd b9 c2 b6 bf b6 ae b0 a5 a8 a8 a7 a5 a7 97 9e 9d 9a 9d 96 9a 9d 96 91 93 94 8a 7f 84 7c 7c 7e 7a 71 7b 76 7b 6f 6d 64 6b 5f 69 64 63 6d 85 85 76 67 4e 40 2e 17 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 04 06 05 06 00 0d 09 15 2a 43 5b 65 7e 8f 9c af bd af 9b 78 70 6c 65 6e 75 79 83 89 8a 92 94 98 9d a7 a5 a3 a6 b0 ae a9 b8 b6 b3 b3 b9 bf bf c4 c4 cd d3 d0 d1 dc dc de e1 e9 eb f0 f9 fd fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 fb f5 f5 ee ec e8 e8 f1 ed ec e3 e7 de e4 e5 de e4 dd db e1 d9 cf dc db cf c8 cd c7 c4 bc b8 ba bc bc b6 b7 b6 b6 b5 b0 b6 b5 b3 a6 b1 a7 a5 a6 a8 a6 a5 aa 9e 9d 9f 9d 94 93 8a 83 86 85 7b 7b 79 82 7d 7b 7a 7d 75 72 70 6f 6f 69 63 67 66 7c 80 87 79 67 59 36 27 16 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0d 0a 06 0b 15 2f 40 5e 77 86 98 a6 b9 b5 ab 81 6e 6f 6e 69 75 74 7c 86 8b 89 94 97 91 96 a6 a3 aa ab ad b2 b4 b1 ba b9
 c3 bb bb c3 c4 c3 c2 cc cd d7 db e4 df e7 e6 ee f3 f0 f3 fa ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f5 ec ec f5 e8 e8 e5 dc ea ec ed dd e0 e8 da e4 d2 d9 d9 d7 d6 d8 d3 d5 d4 ca ca c5 c8 c7 bd be c0 bd bd b7 b7 b9 b5 b2 ae aa af a8 a5 a5 ac ad a3 a6 a7 a6 a7 9a a1 95 93 8d 8b 8e 80 84 77 7d 7e 81 78 7d 78 7a 79 75 75 71 69 72 67 67 66 67 74 82 97 7b 62 59 38 25 12 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 08 00 0d 10 11 2a 3e 5e 7d 87 9e b5 bf c2 a5 7f 76 6f 6c 76 78 79 81 84 8f 93 94 9b a0 9e a6 a5 ab a9 af c2 b0 b6 bc b5 bc b9 bd c0 c4 c4 ce d1 d6 d1 db d6 e2 df e8 ee ec ef f2 f8 ff fd fd f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 fd fb f4 f7 ec f5 e8 ec e3 e3 e0 e4 e7 e0 dc e0 dc df db e1 dd d5 dc d5 ce d0 d2 d4 d2 c8 ce bc c1 c4 b9 ba b6 c0 ba bd bb bd b7 ad b0 a4 ae af af ae b2 af a3 b5 a0 ab 9c 9f 9e 96 9b 8a 87 84 85 81 7d 77 7b 71 78 7a 76 78 80 80 6f 6b 69 65 64 68 62 68 7a 8f 8c 79 6c 54 36 21 03 01 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 00 06 05 04 0b 07 08 15 1f 3d 65 83 92 ab bb c2 bb 99 74 76 75 77 79 7b 80 85 89 89 8f 95 9d 9f 9a a2 a4 aa ab ad bc b3 b1 b9 bc be ba c4 c6 c0 c6 c6 d3 df d3 d5 d7 db d8 e8 ec f3 ef f1 f6 f7 f1 fa ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe f6 ff f3 f2 f3 e6 e8 ea ec e6 e6 e2 e1 de de da d8 e2 db d0 d4 d4 d4 cd cb cf c2 c5 ca c4 d0 c1 bc c2 c1 b9 b7 bd b6 b3 b8 b6 af b7 b6 b0 af a6 af a6 a7 a9 a0 a5 a8 a3 a8 a8 99 a2 92 8f 8f 92 8d 84 79 80 7e 7e 7f 75 77 7b 7b 77 7b 7c 7b 6e 6a 6d 61 70 69 6d 85 8e 97 83 65 58 33 19 07 05 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 08 06 17 19 1c 35 54 79 98 b2 c4 c7 bb 92 80 7b 78 78 7b 81 8a 89 8d 95 92 94 9a 9b a4 a6 a5 a9 b1 af b9 b4 b8 ba c2
 be bb c2 c2 c0 ce ce c9 d4 d3 d9 d8 df df e0 e4 e5 e4 f3 f4 f2 f3 f3 f5 ff fe ff fd ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fc f6 ff f7 f0 f7 f0 e9 e8 e7 de de e1 dc db d6 de db d8 d1 d4 d2 d1 ce d1 ce cd c6 c6 c7 c5 c7 c7 c3 c4 c6 bd b1 ba b5 ba bb b5 ae b7 a6 b0 a6 ad b3 a5 a0 9d 9d a1 9c 9a a2 9f 9e 9c 98 91 90 8d 8a 86 8c 7f 83 7c 7c 79 80 7a 76 7e 79 76 78 6f 71 70 6f 6d 68 6a 6c 70 7b 93 8e 76 5c 47 23 1c 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 06 08 06 10 10 15 34 52 76 9d b6 ca cd b4 8b 7a 7c 7e 77 7f 84 83 8b 91 93 94 9c 9b 97 a1 a4 a8 a8 a8 aa b3 be b0 bb c2 bf bc c4 c4 c4 c8 d2 c6 d0 ce d8 db d6 e2 e5 e3 e6 e9 ed f2 f3 ef f6 f8 fe ef fc ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f9 fd f8 fc f4 ec e9 e0 ea df de df db db e2 d3 d5 d0 cf d1 d2 d1 cd c9 c7 c3 c5 cc c2 c5 c0 c0 bd c4 c4 ba bb bf b4 b2 b6 b4 ab ab b0 ab ae a6 a4 a6 a6 9e a3 a0 99 97 97 95 97 95 94 8e 94 92 8c 89 86 89 82 84 83 7c 73 7b 7a 75 79 75 6c 72 73 7c 73 61 6e 68 6b 6c 60 6e 8d 8a 92 7a 60 4a 21 14 07 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 06 05 03 08 10 07 16 19 2a 51 6f 98 b7 d2 d0 b2 88 7f 74 85 83 85 8b 8c 8e 93 97 98 98 a1 a4 9f a1 a5 af af ad b1 bc bb c7 cb c8 c5 c2 c7 cc c9 c2 ce ce d2 d7 dc da de e2 e4 ec ed e2 e9 ec f1 f2 f3 fa f6 f7 fb fd f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fe f4 f8 ed ee f5 e8 dc de dc dc db da d3 e0 ca ce d5 d4 cf c7 cf c1 c0 c6 c3 c5 c2 c5 bb be be b1 b8 b7 b6 b9 bd b5 bc ad ad b2 b3 ae af b1 a7 a7 a3 a3 a7 9f a1 94 9d 99 a2 a0 93 99 8f 96 91 94 93 92 8b 8b 74 83 79 7a 7f 7a 77 7c 7a 79 79 74 75 77 71 6c 6e 75 6f 6f 66 73 92 9b 91 77 57 3d 1b 09 03 03 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 02 06 10 18 24 2c 4f 74 9c bd ce c6 aa 84 85 83 81 85 89 88 90 8c 96 9d 98 9e 9a a0 9f 9a a5 ac a6 b2 bf ba c1 c3 c9
 ca cb cb c8 ca c7 c6 cd d3 d6 d9 d5 db dc dc de de e3 e4 eb ec ec f0 ee ed f4 f1 f0 f9 f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fc f2 f5 eb ee ef e4 e4 e2 db e3 d5 d6 d0 d1 d3 cd ce c8 ce bf c7 c2 c2 c2 c3 bf c3 c1 c2 b8 b2 b6 a7 b5 bb b9 b0 b7 b4 b4 ab b6 a9 ad a7 aa a3 aa aa a0 a9 a0 9c a1 9b 95 9b 95 96 97 9e 95 92 92 96 92 8f 8c 8f 86 87 7c 81 7b 7e 7f 75 7c 7f 7e 81 7c 76 77 6e 6e 73 6b 6a 6f 86 94 94 8b 75 5d 3c 19 0f 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 15 0d 15 13 2d 4c 6e 9c c0 d0 c7 99 7f 7a 85 81 87 90 86 8a 8d 8e 98 95 93 9c 9b 9c a7 a5 a9 a5 a4 b0 b1 ba be c4 c0 be c2 c5 c7 c9 ca ca c1 c9 ca d5 ca d5 e1 d9 de df de e5 e4 e5 e9 ea ee e9 f5 f3 f7 fb fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 ed eb eb e6 e6 e4 e2 d9 db d2 d1 d1 cc cf cf c4 c8 c9 c5 c9 c6 bb bd be c1 c2 b4 ba b4 bc b6 af a6 ac ad b1 b0 b0 b5 a7 a5 a4 b0 ad a4 a2 97 a0 a2 a3 a5 9f 9d a1 92 96 90 9b 9b 97 9e 92 9a 94 8b 91 87 88 8b 88 87 86 80 7e 7f 78 72 7f 78 83 76 82 78 7b 6c 6e 69 6a 74 6e 83 92 97 8b 75 4d 29 23 0e 0c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 08 05 08 0b 07 0b 10 1f 2d 57 75 a0 c3 d5 bb 97 86 84 81 8f 85 87 87 93 8f 9a 93 9c 9c 9e 9d 9b a0 a0 ae ac a9 b6 b3 bc bc bc c8 c5 bf c4 c5 c9 cb ce cc d3 cc cf d2 d2 db d9 e3 e0 d6 e3 e1 df e5 e7 ec e9 e8 f4 f6 f8 f9 fe ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f7 ee ef ee ec eb de e0 d4 d6 d0 d9 d5 d0 d2 c8 c0 d2 c4 c9 ca ca cc bb c2 c3 b9 b9 bb be bd b8 ba b2 ae ae b0 bb b0 ac b1 a3 a8 ab ad a5 ab a9 a4 a1 a1 a1 9d 99 95 98 9c 97 98 9b 99 94 94 96 95 97 95 95 87 89 86 86 87 85 81 7c 7e 7f 7e 7f 84 86 81 85 7e 75 6f 71 6e 70 6a 6e 86 9b 9f 92 75 58 38 1f 10 09 07 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 09 0b 14 11 23 25 4a 7f 9a bf d0 b6 9e 85 84 83 86 8f 84 86 8f 96 95 a0 9b 9a a5 9b 9e a1 a5 ac a6 b1 b5 ac b8 bf b7
 c4 c5 c3 c5 c8 c5 c9 c9 c7 d5 c9 ce d3 db d6 dc d5 df d6 dd dd e1 e4 e4 eb e3 e8 ed ea eb f6 ff f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f1 eb ed ee eb e7 db e6 da dd da d6 d1 d6 ca d1 cc c7 c5 ca c6 cb cb c5 be bc c4 bf ba b5 b7 b8 b8 b7 b2 b4 af b2 b3 a7 ad ad 9e a4 a6 a6 a7 a7 a0 a5 a2 9f a1 9e 9f 9d 97 9a 95 93 9c 92 92 92 96 a2 94 8b 8e 8d 8f 8d 85 85 85 7c 7a 84 83 81 84 83 80 82 80 7d 7e 7a 75 6f 73 6e 75 82 a4 93 94 70 55 3a 26 12 09 02 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 0a 0e 10 18 14 2c 48 7c 9a c4 d4 b1 96 85 83 8c 87 8d 85 89 88 8b 99 9c 9b 9e 9b 9d 9f 9b a2 9e a4 aa a5 ad a6 b5 b1 bb bd c6 c0 bd c1 c8 c7 d0 d4 ca ce d6 d0 d6 d4 d0 d8 d5 d6 d0 db dd e3 e1 e0 e5 e4 e3 e7 f2 f0 fb fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f6 e5 eb e1 e8 e8 e5 dc dd d4 d3 d3 d1 c7 c6 cd c5 c4 c7 be bf c2 bd c0 c0 b9 be c1 bb b4 b3 af ab ae ae b2 af b2 af a6 ad a3 a3 a6 a2 9a a3 9c a1 a2 a3 96 93 8f a2 96 97 9b 8f 92 92 90 97 97 99 98 99 8a 89 87 84 90 86 85 8f 7d 82 85 7d 7f 83 81 84 89 80 8e 80 7f 7a 76 7b 68 6b 76 84 97 98 95 74 5f 44 27 1c 16 00 06 07 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 04 0a 0c 0b 15 20 32 51 76 9e bf cf b7 91 89 83 8e 8b 8c 8d 8c 8a 8e 8e 98 96 98 a0 98 a0 a2 a5 ad ac ae ad a8 ac ae b3 b3 b4 b7 bd c0 c9 c8 ca c5 c7 cc cb cb cf cf c9 cd cf d8 db d3 d8 dd d5 e9 df e4 e6 e6 e6 e5 ee ee f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f9 f5 ef e2 e4 e4 e0 dc d7 de db d0 cb c8 cb c7 ce c4 c1 b6 c4 c7 b9 bb bd b8 b3 aa b3 aa b2 ad af ab a7 a7 aa ad 9e a5 ab a6 a1 a7 9e 96 9e a6 9b a7 a9 9e 9b 94 98 9f 91 92 8c 8b 8e 91 93 96 94 8a 91 97 96 95 8b 93 84 8c 86 8d 86 81 86 85 8c 86 8a 7d 7f 85 8b 88 81 7d 75 7a 73 6b 6f 6a 85 9f 9e 97 78 62 4e 31 22 0c 00 07 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 05 06 09 04 04 0c 15 17 25 3a 59 74 a9 c7 d3 b3 94 94 87 8a 90 8c 8c 8c 90 95 9a 9a 95 9e 9c 9b 9f a1 a5 a5 aa b0 ab b4 a6 ae b4
 b2 b4 b9 be c7 b8 c7 c2 c8 c7 cb ca c8 d2 c4 cc cc cf d9 cf d2 dd dd d4 dd de dc de e3 ec e5 f0 f0 f0 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 f6 fb f0 ec e0 e3 e2 db dd db d8 d5 cc c5 ce d0 c8 c6 bf c3 be bf bf bb b7 b5 b7 ae b3 aa ac a8 a9 a5 a3 a4 a2 a0 9d 9f 9f a6 a7 ad a6 a6 9e 98 a1 9c a6 a0 96 9b 96 9e 9a 99 96 90 92 91 8f 8c 91 94 86 9e 91 93 93 92 86 8d 89 8f 86 88 85 87 81 7c 7f 85 84 87 86 81 89 7d 7c 75 73 70 6f 68 73 85 a3 a1 8d 84 69 51 36 25 15 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 05 03 02 07 0d 15 22 3e 52 79 a9 c1 cb aa 8f 8b 8c 8b 8c 89 85 7f 84 90 96 a0 99 97 97 99 9c 9d a2 a3 a0 ae a9 a3 af a8 ac b1 b2 bb b6 b7 bd be c3 cf c5 cf c9 c7 c4 c1 cf c3 cd cb cc ca d4 d6 cf d5 d3 da db e7 e0 de e6 ef ef f6 f4 ff f7 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f5 f7 fc f6 eb e8 e0 df da d6 d3 d1 c9 d1 cb c5 c5 bd c5 c5 c4 bd ba bc b9 b3 b5 b4 b5 b0 ae 9f a2 a7 a5 9e 94 99 96 8e 8d 96 8f 98 9a 97 95 9f 96 97 99 97 9d 9f a0 9e 99 91 9a 8c 90 90 8a 8a 8b 8f 8f 87 91 8f 95 95 88 90 83 8f 8d 86 91 82 7e 81 82 84 84 83 8b 8b 8a 85 81 84 7c 76 70 70 6b 69 71 7f 9f a2 a1 86 66 51 31 25 1a 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 07 0f 10 1f 29 47 65 84 af c7 c9 a7 93 90 8b 8d 90 88 94 87 8b 90 92 95 91 9e 9b 9b 9e a4 a6 a6 a0 a8 a7 a7 ab ad a7 af af b2 ae bc bf b8 be c4 c5 c9 c6 c0 c6 c2 c6 c4 c5 ca ca cb cf d6 d5 cf cf d4 d8 d3 d8 e1 e9 ed ed f3 f7 f6 f8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fd ff ff ff ff ff ff ff ff fd f4 f2 ef ee ee e7 e6 d9 dc d0 d8 d2 cd c9 c5 c4 c9 bf c1 ba bf bb bb b7 b7 b7 b3 b4 b0 a8 ab a3 9c a0 9b 99 9c 91 90 96 8d 8e 8e 90 92 97 8b 8e 9a 93 8e 95 94 9c 9b 95 9c 8e 95 8a 90 8b 87 8e 8a 87 89 8d 8b 8c 8b 89 8a 8d 8e 8b 8c 91 8a 89 82 83 7f 7e 80 84 89 83 89 83 7e 85 81 7c 70 77 68 62 6c 6a 85 9c a9 a3 94 78 5b 44 2d 1d 09 06 06 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 09 06 0d 06 09 27 30 44 6b 90 aa d0 c2 a0 94 8f 8b 91 90 8a 8b 92 91 95 97 97 91 9d 9b 9b 93 a1 a4 a1 a3 a4 a9 a6 a0 ab ac
 ac b4 b1 b0 bb b5 bb c5 bd c8 c8 c3 c6 cb cf cb c7 c2 cb c7 cc c7 c7 cb cc cc d5 d1 cc db d7 e2 e5 e0 eb ef ee f4 f7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 eb d5 db cd ec ff ff ff ff ff ff fb f8 ef f0 eb e0 e4 d9 db d0 dc cb d4 d1 c2 cc c2 c4 bc c1 bc b9 bd b6 af b3 b6 ad ad a9 a7 a1 a3 a4 9b 93 99 97 9e 92 90 88 8a 88 86 8b 87 91 80 84 85 85 94 89 8c 8f 94 99 96 93 99 8b 8b 87 89 86 8c 80 8b 8d 90 8b 8f 88 8e 85 8b 8e 8a 81 83 87 8e 84 7f 7f 80 88 87 85 84 8d 83 87 76 74 70 6f 79 67 6e 6a 84 a2 af aa 97 7f 5f 50 30 20 17 09 05 07 05 06 06 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 05 05 07 0d 10 25 35 45 70 92 b9 cf c1 99 91 8b 8c 91 8f 88 91 91 90 95 9c 9b 92 9a 99 9a a0 a2 a4 98 98 a3 9f a5 a9 a8 a5 ad a8 ba ab b4 b4 bf bb b7 c0 b9 be c9 c6 c4 ca c4 c0 cd c5 cc c4 c9 c3 c7 cb d3 c8 d1 d2 d9 e6 e4 e8 e2 ee ef f0 f0 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f0 e9 f1 f3 ff ff ff ff fb fd f1 f0 e9 e2 da d1 ca c5 c7 bc b0 ad 97 be d9 f3 ff ff f9 f5 f0 e4 ed e8 db e3 d6 d4 d9 cd d6 ce c2 c4 c8 c3 c8 ba bf b5 b8 bd b6 b2 af aa b3 a8 af a6 a5 a2 9d 99 99 9a 92 8a 8a 91 86 89 88 80 82 88 7e 7e 7e 7f 86 7f 86 8f 8c 8b 8f 93 92 9b 95 8a 8b 85 88 85 84 86 82 88 7f 85 88 86 8f 87 85 81 87 7d 82 88 7e 7c 82 7e 80 7f 82 82 88 84 7c 7e 7c 75 6d 70 6e 6f 6c 70 7e 96 ab ad 94 85 67 50 3c 25 17 0b 07 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 18 1c 2a 31 4c 6e 95 b3 c4 bd 93 8f 8e 8e 95 99 8c 91 88 8f 92 94 97 98 95 95 97 96 9d 9a 9f a2 97 a3 a3 a5 a6 ab a7 ab b0 ab b4 bf b9 bc ba bf bc bc c7 c5 c6 c8 be ca c2 cb bd c6 c9 c8 d0 cd c3 cb ce d3 d3 d2 de e5 e2 e1 e3 e4 f1 ee fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 d6 c9 c3 c3 c5 c8 d2 d2 d3 d0 ce c9 c0 b2 ba af a7 a3 97 9d 94 8b 84 83 8a 90 a1 c0 e4 f5 f5 e8 e3 e2 da df d8 dc dd d1 ce c8 c9 c4 c2 be c0 bb ba c1 bf a8 b0 b4 ae ae a7 a7 a3 a8 9b 9e a2 9c 99 96 95 96 91 90 8b 89 90 86 84 7e 83 85 81 7e 7d 78 73 77 82 80 84 85 81 8d 95 94 96 90 8a 7e 7f 7a 84 7e 84 8a 87 81 7d 7e 88 88 8c 85 81 7e 82 80 7f 7d 75 7f 80 81 7b 84 84 7e 81 79 7b 6b 71 70 6d 6f 6d 77 76 92 a0 b0 a1 82 6f 4a 3a 25 1d 13 0d 03 04 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 02 06 05 03 09 15 23 31 3e 5e 7e 9b b1 cd b4 98 95 89 97 8e 92 92 91 98 96 95 93 96 9d 9b 9a 92 94 92 9c 9f a1 a2 a9 a8 a8 a6 a7
 af ae ab b5 a7 b0 b9 b4 b9 b5 ba bf be c3 c2 c5 cb c5 cd ce c7 c4 ca c4 c8 c1 c3 c5 d3 ce d2 d5 dc dc e1 e9 ed e2 e9 ea f8 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 d8 b8 ac 9c 8d 97 94 99 9e 9c a0 a1 98 98 94 91 8e 7c 73 79 74 73 77 68 69 65 63 68 78 a4 d8 e7 ed e8 e2 de d9 db d6 d0 d2 cc d2 c5 c6 c1 c6 c1 be be ad b1 b3 bb ab b4 aa af aa a1 a5 a6 a0 9c a4 98 9c 9b 94 8d 8c 8e 83 88 7e 82 7b 81 7f 7f 7c 78 7c 7f 7f 7d 75 7c 78 84 85 81 90 91 96 85 85 81 81 82 82 7c 86 83 7c 7f 84 87 8c 7f 84 84 80 8e 7d 85 7e 7c 82 82 7d 85 7f 7f 84 86 82 82 71 6e 75 77 6e 6e 6f 72 70 8b a1 ae aa 8f 7c 60 44 36 24 18 0e 07 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 0c 10 0f 2b 2b 44 60 78 9c be ce af 9c 8c 87 92 92 8f 90 95 8a 94 94 9a 98 9b 97 9c 98 9e 95 9b 97 92 a0 a1 a2 a4 a5 a9 ae ae b0 ad ab af b0 b8 b4 b8 bc b7 b5 c2 bc c3 cc ca d4 cc c9 bc c1 b9 c4 c4 c1 c8 c0 c9 cf d5 d8 d9 d6 d9 df db e7 ed f2 f6 f7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 ba a1 88 82 7a 6c 76 6f 7e 76 78 79 7d 7b 7c 7d 74 6d 69 66 64 64 5c 58 56 57 58 4a 56 66 9e ce e6 e5 d5 d5 d6 de cc d4 c8 cc c5 ce c3 c2 bf bd b6 b0 b4 b5 b2 b4 b0 ae ac a9 a7 9b a0 9f 99 9b 8d 9d 92 95 93 8a 92 91 89 8a 7f 84 82 7e 76 76 79 7b 79 72 78 78 78 72 77 75 71 7a 81 8c 85 8b 87 83 77 75 7b 7a 7a 7d 7b 7d 81 81 7c 7e 7f 77 81 7e 83 75 75 81 73 7a 80 7d 7c 7d 7c 7f 76 75 76 73 74 6d 74 6b 6c 71 6f 71 85 94 b1 a3 93 7c 5f 48 2e 28 14 11 06 0f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 11 18 1a 1f 2f 49 59 7c aa c1 ce af 8e 90 8a 90 95 90 98 89 92 97 95 98 97 99 97 95 90 96 94 99 98 9d a2 a2 9c a7 a6 aa ae a7 ad a9 a9 a9 a5 b4 b5 af a9 b6 b3 b5 bd c0 c6 c9 d0 d1 c5 c2 be c5 c5 c5 b9 c6 c5 c7 d2 d2 cd d3 d2 de dc df db e3 ef e8 f7 f8 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ba 8b 6b 68 5f 54 63 55 5d 64 6d 66 77 79 88 86 89 85 7b 67 62 54 52 51 43 48 50 48 49 46 57 92 c9 dd db d5 d5 d4 d2 d0 ce c7 cc c4 c6 b9 be b4 b9 ad ab ac b3 ae ae a6 aa ac a9 a9 9b 9b 9c 9d 99 94 94 90 89 8d 87 86 80 80 80 7f 7c 74 81 79 72 76 67 75 6f 72 6f 73 75 76 6c 69 81 7e 81 7d 86 89 84 7e 6e 7a 79 75 7a 77 7b 77 7b 7a 75 74 80 7a 78 7e 79 80 78 7c 7a 7e 76 81 79 7e 7b 72 76 6e 6b 6d 6b 6f 75 73 70 6d 71 79 90 a5 a5 96 81 67 52 44 32 1f 15 04 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0d 0b 12 24 2c 38 49 5e 80 a2 bb d5 b2 92 90 85 8e 8d 9a 97 95 94 90 8a 93 92 97 98 93 9e 97 94 93 9c 94 9b a2 9d a4 9f a9
 a8 a5 a6 ad ad af b3 ab aa b0 b1 b2 b4 b2 b9 c1 bf be ce ce bf c1 c6 b3 c1 bb c1 bf c4 c0 c5 cd cd d0 d4 d1 d2 d8 da e4 e7 e6 f2 f9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 a0 60 50 44 4c 55 4b 55 5e 5d 64 73 78 88 94 95 9a 8e 7f 6f 65 55 4c 46 47 46 49 3f 35 41 59 8c c1 d8 d5 cf cb cd c7 c3 c2 c3 c3 c9 c1 b7 bc b9 b1 b1 ab ab af a9 b0 a2 a6 a0 a5 a0 9c a0 8d 97 97 8d 92 8a 88 80 82 86 87 84 7d 77 78 7d 76 74 73 76 76 7b 68 75 78 6e 71 6d 75 73 78 7d 82 7a 82 83 80 7d 72 77 71 6e 74 7f 7d 76 78 71 7a 78 77 78 77 7c 75 76 81 79 75 77 75 7d 77 76 71 73 67 7a 71 74 70 77 6f 6e 74 75 6d 77 80 97 a9 9b 90 76 59 48 33 31 1a 16 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 08 0b 10 16 0f 22 36 31 4e 6a 87 a7 be c8 b4 93 8c 89 84 8b 8f 8d 8b 90 93 8e 97 8c 8d 96 91 8c 92 92 96 a0 9e a0 a1 a1 9f a1 ad ad b0 ae a5 ad b1 b2 a4 bc af a5 ac b3 af b7 c1 bc c9 cd c7 c1 bf c1 c0 c2 b9 b6 bd bd c3 c4 c5 ca ce c8 d2 d2 d7 d4 d7 e2 ee e9 f5 fa fe ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e1 9d 56 4a 47 42 41 4c 46 4b 58 5e 62 74 84 98 95 9d 87 83 6e 5a 51 48 41 36 34 38 3a 34 38 4b 87 b3 d1 d3 cc c0 ba c6 c0 c5 bc b6 b8 b6 b4 b8 a9 af aa b0 a9 b0 a7 a0 a1 a0 96 a0 99 9d 96 99 8d 89 94 8c 8f 8a 82 84 81 79 7b 70 74 6e 6d 75 70 76 75 6d 71 6a 74 6d 61 65 73 74 73 73 6e 7b 7f 74 7c 81 79 76 6f 71 70 76 75 79 7a 6e 79 76 74 78 7b 77 77 78 7d 77 79 7e 80 72 76 7d 73 7b 78 6f 7a 7a 71 72 6b 78 6e 72 73 71 78 7d 8e a2 98 90 78 60 4a 3e 2c 1f 18 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0b 0c 0c 21 29 32 48 52 6d 8d a5 be c3 b0 91 8f 81 8a 8c 82 91 92 91 92 87 96 8e 90 8c 95 95 8f 94 94 8f 98 99 9e 9c 9e a5 9e a6 aa a2 ad b2 a7 a7 a8 a9 ab a4 a7 a9 a8 ad b1 bb cf c1 c4 c0 be c2 c1 c5 b9 b6 b9 b7 bb c3 c3 c9 c7 ca d0 c5 d0 d4 d5 db dd de eb f1 fb fe ff ff ff ff ff ff ff ff ff ff fe f8 eb dd 9e 4d 37 39 3b 3b 3e 44 4f 55 51 5a 62 7b 89 90 8d 83 76 65 4f 44 43 3e 36 36 32 33 3b 2e 4b 75 aa ca c7 c8 c4 c0 bb bb bc b7 b9 b7 b4 b1 ad a9 ab ae a5 a5 ac a3 a5 a1 9d a4 99 90 94 95 92 8b 8e 8a 8a 88 8a 85 85 7d 7e 79 74 77 6f 6c 71 6e 6b 6c 6b 75 64 71 6e 65 65 6b 6d 6e 73 6f 72 76 78 7e 7f 6b 68 6e 73 72 6f 75 6f 6c 70 71 70 6a 71 71 70 77 67 73 7e 7a 75 74 72 7b 6f 78 7c 74 74 72 75 6b 76 70 6b 75 6d 70 69 6c 7c 82 a4 9e 96 7e 68 5d 3e 2e 22 12 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0b 07 0f 1b 19 24 31 40 59 74 8d ae cd cb af 8a 90 84 90 86 8b 91 86 90 8d 8c 8e 91 8f 8f 8f 8a 8c 95 8f 96 9c 9a 98 a3 9c a6 a3
 a4 a7 a3 a5 ad af a6 b0 a7 a1 a8 a8 a7 a6 a8 af b2 be c2 b3 bb c2 c2 bf bb ba b7 b9 bd c0 bf c3 c3 cd c8 c6 c6 cb c8 cc d1 d9 d8 e4 ef f0 f0 fd ff ff ff ff ff ff ff fe fb eb f1 e6 d5 9e 4c 36 36 30 36 4e 40 3f 50 4a 54 63 78 8e 8c 8e 7e 6a 5a 46 3f 3b 3c 35 31 2a 33 39 32 3e 65 ac c7 c2 bd b7 c3 be b7 b7 ab ad ae b0 ae aa aa ac ab aa a5 a6 97 9f 96 a0 98 98 95 91 8d 91 88 8a 85 86 87 89 84 80 7d 78 7f 72 78 70 68 6d 6c 6b 70 6a 72 66 65 73 6d 67 66 6a 71 6a 7c 79 6e 72 76 7f 6c 6f 71 68 6c 74 75 6c 71 75 75 6f 6d 6a 72 77 70 7e 75 7c 79 71 76 6f 7c 79 7b 74 72 72 7b 70 76 72 7a 74 6b 73 72 69 6e 71 79 96 a1 9c 8d 6c 53 46 33 22 13 17 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 0a 10 13 18 24 3a 4a 5b 71 93 a7 c2 d7 b4 95 86 7e 87 8c 89 8d 80 85 93 8a 8f 89 86 8f 8a 8c 91 89 8c 9b 90 9c 9b 95 9b a1 a2 a1 a9 a7 a7 ab a0 a1 a6 ad a7 a2 a6 a5 9f a3 a8 a8 b6 b1 be b9 b9 be b9 bf b4 ba b5 b0 be bc c1 c8 be c2 c7 c6 cd c9 cb d3 ce d0 e0 e0 ef f5 f3 f6 f8 fb ff fb fc fd f4 ee e9 e4 dd cb a0 46 3b 2c 2a 35 39 33 36 41 4e 58 5a 73 83 86 85 7c 68 4e 41 3d 3d 32 2f 25 2c 2f 32 33 2f 63 96 bd c1 bc c1 b5 b9 b3 b5 b6 af ab ac a7 a6 a5 ac a3 a5 a3 a8 9c a0 97 98 9e 94 94 8f 8b 90 83 8a 88 84 7b 82 7d 75 7d 76 79 71 6d 6e 70 70 71 6b 6f 66 6c 69 68 6b 62 66 6f 70 69 6e 71 71 75 76 78 75 6b 69 6f 71 6f 6c 65 70 6b 72 6b 71 6a 78 6d 76 73 70 76 79 76 72 75 73 76 77 6e 74 74 70 7a 6a 70 6f 6f 71 72 6d 71 71 6f 70 71 88 a2 a2 8a 80 69 53 3c 2d 1a 16 09 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0a 08 16 1f 35 3a 48 5e 77 95 b4 c6 cb b9 8e 88 85 7d 8f 8a 82 87 84 8f 8e 8d 8d 88 8e 88 85 85 90 9a 8b 97 95 9b 8f 98 a7 a4 a2 a6 a7 a3 a3 a3 a4 9a a7 a1 9e 9e 9f a0 a1 9e a3 a6 b1 b3 b7 bd b2 bc bc bb b5 b4 ab a9 b5 b9 be bf ba c5 bf be ca c6 c6 cb c9 cf df da ec f4 f8 f8 f7 f9 f4 f3 ef eb e1 e2 dd da cb 9f 45 27 26 28 2e 29 29 30 3a 40 48 52 5d 78 83 78 75 64 4f 3a 33 31 29 24 24 26 22 21 26 2d 5a 8f b2 b7 b7 b2 b0 b8 ae ac a3 a9 a9 a6 a7 a5 a0 9d a1 a6 a3 9e a1 9c 90 93 8d 8e 8e 86 88 86 84 86 7f 83 78 7a 75 75 71 78 6a 6b 6c 69 65 63 65 61 61 6d 5f 67 66 6c 62 67 6e 64 66 6b 65 71 6d 70 74 6f 6b 69 6e 64 64 6d 6a 6e 73 6b 6e 71 6d 72 6a 72 6f 78 75 75 6e 6f 72 73 74 78 76 6c 71 74 71 75 78 74 71 72 6d 70 74 70 6d 6b 75 7a 91 a0 90 7b 61 58 40 30 1f 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 0d 08 09 16 1a 29 39 4a 61 7b 9c b8 c4 d0 b6 87 82 7e 83 88 84 85 87 87 88 86 8b 8e 88 8e 84 84 89 8e 8f 8b 90 88 9a 9b 9d a9 9a
 9f a1 a0 9c aa 9d a7 a4 a4 af 97 9b a8 a1 a0 98 9d a5 a7 af b0 b1 ba b0 b7 b5 b6 ba b0 b8 b5 b0 bb b8 bb c1 bc be c2 bc cc c8 cd d3 db df e2 e5 ee f6 f4 f2 f0 e3 e0 e4 e0 d8 e1 cd c2 9c 45 2a 2e 27 26 23 35 2e 42 3f 4a 4b 5e 73 7e 7f 6a 58 44 32 37 34 2a 24 1f 24 2d 26 1f 36 4e 8d b2 bd be ac af ac ad a9 a5 a2 ac a0 a1 a2 9f a1 a9 98 a2 9f a0 95 95 8a 8a 91 8c 90 87 84 89 7b 78 7d 7a 70 78 73 6e 6c 6c 6f 72 6c 6a 65 69 65 60 68 61 62 6c 66 69 63 69 71 6b 66 69 6b 6d 71 76 68 71 66 63 66 61 69 67 6e 6b 6e 68 69 66 67 70 6c 73 6f 73 7f 73 73 72 68 76 70 76 73 73 78 74 77 72 6d 74 72 6e 6d 72 6f 6c 6a 6d 76 83 99 9a 81 70 5f 49 30 1e 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 02 0a 18 1a 1d 2e 3b 51 61 82 98 b5 c5 d0 b4 97 8a 7e 75 81 7d 89 8c 82 8a 87 86 8b 85 80 86 8c 85 93 91 96 90 92 97 95 95 9f 9e a1 a3 a1 a1 9d a3 9a 9f a2 9e a2 9d 9d 9c 9b 97 9d a2 ab a5 aa b2 ad b4 b2 b1 b3 b1 b2 ad ad b1 b6 b8 ba bc b9 bb c0 c1 c5 bf cf cd ce db e0 e2 ec df f1 e7 f3 e7 e2 dd df d6 d2 c9 bf a2 4d 2f 28 2c 27 27 27 2d 35 2e 39 4a 54 6e 78 70 64 53 45 34 2d 27 29 1c 29 1d 25 23 21 25 49 80 a9 ac ae ab aa a8 ab a5 a8 a5 a3 a6 a7 9e 98 a0 a3 9b 9b 9e 8f 9a 8c 8d 8e 84 8d 8e 82 84 7b 84 7a 7c 78 75 7a 75 6e 71 6e 6e 68 66 6d 64 6c 66 60 65 67 60 66 6a 5f 5e 6b 66 65 6b 66 6c 73 72 6d 77 6f 6a 6b 68 69 62 6c 6b 68 6f 6a 64 6e 78 6a 70 6e 76 6a 70 6d 73 76 6f 6f 70 7d 75 6f 70 74 72 77 72 73 66 6a 6f 6d 6e 6e 79 6b 77 83 95 9c 8a 77 5f 53 39 26 1e 0b 06 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 0a 19 29 31 40 5b 61 7a 90 b0 c6 c9 b0 99 82 7a 7c 7d 7d 7c 87 7f 78 85 84 84 8c 85 84 86 88 88 89 8e 90 95 99 9a 91 97 a1 9b 9b 9c a0 9a 9f 99 a0 99 9c 9e 9a 99 9a 9c 97 9d 96 97 a2 a5 b2 ae a8 b0 a9 a6 a9 a5 aa ac b2 b0 aa b2 b4 b8 b5 b5 b7 c1 b4 bf c6 c6 d5 d9 e1 ea e4 e3 e7 e0 dc de d5 d4 cf cf c4 b9 9b 48 24 1b 20 25 23 26 2d 31 33 3c 40 4e 60 70 60 60 4b 3d 26 20 21 24 1d 25 1e 18 1f 22 20 42 77 9e ab ae a2 a5 a6 a7 9b a6 97 a4 9a 96 95 91 9d 9a 99 9c 96 96 89 88 86 87 8c 83 7d 7d 78 7b 7d 78 79 72 6e 6e 70 6a 67 6a 6b 66 5d 67 68 62 63 68 5d 63 5f 5a 67 62 6a 6b 68 66 65 69 70 67 7a 6b 67 69 61 68 63 5c 65 63 6c 64 67 6a 70 6a 6f 68 69 6d 6e 71 6d 6d 70 6b 67 67 6c 6f 74 6c 6f 6e 74 73 76 70 66 68 6a 6b 69 69 70 68 6f 77 88 a2 92 7f 68 56 41 25 16 10 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 10 13 1d 2d 43 58 61 76 96 b4 c1 d7 bd 96 84 71 73 84 7a 7e 7e 7d 7a 83 7e 8f 89 84 85 87 8b 87 90 8a 8e 8a 93 92 9e 9e 97
 9b 9f 9e 9b a2 94 9e 92 95 9e 93 95 9b 93 8f 99 95 92 9c 98 ab aa ad ad ae ad a6 ab a3 ab b0 b1 ae ae ae b5 b9 b4 b7 ba ba ba b9 c0 ca cb d1 d4 de e8 e2 dd d7 dc ce cf cb c9 cf c1 b1 9d 45 1a 12 1b 1a 18 32 20 35 31 2f 37 4a 67 66 61 5f 4d 39 2a 1d 1c 16 1a 16 21 1f 23 22 27 39 74 a0 a9 a6 ab a4 a3 9f 9f 9b 9f 99 90 8f 9a 92 a0 96 97 96 91 90 92 86 7d 83 7b 82 84 7d 7f 7c 76 70 75 76 6c 74 71 66 6d 6d 5f 68 66 69 5d 63 5d 61 5b 61 5f 61 66 65 60 63 64 63 66 61 6f 73 71 68 6c 65 6e 65 60 60 65 62 5c 64 68 64 66 62 6e 6a 6c 6c 6c 6a 6e 6b 6c 69 6b 6c 65 72 6e 70 6f 70 6e 76 6e 6d 67 68 6c 69 6d 6d 6a 6c 6e 74 84 97 99 7f 6a 54 3a 28 1a 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 07 1c 19 24 36 4b 51 6d 7b 9b b8 cb cc b9 8e 7c 70 75 7e 79 7f 84 84 7a 7a 84 84 82 81 84 82 86 96 8d 8a 98 94 9c 98 9b 9e 9f 98 98 9b 96 9d 9b 93 95 92 95 99 92 98 90 94 94 98 90 93 95 94 a6 ab ac ac a9 a3 a6 a5 9e a2 a9 a7 a1 af b5 b3 b0 b6 b6 ba bb b6 c1 c5 d1 cc d3 db dc e2 d8 d6 d5 cb cd d3 c1 c7 bf b2 8b 40 1f 23 1b 13 1e 20 1f 24 33 2a 3b 48 57 67 60 55 48 2b 1f 17 1e 21 19 1b 16 21 24 22 2e 33 5f 95 9a 9b a9 9c a5 9e 9b 96 94 9d 99 94 8e 91 97 95 92 96 99 95 94 89 7e 81 87 7d 7e 78 75 76 78 7c 70 71 71 6d 71 5f 6b 66 66 68 64 68 64 5f 5e 5f 63 62 5f 66 6a 62 67 67 6b 61 63 73 6a 6f 67 6a 64 69 6b 66 65 66 66 6d 64 61 67 6b 64 66 68 66 6b 6f 6b 6b 6d 6d 6f 6b 6b 70 6e 72 75 6e 70 6f 6a 6e 6d 6d 71 63 69 6e 66 68 66 64 64 75 7f 8d 9a 89 65 54 3e 29 1f 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 04 00 11 08 17 29 31 47 5f 6f 87 9a b7 ca c6 be 91 87 73 78 7e 7e 80 84 7f 79 82 80 81 87 86 80 81 86 8a 91 8e 93 95 98 90 97 9b 96 92 a1 96 91 97 9c 8f 97 9a 98 8c 8a 90 91 8d 8f 94 8a 86 94 96 9f a7 b2 ab a2 a2 a5 a6 a8 a7 a4 a7 ad ab b3 b5 b0 b2 b3 b1 ae ab b9 c4 c1 d2 d0 da d6 d3 c4 ca cf c4 c5 c8 be bf b7 a0 84 46 29 10 14 1a 14 2b 1e 23 2a 2d 38 3d 48 61 58 51 3c 25 21 16 1c 1d 14 23 1c 1e 1f 1e 22 2d 62 87 9e a1 a3 9c a5 99 93 95 96 92 94 92 97 94 99 95 92 94 93 8b 89 84 88 84 82 89 82 75 76 6f 72 76 70 72 72 6d 67 6e 69 69 65 61 67 5d 62 5f 5b 63 5c 5c 55 5e 6a 65 66 66 57 5d 65 68 71 61 62 63 64 5c 6d 5c 63 5a 5e 67 64 61 60 67 66 63 65 5d 68 65 6e 69 6a 6d 6b 6f 6c 6a 64 6a 6e 6a 6d 67 6c 6b 6d 6b 6f 61 62 69 66 6a 62 6b 65 6b 79 8b a4 8c 7a 5b 41 2c 1e 0d 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 12 24 2b 37 4b 52 69 84 a2 b2 c4 cf bc 99 80 73 76 7a 7b 7b 77 7e 85 85 83 83 80 82 83 8b 89 8c 8e 90 91 95 93 95 96 90 98
 95 90 96 93 8f 91 8e 92 93 91 90 86 8d 92 8d 91 90 83 86 94 90 a2 a6 9d ae 9d a9 9e a5 a5 a1 a1 ad ab aa b1 a6 ab b6 aa a9 b6 b2 c2 bd c6 c8 c1 d2 cc cd cc cb ca c3 bc b9 ba b7 b5 af 88 50 26 19 17 18 18 21 1e 28 27 29 2f 35 45 56 56 4f 41 32 16 19 10 11 20 1c 0f 15 19 11 1a 24 59 87 99 a0 92 96 93 93 92 94 8f 99 90 89 8f 92 97 8c 8b 8b 8b 90 89 87 7c 85 84 7b 73 78 80 73 74 67 72 6a 6f 6b 67 72 60 63 62 65 66 63 67 5f 5f 5a 65 5d 61 63 63 63 5a 5f 60 65 6f 64 6f 67 6a 65 6a 64 5d 64 62 5e 62 65 61 65 60 5e 63 5f 6a 67 68 6a 69 6f 64 6f 5c 62 6f 66 5f 6c 64 5b 68 6f 62 67 6b 6b 69 61 6e 6c 68 65 66 61 65 6e 76 87 9a 91 7e 60 4a 32 24 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0c 24 24 42 50 5c 68 80 9f ae c7 c1 b7 98 7b 78 74 72 79 7b 80 78 7e 85 7d 80 83 83 85 85 8c 8d 8c 8e 8f 94 91 8f 95 96 92 93 95 93 8d 96 95 9b 8f 91 8e 90 8e 8c 8e 84 86 88 92 8e 8d 8d 96 9c ac a2 a7 a9 9f 9d a1 9e a5 a3 aa b1 b0 b0 b2 ae a9 ad ab b8 b9 c1 c6 be c3 ca c2 c2 bf bf c0 b5 b7 b9 bc b7 b2 a8 95 54 22 12 10 13 11 18 18 26 24 2b 2e 31 43 4d 58 4a 3a 25 1b 0c 14 1a 14 1c 15 16 18 1a 1e 21 4a 7f 8b 95 91 91 93 93 96 87 89 8e 8e 8b 8b 8d 95 90 90 8d 88 87 8d 7b 7e 7d 7b 7c 75 73 72 6f 6f 6c 77 6e 6b 6e 64 69 6b 69 60 5f 60 5a 61 5e 62 60 64 65 61 67 60 5e 61 64 5c 6a 63 76 6b 66 6a 62 63 5d 62 67 66 64 5e 66 63 66 6b 66 66 59 67 64 67 61 66 64 66 63 63 65 6a 67 68 65 68 6a 6f 72 67 6c 66 6f 6a 65 64 5e 67 6f 67 6f 6d 65 73 80 98 93 7a 61 48 38 2c 0e 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 15 21 2b 39 4c 5b 74 85 9e a8 c4 c4 bf 8e 7f 70 71 78 7c 7c 7a 79 7b 82 82 84 7f 84 88 89 85 8c 8a 8e 96 8d 93 92 8b 8e 8d 8c 8a 90 8a 8a 93 87 8c 90 94 8d 88 88 89 8b 87 88 83 88 88 88 94 9e a5 9e 96 9c 95 92 8c 97 9e a6 aa a5 af ac b4 a0 ac ab a6 ac b3 b8 bd c2 c4 c6 c1 c2 b4 b2 af ae b1 b1 ad b4 aa a2 a0 5c 1c 12 13 16 11 15 1b 1a 21 20 30 37 33 4a 48 41 35 20 19 0e 0d 11 16 10 14 0f 21 10 19 21 42 74 8d 8d 94 92 87 81 83 8d 8a 8a 84 8a 8b 89 8a 8b 8d 8a 8a 89 83 7f 77 79 7b 77 73 74 77 75 74 68 75 67 73 70 5e 69 63 67 66 67 60 5c 62 5f 5f 60 54 65 61 68 60 5f 5f 5f 64 6e 69 69 5c 5f 64 61 61 5d 60 62 5e 5a 5b 5d 64 5e 5c 61 5d 61 5d 6a 64 67 64 65 6d 61 69 6a 64 64 63 66 64 68 65 69 64 66 65 66 6a 69 64 65 68 68 66 6a 60 67 6d 7d 92 8d 7c 69 4a 37 22 10 06 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 06 14 13 1f 2f 3c 4a 57 71 7f 98 af ba c7 b4 98 83 67 6b 72 72 73 7d 80 7e 75 7f 7a 76 8b 81 87 82 87 8d 8e 93 8e 92 95 8f 89 8d
 89 94 8f 8e 84 8c 87 83 8b 85 85 8d 8b 7b 8b 88 81 89 86 8f 8a 91 9c 9b a0 a3 8f 89 90 90 91 96 9f 9f a9 ad a8 ac a6 a1 a7 a4 ac b5 ad bb ba bf b8 b1 b8 b6 a9 af b1 a7 af af b1 ad a0 99 5f 20 13 0e 0d 13 0f 19 1e 23 20 26 2a 33 3f 3e 3e 32 1d 13 12 0a 0a 0d 0e 14 11 10 0e 16 1f 37 7d 8c 91 8d 8c 8f 87 88 89 88 8d 8b 8c 8a 8e 83 86 8d 88 8c 86 80 7e 86 7a 7b 72 79 6c 75 67 76 6b 71 66 6f 70 67 70 68 65 6b 5a 64 65 5f 65 59 65 63 61 62 6a 5f 60 5f 63 68 6d 6f 63 64 5f 61 60 6a 5d 55 59 5b 5c 60 5a 59 61 5f 62 5e 5c 61 62 62 6a 6b 62 62 5e 61 64 65 62 68 60 5f 64 63 63 66 63 64 5a 66 5f 68 60 64 66 62 62 63 63 70 72 8f 92 7f 69 4f 39 2b 10 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 10 15 24 2b 3f 55 5d 75 83 99 af c2 ba b4 97 79 6e 72 71 71 7c 73 81 77 75 74 79 82 85 83 89 88 7f 91 8a 86 92 8e 8b 8b 8d 93 89 93 89 86 8c 8d 8f 8a 85 84 85 84 83 8e 84 85 7d 83 85 84 87 8c 94 96 a4 99 87 8f 8a 8b 91 9a 9d a8 9f a2 a0 a3 a1 a5 aa a3 ab b5 a6 b0 b3 aa b5 b1 b2 a9 a7 a1 a4 aa b1 a5 ad 9e a8 94 67 24 14 15 12 18 19 18 17 1a 17 1f 26 38 3a 44 3a 2e 16 0f 17 0e 13 11 11 10 10 17 15 19 1f 33 6d 88 8a 84 87 84 86 85 7f 8c 89 89 86 8a 8f 8d 8c 84 89 82 81 82 79 76 71 75 75 73 71 7a 6e 78 71 6f 71 6e 6c 6d 64 69 65 65 5b 60 64 62 5f 66 5c 69 6e 62 62 64 62 66 6c 69 6b 70 68 66 67 63 5b 5a 5e 63 5c 63 58 5a 5d 62 64 60 65 5e 5d 60 66 64 65 6e 5d 6c 63 62 6a 61 67 64 5d 67 64 6a 65 6c 6d 64 65 64 65 62 62 67 66 65 67 6a 62 69 7c 84 8e 83 6c 4a 32 2d 11 0d 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 12 2d 32 46 55 5c 71 7f 9d af bc bd bb 9c 81 76 71 73 7d 7d 74 77 76 72 80 7f 7d 80 7d 83 86 84 8a 8c 82 86 85 8f 8b 8e 88 89 89 8a 8b 86 83 86 8c 86 8a 82 7f 85 81 83 82 7e 85 81 83 84 87 98 90 9c 91 85 89 86 83 90 96 98 a0 a3 a2 99 9f 9f 9e 9e 9c a6 ab b4 b0 b2 b3 ab a7 a7 b0 a7 a9 a7 ae a9 a0 ad 9e 98 98 73 2d 14 0c 0e 0a 11 16 18 19 18 21 26 2c 37 3c 3e 33 19 13 06 0d 08 0c 15 0c 12 0c 11 17 14 3a 65 80 8c 82 82 81 7f 85 87 86 84 8c 85 87 84 8a 90 88 87 7c 81 78 7e 7d 7b 7b 6c 6f 6f 6f 71 69 6b 6f 6f 6f 6b 64 68 60 60 60 6c 63 66 64 63 5e 60 58 64 60 5e 6b 56 66 67 6c 70 69 65 62 5d 59 5f 5f 5e 60 64 5d 59 5d 65 60 5b 5f 62 5a 5a 67 61 5d 61 69 63 5f 5e 62 68 5b 62 62 5f 64 60 64 64 64 69 5f 66 62 5a 66 63 6f 62 63 62 69 62 67 75 84 90 80 6b 4f 33 26 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 06 06 1a 1c 29 40 50 58 6c 83 99 a5 b0 be ae 91 83 6f 6c 67 75 74 70 79 73 76 79 74 7d 76 7b 80 7a 84 83 88 8a 86 87 8e 8a 88 84
 8d 86 84 83 80 83 84 86 7f 84 7c 87 7e 7c 7c 81 78 7a 7e 7f 80 84 92 9c 9f 91 80 83 84 88 8a 90 92 90 8e a1 9e 95 94 96 a4 8f a8 a0 9e a9 a5 ae a4 a0 a5 a1 9b a1 a0 a2 a8 9f a0 9a 96 91 61 26 13 10 06 0c 0a 10 0d 18 1a 19 1a 24 2a 31 36 2b 1c 0e 06 05 0a 0a 08 07 05 10 0c 0f 14 2c 5d 7d 83 7b 80 80 7f 80 81 83 83 7e 7c 81 81 8d 89 8b 85 81 7c 78 72 7b 74 75 74 78 6a 71 6f 6f 64 64 6b 6c 67 65 64 6b 6c 67 60 5d 61 61 5c 61 5e 62 5d 58 5f 63 62 68 71 6f 64 65 65 5f 57 5e 5e 59 5f 58 59 64 53 52 5d 5e 62 59 52 5c 57 61 5b 62 5d 64 5a 68 54 60 5d 5c 5f 65 5c 63 5c 61 65 63 5e 5a 62 67 58 5d 5d 64 64 65 60 64 64 69 6c 7c 8e 7f 6b 51 38 29 09 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0e 1a 1e 2f 40 51 5e 74 7e 94 a8 b5 b2 b4 92 85 6d 71 6a 6f 76 76 6e 76 77 7a 79 74 73 73 7a 7c 80 87 84 85 83 86 88 8a 89 8a 84 8a 79 86 88 7d 88 84 87 7f 7d 82 7d 7c 83 7d 73 7b 7a 79 7a 81 89 95 94 8a 8b 81 83 80 7c 87 8f 93 99 98 94 93 92 90 9a 9d 9a a0 9d a9 ac a8 a7 a3 9a a5 a2 95 a0 a2 9b 99 99 98 8d 92 6d 30 0e 07 0a 0d 10 14 15 19 11 1e 17 26 31 2e 2f 2a 19 08 0a 05 04 06 0d 05 08 11 08 0f 19 21 5e 7e 7b 7d 79 7f 7b 7f 85 81 88 84 84 84 88 8c 8a 7f 78 7b 77 79 77 70 73 71 70 6a 69 6c 6e 71 6a 71 63 6b 63 6e 65 63 60 65 66 62 62 56 5c 67 61 5f 64 60 64 64 5d 67 6c 6c 69 65 5c 5f 60 5f 5c 60 5d 5b 5a 5a 62 5a 64 5d 5e 5d 62 65 60 5c 62 61 5c 5b 69 62 57 5c 5e 62 63 5e 61 61 59 5c 60 5a 5a 5b 62 60 65 63 64 60 65 61 69 67 5f 60 66 75 8c 7e 68 52 37 2a 13 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0d 1c 16 2c 40 4d 5a 70 7a 93 9f af b7 af 99 81 72 69 6f 66 6e 70 6d 73 72 72 75 75 77 77 73 7d 80 83 89 87 84 83 85 80 84 83 85 87 87 7e 7c 80 81 7a 7a 82 7c 7e 7e 82 7a 75 7a 7a 7b 7a 7c 81 8e 92 8c 88 83 7a 75 7b 86 85 90 8a 92 8e 92 91 95 94 96 95 9a 9c 9c a1 9c 9d a3 9d 9c 98 97 9a 9e 9f 99 98 98 92 8b 93 71 2a 0c 0b 08 05 0a 0e 0e 10 0b 15 13 1f 24 35 31 25 0d 0d 06 05 03 04 06 10 05 0f 16 09 11 27 4c 7a 7a 82 76 82 7b 7a 86 7e 7e 8a 7c 80 7e 82 85 8c 81 7f 76 76 6a 6b 74 75 6a 70 6d 71 6b 6c 6c 6c 63 6a 63 69 6b 65 5f 66 6a 63 64 61 5c 5b 61 5f 62 5f 66 61 71 6f 68 69 63 60 61 57 60 60 60 5d 5c 5a 5b 5a 5a 62 64 56 55 5e 60 6e 5d 63 5c 5d 58 64 65 69 63 58 5b 55 5d 5e 5a 64 5f 62 61 5f 65 5a 5f 65 62 5f 60 63 62 5e 62 64 62 60 65 71 80 76 6c 53 3d 2d 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 02 06 1a 19 2f 45 4b 60 6b 85 88 a3 af a9 a2 88 7b 74 6e 70 6b 74 68 71 67 71 6c 6e 79 73 77 75 78 82 82 7e 82 8b 8c 88 83 8a 84
 81 7d 7d 7a 7d 76 7d 80 7d 7c 7b 78 74 7b 74 7b 7e 76 70 79 74 7b 89 90 91 86 7e 72 75 7b 7d 7b 81 82 83 8c 8a 90 84 8b 8d 8b 8c 97 94 99 94 9b 9e 99 97 96 8e 9a 94 98 92 8e 96 91 96 87 72 31 0a 06 10 0a 06 0f 13 1a 0a 0d 0d 17 2b 30 25 23 0a 00 06 05 03 06 0b 05 0b 06 0b 0d 0d 21 50 6b 7a 76 75 78 6f 7b 80 84 81 7e 83 83 81 85 89 83 7f 7c 78 74 73 67 6d 6b 71 75 73 70 73 65 6c 6d 60 6e 66 6b 69 65 68 6b 63 61 64 64 59 5d 59 5c 61 5d 67 66 6e 6a 66 65 61 60 5c 5d 61 5d 56 61 60 5c 65 5c 5c 5d 58 56 5c 5f 58 5b 5a 5b 52 5c 61 5b 5b 59 57 5a 62 52 59 5b 61 51 64 64 5b 60 5c 5b 64 5e 5a 57 61 64 63 5d 54 61 5a 62 60 6f 7e 79 70 4e 3b 2f 17 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 06 0b 16 21 2d 40 4b 5e 6e 82 97 a1 a6 a8 99 8a 77 70 6e 6a 73 6b 6d 6e 72 7b 6e 73 73 70 78 74 75 81 7e 80 81 82 84 89 86 81 83 83 82 84 7d 83 7b 7f 84 77 80 79 79 7c 7d 6d 76 7a 71 80 77 6f 75 80 84 8a 90 7b 81 77 77 7d 7d 85 8d 89 89 7e 82 85 85 86 8a 8b 91 8e 90 95 98 9c 97 96 95 92 91 8f 8b 95 90 85 90 8a 85 6f 2c 0d 02 0b 14 0e 09 14 0a 0b 09 16 16 1c 23 2b 20 0c 09 07 05 03 03 0c 09 08 0f 07 13 0d 19 47 6c 7b 71 7a 75 74 7a 7b 7b 7f 7b 7c 7d 79 86 86 82 82 81 79 7c 6c 70 74 6c 73 66 6b 68 6b 6f 6a 6d 67 67 65 66 63 62 5c 5f 5c 5c 68 65 64 66 60 67 62 68 71 67 6b 66 61 5b 64 5e 5f 5e 60 5f 5c 5c 5e 5a 61 56 55 5a 5b 58 60 5e 5c 5f 56 5c 5c 5d 65 5e 59 5a 5b 54 5e 57 5e 5f 5d 56 5a 5a 5f 66 5d 60 63 64 5c 5f 5f 5f 60 5f 5d 60 56 60 62 64 7f 86 71 59 42 2f 15 10 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 06 01 0e 0d 22 29 43 4f 62 71 78 87 a2 a2 9e 92 80 78 76 72 75 72 71 67 77 6b 77 69 6f 74 78 6d 71 77 75 7d 80 7f 80 7e 7c 7f 7a 82 7b 81 81 7b 7c 77 7c 75 81 7a 6f 77 76 77 70 79 77 78 73 7a 74 7d 7e 83 7c 83 84 7c 7b 74 78 7f 78 7b 86 81 85 8c 81 84 8d 84 8d 8a 8f 8f 93 98 91 91 8a 90 96 98 94 92 99 96 9e 8e 88 89 70 30 0f 04 06 08 07 00 0b 0a 06 0b 11 1e 1e 24 25 1d 09 0d 06 09 03 05 06 0a 07 09 0f 09 10 10 3e 6f 78 79 79 76 76 6c 7a 7d 7b 81 79 83 7b 86 89 86 79 7d 7a 70 6c 6c 72 71 65 6d 6f 6f 67 72 6a 6c 66 68 66 68 61 63 6b 62 61 64 62 59 62 60 63 64 67 69 68 7c 74 65 66 65 5e 61 67 56 5d 61 61 64 62 64 5d 55 54 5b 5f 58 5b 5e 5c 53 57 59 5d 56 56 61 5e 64 5c 60 5d 5c 5f 5e 58 5c 59 5c 61 63 5f 5e 59 64 66 60 64 5f 63 5a 66 5c 60 58 5c 67 6e 7a 68 55 44 2e 1d 0c 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 14 1e 30 38 56 5c 67 80 8d 9c a2 a0 85 73 6f 6e 70 6f 69 72 64 61 69 6b 6e 71 65 70 6f 6f 70 73 79 7d 7c 80 87 73 73 77 7b
 75 7e 75 78 7a 7d 78 7d 7b 79 6d 7b 73 67 76 74 73 74 71 73 76 6d 7c 7d 86 7d 7b 75 71 74 7d 78 78 7a 7a 84 7b 80 7e 7c 8b 78 81 84 8d 90 8d 92 92 89 8d 8c 8e 95 94 93 96 89 8c 8a 82 82 75 33 0d 05 08 07 09 01 0c 08 07 0b 06 0f 21 1a 17 16 09 00 06 05 03 00 07 05 0c 0f 06 05 0b 12 3b 67 73 79 6e 71 6a 78 73 77 7b 76 7e 7c 73 7c 81 7e 81 7d 6d 76 72 6a 6a 64 6f 6c 6a 70 70 66 67 68 5e 6b 64 67 65 62 65 64 61 68 5c 5e 5f 62 5d 64 61 6e 75 72 6b 64 69 6a 60 61 5c 5e 4f 5f 5d 5a 5a 56 57 64 55 58 62 55 5d 5b 5c 58 5f 58 64 59 59 61 5d 58 5c 56 55 59 5f 59 5c 55 5b 5d 5c 63 5d 56 64 5b 64 5e 5d 5a 5b 5c 60 5a 58 5a 5a 61 79 71 78 56 3f 30 18 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 15 1b 2e 3d 49 65 66 7e 8d 9a 9c 91 7f 74 62 6e 68 6c 65 6b 6e 6e 6f 6b 72 75 6f 69 6e 7c 73 75 7b 73 7e 7d 81 7e 7d 80 7c 7b 73 76 76 6c 73 71 75 79 76 75 75 72 76 67 73 74 66 71 6e 6d 78 70 7e 7d 88 7d 7a 71 74 76 75 71 77 75 7f 77 76 7e 80 7a 82 8a 82 80 85 83 88 8e 87 8c 8b 8d 8a 8d 8e 95 95 94 8a 82 83 6d 3f 12 0e 07 05 06 06 06 0c 03 09 0d 0d 15 12 16 14 05 07 06 05 03 00 08 09 05 09 09 0f 05 11 3a 67 71 6e 6d 6e 73 6d 77 78 7c 77 72 81 78 84 83 7c 80 7c 79 76 6c 6b 6d 6b 6f 6a 63 68 63 6d 5f 65 69 6b 62 6d 5f 65 63 60 58 63 5e 64 65 68 66 6c 6c 66 72 72 62 5d 5f 5a 61 61 5e 58 5e 60 5c 61 58 54 5e 57 57 5c 5d 5a 61 5e 59 53 5b 54 56 62 57 5c 5c 57 61 59 54 53 55 59 55 55 52 56 60 5e 62 54 5c 61 5e 5e 5e 5d 58 55 56 57 63 5a 5f 65 6a 78 6b 58 3f 2d 1b 0e 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 12 1e 2a 3e 53 62 6b 7f 8c 93 a4 93 7e 6e 6c 64 6d 6a 6f 6b 71 72 73 72 6c 6a 75 75 6c 73 68 70 77 7a 7b 7f 82 77 78 77 79 79 7e 7b 75 74 6f 7b 78 72 7e 7a 74 6f 70 6c 69 6c 73 6d 74 6d 72 7b 7c 8a 7c 79 78 7c 70 76 76 6f 79 72 7f 7c 7c 76 80 7a 83 7e 85 85 80 88 8a 80 8f 8c 84 86 89 8e 93 8e 8e 93 92 84 86 76 3e 10 07 06 05 07 0a 09 07 07 08 0d 0c 12 14 19 1c 0c 0b 06 0a 03 00 0b 0a 03 05 06 09 0c 0d 2d 59 76 6f 75 78 77 7a 6a 75 7f 74 72 79 73 7e 83 87 77 80 80 7a 72 71 78 6f 6d 72 6a 69 6c 68 66 6b 67 5e 70 6b 63 67 68 68 5f 62 65 64 65 66 66 69 6a 6e 72 7b 69 5e 67 5f 65 61 5d 56 53 5e 5c 5b 5e 59 57 5d 54 5b 5f 5f 61 5f 60 5e 60 5f 69 67 5a 5e 51 61 5e 5b 5b 5f 4f 5a 5b 5a 61 54 5f 5b 56 59 57 5d 5e 58 65 5c 5e 65 5b 5e 5e 5f 5b 67 68 70 65 54 43 2b 19 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 16 1a 28 42 4b 5b 72 7e 84 91 95 94 7a 69 6b 61 63 6c 6a 63 72 6e 71 6f 71 72 6f 6e 6f 6e 6e 70 6b 70 72 77 82 73 71 6e 75
 7c 7f 75 73 77 6d 74 74 72 72 69 75 75 6b 70 70 66 70 69 71 67 70 71 74 7b 78 7c 7d 6c 6d 70 74 6c 6f 6b 6d 77 7a 6b 7d 76 7e 81 7f 82 81 7f 75 8a 80 85 8b 86 87 8c 92 93 91 82 82 80 7d 75 44 16 04 06 05 03 08 06 09 08 03 06 05 15 0a 0e 0e 03 04 06 05 03 04 06 09 04 0e 08 08 08 13 2c 5f 6c 72 73 6e 69 78 6c 7b 73 80 7a 79 7a 80 7e 76 80 7a 7c 7c 74 6b 6e 61 6a 6b 6c 6c 6a 65 61 6a 60 69 65 67 6a 66 65 64 63 5d 65 64 6f 6e 68 66 69 62 71 70 62 5f 61 62 5e 5c 58 56 5a 53 5d 5b 5c 58 59 5c 5b 53 53 59 64 61 65 5a 5c 57 5b 62 60 5e 5e 5c 54 55 5c 4c 53 55 5a 5a 5d 55 5b 5c 62 56 5b 59 5b 58 5b 5b 5d 57 61 57 5c 5c 4f 65 64 71 6c 55 42 2f 13 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0d 25 36 4a 5d 69 7a 86 96 97 8d 7b 65 6a 66 65 65 5f 6b 66 6c 72 6e 76 73 70 6f 7a 6e 71 72 71 6a 75 6e 76 76 79 7e 75 71 76 6b 74 73 73 71 73 75 77 6f 6c 6b 6b 6e 6e 6f 68 6f 6b 6c 63 69 6a 78 75 7a 77 72 6e 6d 69 70 74 72 7d 78 71 70 7c 78 7d 7f 71 79 7d 79 83 7f 78 7c 85 84 89 86 8e 8a 95 92 88 83 82 7d 41 0e 05 08 05 03 00 07 05 03 03 06 05 07 10 12 08 05 07 06 05 03 00 06 05 07 03 08 0b 04 0a 2a 54 73 70 79 78 70 6e 76 72 7e 7c 71 75 72 70 78 7e 7a 79 7a 77 7b 70 6d 6c 69 6a 6d 68 6e 65 66 65 5f 62 70 66 65 69 66 68 64 64 72 6b 69 69 6c 68 65 65 79 69 61 60 64 5f 60 5a 5c 62 5d 5f 5c 59 58 56 5e 54 55 5b 63 54 57 59 60 59 59 62 5c 5c 61 5c 5c 60 58 5c 54 53 59 4c 55 53 57 59 59 5b 53 5e 53 56 51 56 5a 5f 5b 5b 60 56 52 5d 5e 5b 5f 6e 66 5a 42 30 16 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0f 20 39 51 62 70 81 84 91 93 82 76 64 65 5d 6a 62 6d 62 69 67 69 73 6c 6e 74 70 6c 6c 70 74 75 7e 77 72 75 6c 77 7c 70 75 78 76 71 6c 69 67 6e 67 76 6b 6e 75 6b 73 66 69 6f 73 6f 6a 6a 67 70 73 78 81 78 79 74 65 6f 72 6b 73 77 6e 75 78 74 78 70 73 76 7b 75 7c 80 80 81 7f 76 80 8a 91 8a 96 97 92 94 8f 86 78 4e 08 07 06 05 03 0a 06 05 05 00 06 05 10 0b 09 05 0b 00 0a 05 03 00 06 05 04 07 06 05 07 0e 28 51 64 73 72 74 72 70 79 7c 7f 75 7a 71 6c 75 78 7c 7e 83 77 77 79 7c 76 71 72 6f 69 6f 65 66 62 6d 6a 67 60 69 64 62 6f 64 63 67 66 66 6a 6e 6c 5f 61 64 75 69 62 67 5d 69 63 63 5d 5a 54 5a 5b 5e 64 57 57 57 54 58 5e 5a 5c 66 65 65 59 5f 5e 5c 64 6d 62 64 55 59 50 58 54 58 56 54 55 51 5f 5c 59 50 5f 5c 4c 58 5a 59 64 5d 5c 5b 5c 61 60 5b 68 66 67 59 3d 2b 18 06 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 24 2f 47 5b 69 81 84 8f 94 84 70 64 66 5b 66 62 69 68 61 64 6e 69 73 72 74 77 70 70 71 75 75 77 6f 6e 6c 6e 71 71 73
 6f 76 71 6c 73 70 6e 6e 73 65 6e 67 6f 72 68 67 72 69 69 67 6c 6b 67 70 74 74 71 6f 75 6d 6a 73 75 74 6c 72 63 70 75 70 79 6e 75 74 7d 71 73 78 7d 80 78 83 7b 80 8a 85 97 94 8f 8c 87 8d 78 4b 15 0e 06 05 03 00 06 05 03 03 06 08 05 09 08 07 03 00 06 05 03 00 06 05 07 00 0b 0b 03 07 25 47 62 70 73 72 77 75 76 7d 75 7c 79 76 6b 7c 7e 6c 83 7b 87 7f 7b 79 6e 6e 67 60 66 60 63 61 63 65 5d 67 62 6d 69 67 64 5e 63 6a 69 6f 6c 6a 65 63 64 67 6c 68 60 5d 62 64 5e 60 5a 5a 60 5d 61 5b 5c 58 55 60 57 5f 5f 64 5d 61 60 55 55 59 5d 58 5e 65 5d 5c 54 58 52 53 53 53 50 51 4e 5d 56 59 53 57 58 5a 4e 52 60 5d 5c 59 5f 50 56 60 57 5e 63 63 65 51 39 26 11 0a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1a 2b 47 54 66 79 84 87 90 7e 70 5b 5b 62 65 65 6d 6a 66 6b 6d 6d 6e 6d 71 72 74 6f 78 74 6d 75 6a 71 71 73 75 72 65 6a 6f 6a 63 6b 6a 69 64 68 69 6f 61 66 66 63 6c 6a 69 66 64 69 65 72 62 6e 6f 75 72 72 6f 6d 76 72 6f 75 68 73 70 73 6f 74 6e 77 76 6b 70 75 79 77 7a 72 6d 7a 7a 86 8f 90 96 93 94 7e 83 7c 56 15 02 06 05 03 00 06 05 03 00 06 05 03 08 06 0d 03 04 06 05 03 00 06 05 03 00 06 05 03 09 19 4d 6f 74 76 76 79 6e 77 7a 7a 75 74 72 72 7b 73 77 73 7d 76 7b 79 7c 77 6e 70 73 6a 70 69 6f 65 67 62 60 66 66 5f 64 6c 6b 69 6e 6c 6a 63 6d 62 67 5f 60 70 6e 64 5f 63 63 5e 56 56 58 5c 5f 5a 5e 59 5a 54 59 58 60 57 55 5d 5c 59 5e 58 5f 65 64 67 5f 61 59 5a 5a 5c 54 54 54 50 55 56 52 5a 51 50 4d 54 55 57 53 5e 50 53 55 58 60 5b 63 56 5d 62 60 66 47 32 21 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0f 2b 3c 59 60 70 84 8d 8e 7b 6b 65 59 56 5e 65 65 64 63 62 69 70 6d 6e 74 72 71 6c 68 74 71 72 71 6b 6c 71 72 6d 6c 73 6f 68 6b 69 6f 66 71 67 6b 65 65 6b 6a 62 62 6b 66 6a 64 64 6b 67 6e 6c 6f 74 6c 6a 77 6c 73 71 68 66 72 6e 71 73 63 6f 75 78 76 72 7a 6c 74 73 6d 76 80 78 7f 8f 8a 91 8c 98 95 82 7f 73 4f 13 0a 06 05 03 00 06 05 03 00 06 05 05 00 06 09 06 00 06 05 03 00 06 05 03 01 06 05 05 05 10 4b 6d 6b 79 75 77 6f 73 75 7d 75 7c 77 77 77 74 78 70 7d 7b 7d 7d 75 78 76 70 72 69 64 6d 66 63 6d 64 65 62 72 61 6f 70 6a 70 70 6f 70 65 68 62 66 61 69 6f 66 62 66 68 65 5d 60 5e 64 61 5e 59 58 57 54 56 5c 56 60 59 5f 5d 61 5a 5c 5f 5d 5f 5c 65 63 5a 61 59 5b 57 56 5a 51 54 57 4d 5d 4f 56 55 50 55 55 47 56 5b 59 59 57 59 53 5a 62 60 57 61 68 60 4f 35 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0d 0a 22 35 4b 6a 76 7a 80 85 7c 70 62 5b 62 5d 63 6e 62 65 6b 67 68 70 72 71 70 66 71 6c 75 78 76 6f 74 6f 6d 69 69 6c
 69 6d 6e 6b 69 68 69 6b 64 69 68 6e 6d 67 67 5d 6c 63 60 68 61 62 5b 64 65 6b 6d 78 6d 6f 6d 6e 70 6c 64 6a 6a 66 65 69 74 6c 70 79 76 68 76 76 74 76 76 81 7c 86 91 8d 87 91 93 95 87 82 75 57 1a 0f 06 05 03 00 08 05 03 00 06 05 03 00 07 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 08 15 44 67 73 76 74 70 78 7c 75 76 78 76 73 6b 70 76 78 78 78 74 77 7a 77 7f 7a 77 79 75 73 6a 65 6b 6e 5f 69 75 67 6c 64 65 6e 66 6b 73 6a 74 71 6d 69 6a 6c 75 73 64 5c 6c 67 62 62 59 65 61 5f 52 60 5d 56 5d 57 58 57 57 59 5d 62 5b 5e 5e 64 5d 60 61 64 5e 59 65 58 51 50 58 5a 54 58 4e 54 55 55 5d 58 53 55 4f 5b 52 50 5b 5b 62 5c 5c 57 54 53 5f 5e 5f 41 21 19 07 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0b 0f 16 2b 3d 59 70 7a 87 8e 7e 69 5a 5e 56 5f 5b 61 5a 69 61 69 73 6e 6f 6f 69 67 6c 66 74 72 6d 5f 62 6c 70 68 66 6f 6a 6c 65 62 66 6b 62 60 65 65 67 5d 6a 63 72 67 60 5d 6c 5e 63 61 62 68 6c 6f 67 75 6a 6f 74 70 6b 69 68 6a 6a 6e 6e 68 6f 6b 75 6e 6c 74 75 70 6f 79 7d 76 7e 83 89 86 84 86 89 8d 7c 7f 74 57 1a 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 03 06 05 03 05 11 34 62 6b 72 71 70 75 6f 76 6b 7c 6c 6b 6e 70 78 76 79 79 76 7a 81 78 83 83 75 7d 79 75 72 6e 6c 71 72 69 6e 66 6a 66 6e 71 70 72 75 68 6d 6c 67 68 66 6d 70 70 6c 6a 63 65 62 5e 60 61 60 56 53 5a 56 5d 5b 54 57 5b 57 5d 5e 60 56 59 5c 60 5f 60 57 5f 5f 60 5c 53 4e 52 57 4f 4f 53 4f 58 5b 51 50 51 49 54 48 4e 4f 54 5d 56 61 53 51 55 55 5c 5e 5e 49 38 22 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0a 0b 13 21 3f 5d 6d 71 91 8b 7d 6d 5c 57 58 60 5f 5d 62 61 64 62 68 68 69 6b 6d 6f 67 68 6d 70 70 6a 70 72 61 6a 68 6b 74 69 66 65 63 68 66 64 69 69 61 69 5a 70 66 64 66 60 5d 65 5d 58 66 60 63 65 72 74 75 7a 7d 7a 79 71 6d 68 62 61 69 6d 70 6f 6d 6d 6d 70 73 6a 76 70 7b 7a 7b 73 77 74 73 85 87 84 7f 82 77 59 1b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 10 05 00 06 05 03 00 06 05 03 01 06 05 04 06 10 30 65 67 74 70 67 76 77 76 79 71 77 70 71 77 73 75 7b 7b 7c 7c 84 80 85 7d 87 7c 77 7c 7e 77 77 76 74 76 72 77 78 6c 70 6b 6e 6e 6b 6c 73 6e 6b 70 76 75 7d 75 78 78 6b 65 64 5f 59 63 5e 53 5e 59 57 53 56 5b 55 58 57 5c 5e 5f 68 5c 5c 5c 59 56 5a 6c 5b 5c 59 5f 5a 54 55 54 57 51 51 51 56 51 5d 4e 48 54 4e 55 5a 5d 5e 5b 5d 61 54 59 5a 53 56 58 46 32 1e 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0c 21 3d 50 6c 77 80 8e 7b 71 5d 5d 58 5b 63 61 62 63 57 5f 65 75 66 72 70 6e 6a 66 72 6d 6a 6a 6c 68 6b 64 5e 6a
 6a 5c 62 60 62 66 59 5d 66 63 6a 6b 62 60 66 5b 61 60 5c 68 5f 5d 63 56 66 65 68 75 79 89 8f 87 83 75 74 6c 65 6a 68 6d 6b 69 67 6b 6f 68 72 71 76 79 79 71 74 75 6e 77 75 84 85 87 78 7c 70 58 25 0c 06 05 03 00 06 05 03 00 06 05 03 00 07 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 2a 61 69 6f 68 73 6e 70 70 6f 7d 6c 73 62 6b 73 71 75 7b 82 7f 7f 83 81 7f 7d 81 82 7a 7c 78 7a 81 77 72 6d 6f 71 6f 75 75 6f 73 7b 75 77 6d 72 6f 74 6e 76 79 71 7c 6f 6f 64 61 64 5b 64 59 5e 5e 57 57 55 53 57 5c 59 5b 5e 65 5d 65 5e 5f 54 56 61 62 67 62 5d 60 53 54 50 4f 51 5c 56 54 59 54 52 4e 47 56 52 55 4e 5b 5c 59 5a 5c 59 57 53 52 57 4e 3d 25 17 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 07 12 19 28 46 61 75 81 81 77 6b 5d 5a 5c 5b 5e 61 65 64 63 61 63 63 60 6b 6a 68 67 60 61 6f 61 63 69 64 62 60 66 66 62 65 5e 5d 59 5b 5b 60 5d 5f 55 67 61 5b 5d 61 5a 60 59 62 56 5c 5f 68 65 66 71 78 7d 7e 8b 84 7c 79 66 61 66 5f 5f 64 67 64 67 68 66 73 75 73 75 72 74 70 6e 6a 71 6e 71 76 7f 84 7b 7e 70 5b 1e 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 31 52 63 76 72 69 71 69 69 6a 6c 72 76 74 6e 7a 6f 7a 7e 7e 7c 7a 7d 78 76 7e 75 78 75 72 7b 75 7c 79 70 71 7a 6d 78 72 6e 75 72 75 73 6f 72 71 72 6d 60 62 73 6f 73 70 72 66 5e 67 65 5a 62 5a 57 57 59 54 50 5a 5c 5f 5e 60 56 55 5f 58 5f 5d 5c 5c 5c 53 60 58 60 5d 56 5b 55 5a 5e 57 5a 57 4e 4e 4d 50 59 55 4f 4d 59 59 5c 58 5a 5d 55 50 49 50 3f 29 1d 07 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 06 06 07 09 0d 1d 24 42 56 66 85 7f 76 6a 5b 59 5b 62 61 5f 55 5e 5e 5d 62 63 66 63 70 64 68 6c 68 64 62 6d 69 69 6b 5c 67 67 64 61 61 5e 5c 60 5a 5e 61 5d 66 5c 5b 5e 63 5b 56 5d 5f 60 5a 5c 5e 61 5d 60 6d 75 84 85 8a 86 80 74 64 64 62 65 69 66 6d 61 68 65 64 6c 71 73 6d 6e 6e 6e 63 75 6d 6d 77 71 77 74 7f 74 78 5b 1e 03 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 05 04 09 2d 59 61 6e 6b 6a 5e 6f 6a 6d 66 6d 70 65 73 78 77 6d 73 79 7c 7a 77 78 6e 73 79 72 71 69 78 72 72 73 71 6d 73 77 75 77 73 76 76 7b 76 66 7a 72 6c 6b 62 5b 6b 66 67 6f 70 64 65 6b 61 5d 62 56 5a 5c 5b 57 55 5e 58 5d 5b 57 5d 56 50 60 62 5b 5b 5c 61 5e 5d 5b 59 59 56 5d 53 5f 52 5a 54 5a 53 52 50 56 57 54 4d 56 56 5c 5c 57 5b 48 58 55 4b 4f 2e 22 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 03 0a 0a 17 17 2a 4a 6a 77 8e 7c 64 63 5f 5a 56 5f 5d 5c 5d 58 5d 59 58 6b 67 6a 68 5e 60 69 66 6f 69 6a 68 61 69 6b 6a
 6a 63 5f 64 67 60 5c 63 61 62 5c 5a 61 63 60 6b 61 5f 5b 5e 61 5c 57 5a 62 66 66 74 7a 82 87 7f 77 69 5f 6e 60 6b 63 69 6c 69 67 67 69 69 72 6d 79 71 6c 69 6e 6b 64 6c 73 70 7d 7c 6b 79 72 60 30 0a 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 01 0a 25 52 5f 67 61 61 69 68 6a 69 71 6d 72 69 6f 71 71 77 78 72 7b 7e 71 74 72 6f 70 6b 6c 6f 75 62 79 68 74 6e 76 72 75 77 7b 78 6f 76 78 71 6f 6c 67 64 63 5b 5b 60 65 70 67 74 70 67 6a 63 64 53 56 65 58 58 51 5c 5e 5b 54 5b 58 61 5f 55 5b 5d 53 5e 65 54 5f 60 5a 5d 4d 59 5a 5f 55 58 53 5b 58 51 4f 59 50 54 58 58 5e 5a 5e 5a 56 57 54 52 46 44 2e 15 0e 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 03 02 0c 09 1d 24 3e 5d 75 7f 75 68 5f 5a 54 56 5e 5b 58 53 5e 60 5a 54 59 61 66 67 63 61 68 6c 64 65 69 5a 5f 5e 5c 63 61 66 60 61 5b 58 58 62 64 54 63 5b 5a 65 5e 63 64 5e 64 5f 52 62 5d 5d 57 5f 69 68 6c 71 78 72 72 6a 68 6b 65 71 71 6b 72 67 66 6d 70 6d 71 71 73 68 71 66 65 6b 72 6f 73 6f 75 71 79 6d 72 66 35 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 05 06 1b 44 5c 63 62 66 5f 62 69 6c 67 6f 76 6a 72 72 74 6c 79 77 7c 72 6f 6f 68 70 74 71 75 65 6f 69 71 6f 6c 6e 69 6b 6a 70 70 69 72 6e 6f 71 6c 68 6a 71 60 61 63 5b 60 64 60 62 6b 72 73 68 60 5d 59 5c 5b 53 5a 54 5a 56 58 5b 59 60 5b 55 58 5c 5f 5f 53 5f 59 52 5f 5d 55 5d 58 5c 55 55 58 56 4c 5e 50 56 58 53 5b 55 5d 5b 5b 68 53 5c 4f 47 47 3c 24 1c 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 06 00 06 0c 0d 20 39 58 71 78 82 6d 5d 54 57 58 5f 61 56 5b 53 5f 59 56 5b 68 63 65 65 64 69 65 62 62 65 64 60 61 61 64 60 64 5f 54 5b 5d 64 5f 56 61 50 5d 5d 5c 68 64 62 5e 60 5a 52 58 5c 58 59 60 66 68 66 6c 74 73 6f 6a 65 69 6c 6f 79 70 6b 6b 68 6b 70 6e 65 73 74 62 6a 67 6b 65 68 6d 71 73 76 7b 72 7a 66 64 2c 09 06 05 03 01 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 1c 43 5f 60 64 5b 67 68 68 6b 6a 6d 66 68 75 76 6d 6b 68 75 71 6b 72 66 69 69 70 72 72 6d 6b 6a 78 67 6d 69 71 69 6a 67 78 71 6f 75 64 6d 6c 69 6d 69 66 5f 65 66 62 66 64 5f 69 67 72 6a 6d 69 62 5d 56 59 5d 54 5a 56 57 5d 51 5b 53 59 57 65 58 59 5a 5e 56 64 63 5a 5b 4e 58 54 55 57 55 56 55 54 4f 5c 56 54 50 56 56 62 5f 64 5c 53 55 4a 4c 2d 1e 1a 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 04 04 13 0b 0d 1c 2b 43 65 78 85 6d 63 5a 55 57 5e 5b 53 59 61 5c 5b 61 59 59 62 62 64 60 68 60 64 66 64 5e 63 60 65 63
 67 5b 5d 58 64 58 52 5d 56 5d 61 5f 5c 62 5b 54 60 5d 5d 5c 5d 57 5c 54 61 63 6d 64 66 6b 61 65 5a 5d 5f 68 67 6e 6d 65 67 63 6a 6a 70 6e 71 6e 69 67 6a 63 6f 66 6d 70 6d 70 75 6f 6b 70 6e 64 2f 0a 06 05 03 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 4a 5b 67 69 5c 69 64 5e 6c 76 68 66 66 6e 6d 66 6c 6a 72 70 70 6f 6f 70 73 71 6d 75 70 6c 6e 6f 6e 70 6e 67 6f 70 6d 70 72 66 63 70 6a 6e 6d 65 66 68 69 6b 6d 6f 6e 65 60 64 6e 72 73 76 67 64 6c 66 60 4f 51 56 57 57 59 55 5c 58 5d 6a 5a 54 55 5e 5e 64 56 61 58 51 5d 52 5d 51 58 4c 56 54 51 57 57 5b 56 55 55 5a 62 5a 5e 53 51 4f 4b 46 2b 19 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 06 0e 0e 1a 23 35 55 6d 7d 6f 59 61 57 52 5e 5b 58 56 54 5f 55 58 5b 63 60 60 5f 5f 66 65 62 63 5f 62 58 5c 5c 66 5c 5b 5c 56 5b 5c 56 62 59 5c 62 5f 5a 50 62 5b 59 58 58 5f 5c 52 58 59 59 63 63 64 5b 61 67 5f 5e 5e 54 58 6c 65 6a 61 65 6b 72 70 6d 66 6c 69 6b 67 66 69 69 63 6d 6e 6b 6c 70 67 69 6a 6d 62 3a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 11 40 5d 63 62 60 68 64 6a 66 6e 67 65 66 6c 6e 63 6c 66 66 70 69 69 6d 64 61 6f 6d 71 62 76 68 74 6a 6c 69 67 62 6a 6e 68 6b 6d 6f 6d 68 74 67 64 72 66 67 71 6a 6a 66 67 6a 5d 66 64 6e 73 73 68 61 63 5e 5b 51 53 53 58 59 5d 5a 57 5a 50 5c 55 58 60 5d 5a 5d 5a 5f 54 53 59 58 59 54 56 5d 51 4f 57 56 5c 54 53 53 52 5b 60 5e 57 5a 50 54 34 28 11 12 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 05 0b 11 16 24 38 5b 69 75 62 56 5d 4c 5b 57 59 53 53 57 54 5c 62 54 5d 5b 5c 65 5d 64 61 5d 61 63 5e 61 63 63 5c 60 5b 54 5a 53 56 5a 56 60 58 57 5d 57 5a 5b 5d 60 5d 5e 4f 5d 52 58 63 62 63 61 5a 5d 55 58 58 4d 5d 5e 5c 5b 62 57 59 5e 62 66 6f 5f 64 61 63 5f 62 66 63 66 65 6f 6a 5f 6c 6a 66 6a 64 5e 39 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 41 59 68 63 60 64 5d 60 65 67 60 61 67 68 64 66 61 6e 63 66 62 65 66 64 66 6a 6f 6a 6c 6e 6a 6a 6d 6c 65 6b 63 71 68 6a 69 64 69 68 6b 60 63 65 65 66 5d 63 60 65 63 5c 6b 59 66 6d 62 6e 68 6d 65 61 59 55 57 5d 54 53 56 5b 57 5d 56 54 55 57 5a 5d 5d 61 53 56 4f 51 55 52 59 53 55 55 57 54 56 51 55 54 55 56 53 51 58 58 53 4e 4b 4e 41 33 24 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0f 09 11 0b 15 1a 20 38 51 65 6d 63 5b 59 56 57 52 59 58 54 59 60 5b 50 5c 5f 57 61 61 65 6d 62 63 65 64 5b 5f 5e 5d
 58 5e 5d 63 5f 5d 59 59 59 5b 57 5c 5f 56 58 5a 60 61 59 5c 58 59 65 5b 6c 62 66 60 52 55 54 5a 59 50 53 58 58 5f 56 59 61 5e 5b 67 66 5e 60 62 67 61 67 64 65 63 71 67 67 68 6d 6e 68 62 62 52 3f 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 0d 40 55 62 5d 62 5f 64 60 64 5f 62 62 63 64 64 5a 68 60 6b 6a 61 67 6b 65 6a 6b 64 6e 67 66 6b 66 68 66 69 6c 66 66 66 68 64 6a 68 68 62 5a 66 5c 62 67 62 61 5e 64 64 66 5e 64 64 5c 66 6d 66 71 65 5f 5f 5d 5d 57 57 5d 58 5a 57 59 57 5e 51 5d 5f 58 64 5d 58 5d 5c 5e 5c 54 5f 5a 53 5e 55 5b 5b 52 57 54 51 56 58 5a 61 52 55 56 4d 4f 3b 2f 17 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 0b 10 12 0c 18 1f 35 47 60 64 5f 5c 5b 56 5a 57 55 50 52 5c 55 4e 55 56 5c 60 5d 5b 5e 62 5f 62 62 67 5e 64 60 5e 5d 60 52 5b 59 5c 55 59 57 54 51 53 53 5f 59 5e 5a 59 5b 5a 5c 5c 61 63 63 64 6b 5a 4b 4c 55 57 4f 53 57 54 58 54 5e 58 5d 5e 5c 60 5d 61 65 63 65 60 62 64 63 69 66 64 63 6a 6d 67 60 6b 61 5e 3b 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 34 5d 5b 63 62 5e 5e 54 61 5c 61 64 60 64 66 67 65 63 61 61 5f 6a 5d 62 6b 6a 67 64 61 6a 63 69 67 5f 66 62 60 65 65 60 61 60 62 64 65 65 5e 5d 62 5f 5d 5e 60 5f 62 65 5d 65 59 5e 60 67 65 73 62 62 60 58 57 57 5d 5e 5b 58 59 5b 59 56 5d 62 5a 5d 60 66 5e 59 59 57 62 5d 56 56 51 52 5a 55 57 54 53 4f 55 59 55 52 58 5f 58 4b 4d 41 3d 2d 11 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 0d 05 04 11 0f 19 26 32 58 5d 60 56 53 54 5a 5b 56 5b 51 52 5e 50 51 5c 59 5b 57 5a 56 56 64 64 5a 66 5e 60 5c 61 5e 5a 52 57 59 5a 4c 5a 52 67 52 53 5d 65 59 56 52 5b 55 5d 60 5b 64 61 67 62 62 45 54 50 58 59 4f 4f 4f 5e 52 51 56 59 61 5b 58 60 5d 65 5a 66 67 5e 60 66 5b 67 62 65 6a 67 66 67 64 5e 63 5d 3e 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 32 52 5b 5e 54 5e 59 5b 56 5a 5d 5c 50 63 59 5a 62 62 60 62 57 5d 62 64 68 63 66 6b 65 60 5c 65 5f 67 6a 68 67 63 69 62 6f 5f 65 67 61 61 5d 5e 5d 60 64 64 53 55 5c 57 60 55 65 61 5f 66 6d 6c 64 5f 55 5a 53 58 5a 57 5b 58 58 5b 54 57 57 54 5e 61 62 69 56 5d 57 58 5c 56 5f 5f 52 5a 55 59 58 55 51 56 5d 54 57 52 56 4f 4e 47 44 42 31 1b 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 06 11 15 13 14 1f 29 39 44 55 57 5c 55 58 5a 5a 59 57 52 5c 5e 58 52 59 54 5d 5f 59 60 5f 5f 60 61 65 57 59 58 5f
 5a 5f 5c 5a 57 5a 58 63 54 53 5e 5b 53 57 59 5f 5b 5e 55 66 62 69 63 5b 64 5c 55 58 55 55 58 59 58 52 4a 54 4b 55 5a 56 59 54 59 5a 56 5f 5a 60 60 61 64 67 5d 6c 65 61 62 5f 6a 63 64 59 5f 55 40 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 29 4d 57 59 5a 58 53 56 60 65 54 55 54 5f 5e 57 5c 5c 5d 64 5c 5c 5c 61 63 5f 5a 65 61 6a 60 63 62 60 63 69 64 62 66 63 62 61 60 63 5e 5e 5c 62 5c 5d 62 63 5d 5e 63 5a 5b 52 61 5d 58 5b 5d 68 6c 64 63 5e 57 57 5b 54 55 5f 5e 5e 59 59 5a 5d 55 5c 62 62 5e 5f 56 59 5d 55 55 5b 57 5b 50 53 5a 51 53 58 5a 52 54 59 51 54 53 46 45 3e 26 1a 0a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 0c 0d 0c 16 17 19 25 30 34 4f 5a 56 4f 57 60 5b 55 59 55 53 54 5b 5e 52 5c 5e 54 57 57 62 5e 67 5e 5e 5d 59 5f 59 5a 61 5d 59 59 50 52 5e 55 5b 56 5c 57 5a 5e 56 5f 5a 58 60 5e 64 64 62 5f 55 52 5d 5a 56 59 52 58 58 54 56 57 4e 51 54 5c 58 5a 5d 51 5c 59 58 62 5d 5f 60 52 62 63 66 57 61 66 60 62 5b 58 55 39 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 25 50 51 57 52 55 56 52 5a 53 52 57 55 5e 5a 55 54 5f 55 60 5e 5f 5e 60 67 61 61 64 65 60 5c 64 64 69 67 64 63 66 64 60 5e 60 61 63 5d 5b 5a 5b 5a 5f 5d 5e 5a 58 63 61 5f 5b 5f 59 56 5f 5d 61 6d 62 5f 58 59 59 50 59 5c 56 5c 55 5c 59 5c 5b 5b 66 61 66 57 54 5d 5a 54 5b 5a 5e 4d 5d 61 55 57 55 55 50 4c 51 5a 5b 55 53 51 47 3b 2f 25 0d 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 07 09 11 11 14 28 2a 3b 44 52 59 53 5c 55 51 59 54 53 5d 53 58 4a 4d 59 53 62 5c 5c 54 5a 59 59 5d 57 5c 59 60 54 61 55 5d 53 50 53 53 52 54 5a 51 58 53 4e 62 58 5e 62 67 5e 64 5e 5e 5b 57 4d 5c 4e 50 52 55 4f 50 5a 54 5d 4c 51 57 53 56 51 4e 4f 54 5a 56 61 58 5f 5a 55 5f 59 5a 5b 5f 64 62 5b 54 55 56 44 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1a 49 4c 54 56 58 56 4f 52 59 4b 60 4d 56 52 51 57 56 59 5e 5e 58 5d 58 5b 5c 58 66 62 61 64 61 68 60 65 64 64 64 64 5c 5e 5c 5d 68 5f 5a 61 65 54 5a 60 61 5c 5d 60 5b 5a 59 63 5a 57 5a 5a 65 65 64 67 60 55 57 63 58 5e 5e 5c 5c 50 58 58 57 5e 5b 56 64 51 56 5f 5a 5a 58 56 5e 5a 5e 5b 4e 5d 4a 50 56 51 53 56 51 55 51 4e 47 37 2f 16 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0f 15 14 15 22 32 36 43 4f 57 4e 55 59 50 5a 54 53 5a 56 60 4d 55 56 54 5e 5d 55 52 62 58 55 5b 57 65 5f 63
 52 59 56 5a 5c 59 52 57 5c 56 5e 58 58 5d 5e 5c 5d 5a 5f 64 66 5f 57 62 5d 57 55 50 55 55 59 4b 54 55 4f 55 4b 50 55 56 5a 50 51 4c 55 54 54 57 5e 59 5c 5c 57 60 61 57 5b 60 5e 5c 5a 5f 60 58 3f 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 3e 4f 58 51 58 4c 57 58 5a 53 52 52 59 5a 58 58 57 5f 5d 62 5d 57 63 57 5b 5b 60 5c 5f 61 68 61 61 60 5e 68 63 5b 60 5e 58 60 61 5d 56 5d 61 68 61 5e 5d 5c 5a 65 66 5e 5b 53 5d 5c 5b 5c 65 65 60 64 56 52 5b 5c 52 58 60 53 60 5e 62 5c 5f 5f 64 5b 64 5b 5a 61 58 5c 5e 5b 60 57 58 60 58 5d 56 57 53 4b 4d 55 55 4d 55 4c 44 34 21 14 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 03 11 1f 21 23 27 40 47 54 56 50 55 53 54 55 58 56 4a 4e 55 59 56 56 4e 56 55 5d 55 61 5a 60 5f 5f 5e 56 5b 5d 57 58 5d 56 4e 58 53 53 52 5a 5a 54 5c 5d 60 5d 66 5c 5b 5e 5c 59 59 57 56 54 51 4e 56 53 5a 54 4d 4b 50 53 5a 53 55 51 56 52 52 55 53 54 5b 52 59 61 59 59 5a 5a 58 5b 5e 64 57 5b 59 50 48 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1b 45 45 4b 4b 57 52 4b 50 54 51 51 54 55 5d 50 56 59 51 63 5b 58 56 61 5c 5d 59 5b 5e 60 5c 5e 5f 63 60 5b 64 61 5e 63 5b 5f 5e 65 5c 5f 56 63 60 57 58 5f 5c 53 59 5a 57 55 61 5e 5d 59 5a 64 5f 5f 65 5a 4e 4f 5c 5a 5c 57 5d 63 52 5f 5a 5c 5e 68 61 66 57 5d 50 53 62 51 54 54 59 5b 55 54 5a 50 55 51 4e 4f 51 50 57 44 4e 34 2c 1c 0d 10 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 09 0c 0f 10 17 1e 22 32 37 38 48 4d 52 4e 4d 51 58 58 51 5b 57 59 4f 5b 57 51 52 5a 5e 57 57 61 64 56 5b 59 53 59 55 57 57 50 52 5b 53 5c 5a 57 55 5a 5b 57 5e 61 61 64 5a 51 5f 5d 59 62 5d 53 52 53 54 55 5a 59 46 4d 52 53 47 4d 4e 4b 53 55 51 53 53 47 54 59 56 57 54 58 58 56 5e 52 5b 52 56 55 57 52 50 41 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 3e 44 4f 4d 4d 53 4e 55 52 4f 47 50 53 54 54 56 52 5d 54 5c 5e 58 56 59 56 5a 55 61 58 5d 66 62 65 5e 62 60 54 61 5d 52 59 59 57 52 5a 56 56 58 58 59 57 5b 5e 5b 50 5c 5d 5b 53 5b 60 55 6a 68 63 60 64 5b 57 58 54 5b 59 5a 5b 55 5d 5f 60 5c 5e 5a 5a 5f 55 5b 55 55 55 56 5a 55 54 58 55 5d 57 4d 53 52 4f 4a 50 4a 4d 3e 2e 18 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0a 15 13 14 21 2b 30 38 4e 49 4e 53 4b 4e 54 52 5a 56 57 5a 53 54 49 52 52 55 5c 5f 5a 5d 5e 64 59 60 5e
 56 5c 61 4d 57 53 58 5b 5b 54 5d 5e 61 5e 5a 5e 5f 60 61 5e 55 57 5b 51 5a 54 54 50 53 50 5c 44 2a 3b 57 55 4f 4c 47 4d 50 53 52 4b 47 4d 4c 50 58 53 5a 53 4f 51 55 50 5c 53 54 55 59 5e 4e 4d 4a 20 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1d 3f 53 56 4d 51 4b 4c 54 4e 54 53 50 4e 56 52 51 54 53 5a 52 59 5e 5b 4e 5f 61 58 5a 60 5e 61 58 5f 65 5c 59 5c 55 54 5c 55 5f 55 53 4d 4f 59 5f 53 53 62 56 5a 5e 5c 5c 5d 5a 59 5a 58 5c 68 5f 62 61 5e 5e 56 58 54 54 54 61 5d 5f 5d 60 65 5c 56 5e 5a 58 57 5b 57 58 54 57 5d 5c 58 5a 59 57 4f 51 4b 4b 57 4c 4e 4f 42 40 1e 13 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 08 11 11 14 1e 1b 25 36 34 42 4a 4b 50 54 4f 56 4e 53 59 58 59 5b 53 5a 56 5a 59 59 5a 5e 59 5b 5f 5a 5e 59 59 5a 59 5b 59 5a 59 59 59 5c 62 5b 67 5f 57 61 65 57 5f 56 5d 5d 58 50 5d 53 50 58 4f 54 50 4d 54 55 57 4d 4a 4f 4f 4e 54 4d 4c 51 4b 4e 50 49 4d 4d 4d 55 5b 5c 56 60 55 5b 59 58 4e 57 52 52 47 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 32 4a 4a 48 4c 4c 4b 4d 52 4c 4e 49 52 55 46 54 54 52 58 55 5f 5d 54 58 53 56 52 57 5e 64 5c 60 61 5f 57 58 5f 64 5a 51 58 5c 58 57 59 5e 60 5a 59 5b 54 50 5e 5e 5b 54 59 51 64 54 57 5f 6b 5b 63 62 5f 61 59 60 5a 53 5a 55 66 54 5f 51 63 5c 5e 66 5f 5a 5c 5d 52 57 55 5b 56 53 60 55 52 56 54 56 4a 51 52 49 54 51 46 3e 23 13 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 04 0c 10 16 21 23 2c 2f 41 45 49 55 54 4f 56 54 4b 55 54 59 58 5b 5b 58 53 59 55 5b 4e 5b 5a 56 5f 57 59 58 55 56 53 57 60 55 58 5c 58 5a 55 60 66 5c 5f 61 5c 5a 54 59 5d 55 58 59 59 51 57 52 4c 5a 52 4c 49 4a 51 44 4b 4f 45 52 52 4f 50 49 50 4d 50 56 52 51 4f 55 54 4f 59 4f 51 53 4d 53 59 49 53 49 27 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 33 49 4d 49 54 52 44 52 48 4c 55 49 51 4b 50 4d 54 51 5a 4e 59 53 54 56 58 5b 57 56 61 54 5e 5e 5e 5d 5a 50 56 56 58 57 54 5c 50 56 52 54 52 5a 5e 52 58 4b 58 5d 5c 57 57 57 58 54 55 58 63 59 5f 58 59 55 60 52 5d 51 5b 5f 58 5b 5d 59 5c 5b 60 60 5e 54 57 55 56 56 4d 58 58 52 5c 4f 56 53 4b 49 54 49 4b 4c 4c 4c 34 29 15 10 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 15 1d 2f 1f 25 2b 3e 40 48 4e 4e 53 4e 4e 4d 56 4f 58 52 59 50 4b 57 59 60 58 5d 59 55 59 50 5e 5c
 52 57 62 53 5d 56 5d 5a 59 5e 5c 5c 58 63 63 62 57 58 57 62 4f 55 4e 53 57 5b 4d 49 51 48 4f 52 50 4a 4c 4f 48 47 47 4a 46 4f 55 54 4d 4d 44 4d 51 56 53 54 50 58 4e 54 57 50 53 59 54 50 56 4a 43 23 06 05 03 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 30 46 52 49 4b 47 48 4b 51 4c 4b 46 50 4f 54 4f 51 4c 4f 56 57 57 54 59 5a 5a 54 55 57 52 56 56 57 52 58 58 5b 59 56 54 56 58 53 4f 51 55 54 4c 5a 5a 58 53 57 53 51 58 5c 53 57 5e 5d 62 5b 5e 60 5d 5d 53 50 5a 5d 58 5a 5e 5d 54 5f 5a 5d 5f 61 61 64 5d 51 55 4f 56 55 57 57 57 55 51 53 4f 4f 50 4b 4e 57 49 48 3e 35 25 1b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0c 15 0e 13 22 28 2c 34 3e 40 43 4e 4d 52 4d 50 55 4d 4c 56 53 55 54 51 5c 56 5d 52 5b 59 56 5c 54 5a 5b 5a 55 5d 58 59 58 5d 64 60 5e 5f 66 5e 5e 5d 5f 5b 60 56 59 5a 56 56 58 55 4a 52 54 50 4f 50 4e 50 4f 59 50 48 51 4c 57 5a 4b 52 50 4c 4c 56 49 47 46 54 56 5a 59 58 54 56 50 52 55 46 4d 51 4c 44 2e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 2c 3c 50 51 51 45 4d 51 4e 41 4c 4b 54 49 58 4d 50 52 64 54 51 55 59 4f 53 52 56 58 5e 5b 60 52 59 5e 57 59 55 54 55 56 57 52 52 53 4b 55 52 52 5c 53 50 54 5a 4d 56 5b 55 62 57 52 5b 59 5f 53 5c 5b 59 57 5a 5c 57 60 60 65 62 58 60 58 61 5b 5f 59 59 5a 5c 58 5a 59 57 55 53 53 57 51 4f 4f 48 4a 50 55 54 4c 43 4a 37 21 17 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 10 1f 1a 25 35 36 3f 47 4a 4a 44 4f 45 4f 57 52 58 53 5c 53 5a 55 59 54 59 56 5d 5d 58 5b 55 61 5d 54 54 59 5a 5e 60 61 57 61 64 5e 5e 5e 5a 59 5f 58 64 5d 59 5b 58 54 53 56 59 5e 4a 45 4c 49 51 50 4d 4b 49 4c 4d 4c 5a 4c 47 4b 4d 54 52 53 4d 52 57 50 4c 4d 4f 4a 4e 50 56 5b 52 54 47 4c 46 2e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 22 48 4d 49 41 4a 4a 4d 49 41 49 4c 56 4b 4b 4c 4c 4e 52 52 52 4e 59 4f 52 56 5b 59 5f 57 55 4e 59 4c 58 5d 59 5d 58 4e 5c 53 4c 55 53 58 57 58 55 53 59 5a 55 5e 57 50 52 55 5c 4e 53 51 5e 58 59 59 55 53 5a 56 5a 5b 5c 5d 64 5b 5d 5e 58 64 5f 57 61 53 5a 54 58 5a 57 4f 5d 53 50 4d 44 4d 50 49 46 45 53 4d 46 40 27 1f 12 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 13 13 19 27 2f 36 40 47 48 4b 53 59 4e 53 4b 4e 52 53 55 58 57 4f 5b 54 62 55 58 5a 5a 56 53 51
 52 57 5a 50 5d 58 5a 5a 5e 5c 5e 5e 56 5b 5b 5b 69 5d 56 61 59 58 5c 55 5e 4f 4b 4e 4d 4a 49 48 54 49 4b 50 52 49 4d 53 52 48 52 47 47 51 48 52 4e 4a 52 55 59 50 51 52 56 4e 4b 4f 4e 50 46 4d 45 34 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 2a 42 4b 45 47 43 42 42 47 47 50 46 57 56 54 4b 50 54 52 5c 54 56 54 52 5f 52 58 56 56 56 56 55 56 57 51 59 51 4d 52 50 59 5c 57 49 52 5d 50 54 56 4c 58 55 4e 5b 51 57 55 57 5a 51 5c 58 5b 5a 5b 61 58 54 55 56 58 5d 63 53 5d 58 5b 5b 57 56 5a 67 5f 5b 53 58 54 55 56 57 51 4d 4e 4e 54 4d 42 50 4f 4c 4d 49 3b 36 20 19 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 09 0d 10 20 23 20 28 3c 35 41 4d 55 4c 4f 52 58 4a 51 4e 5d 4d 4f 58 4f 5b 59 62 5f 5e 5c 59 58 58 50 59 5a 57 5e 59 5c 5c 5c 58 5b 60 57 58 61 5b 5e 5b 57 5f 61 58 60 60 59 59 52 53 4e 52 4a 4b 49 4d 49 49 4c 4d 4c 4c 50 4f 49 4f 52 4d 4d 4d 57 4f 53 4f 52 4b 5d 51 4e 4b 53 51 53 52 51 4e 4d 41 2c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 22 3b 49 47 49 4d 47 50 4f 47 4c 48 4b 4c 4b 52 54 56 4f 52 5b 54 58 4f 5e 5b 64 4f 50 59 57 50 59 56 5c 55 50 57 58 54 58 54 5c 51 5c 50 58 5b 56 58 52 5e 57 55 58 5c 54 57 51 52 5b 4e 5b 5a 57 65 57 4d 54 56 65 65 63 5d 5a 53 5f 5a 5b 5e 59 5b 5f 56 55 5f 57 52 4f 52 57 53 4f 52 53 54 48 52 4e 49 48 44 3c 33 22 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 17 13 20 27 2a 38 3c 3f 4c 4c 4d 55 52 50 4c 46 55 55 54 56 52 5c 5a 5d 5e 59 61 5a 59 58 5f 51 4f 60 58 5a 5d 5b 59 5c 62 5f 5d 64 63 60 5c 63 5a 55 58 57 50 5b 56 5a 53 51 56 51 4d 4e 47 4c 53 51 53 53 56 49 48 4a 4a 48 53 49 4d 48 4b 4d 4a 51 53 52 4c 54 49 52 4e 4d 4d 50 4f 4d 4f 4c 47 32 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 43 43 4a 4f 4b 4c 4a 48 4a 52 4c 4f 4f 4e 55 4b 51 53 51 59 56 5a 50 5b 57 5b 56 4f 59 55 50 4f 51 59 4b 5b 53 5c 55 58 58 55 57 55 4c 54 55 56 55 56 4f 50 62 5d 58 59 55 4f 55 59 57 56 56 50 4c 5a 56 64 55 5e 5c 5d 55 62 58 54 56 58 66 59 5c 63 55 50 53 4c 4e 4b 49 4f 51 50 55 5c 51 4f 54 4a 48 46 40 3d 2b 1e 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 0b 15 18 1f 27 32 42 3d 48 4e 46 50 4e 51 50 50 48 58 4f 54 54 5d 5c 56 5f 5a 60 5f 5d 5b 54 59
 60 5b 55 59 58 60 5d 60 5c 5b 63 65 58 59 5e 65 59 5e 5d 61 52 5d 57 56 57 51 51 55 50 4c 4b 4c 4a 4f 4d 4e 4a 48 4d 4e 4a 4a 4f 4a 48 47 49 4f 4e 49 4f 4e 4a 4f 57 4c 4f 4f 53 54 4f 54 41 4b 3f 37 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 44 3b 48 43 4a 51 46 4c 4a 4a 4c 4b 4b 4f 4b 56 4d 5d 47 53 55 53 55 51 53 51 51 58 54 50 52 54 4f 4a 4b 4f 59 52 52 52 53 4e 58 50 50 54 50 51 4f 52 54 55 5e 5d 57 50 4b 4b 4d 5c 56 58 5f 5a 58 5e 53 53 50 57 5a 60 5b 5c 5c 59 58 62 5f 59 5d 53 54 57 50 52 53 55 54 4e 52 52 51 47 52 4d 53 53 4b 44 3d 30 2e 19 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 11 10 1d 1b 28 33 3b 43 48 47 48 4a 52 4e 4f 51 4f 55 4f 52 5a 5a 5b 5b 57 56 5d 5c 5a 5c 5c 63 56 54 58 56 56 5f 5d 61 62 68 64 5b 55 61 63 62 60 56 5d 65 5a 53 5c 53 51 55 52 56 4f 50 4b 56 4f 4f 49 47 4d 4d 4a 4e 4e 4a 4d 49 47 4f 41 4f 4d 47 4a 51 50 53 53 4b 47 50 48 52 4d 50 4f 4b 47 3c 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 16 41 45 4c 44 4d 48 47 4b 4d 53 49 48 4d 4b 4f 51 4f 4f 4b 52 4d 54 55 55 5b 4c 52 59 58 5d 53 62 4a 4f 51 52 59 5a 52 50 55 4d 51 58 5a 59 58 5b 4c 56 54 5b 67 60 58 5b 57 5c 55 57 57 5e 5e 53 58 58 54 5e 56 5d 5f 60 5a 64 5b 59 61 56 52 5f 5a 5f 51 59 5c 55 56 58 4a 55 4c 55 4f 53 56 4d 47 45 40 4a 3c 32 2e 10 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 0a 13 24 27 33 33 37 49 44 42 49 41 4c 48 51 4a 4b 55 54 50 4f 58 5c 53 5d 5c 59 5b 56 56 61 60 62 53 5a 60 63 61 62 64 69 60 65 64 62 64 61 61 5f 5d 61 54 5a 58 51 54 51 4d 55 51 58 56 50 4f 4e 4f 47 49 46 49 51 4c 45 4b 4e 4a 51 43 4d 4c 47 49 4d 41 55 4a 51 4b 50 50 4c 54 4a 44 3e 41 31 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 37 49 45 4a 45 45 4a 49 47 4a 48 47 51 4e 48 4c 45 4f 4b 51 57 52 51 50 55 59 51 52 5a 55 52 5b 52 54 4f 56 50 5b 4c 59 58 4f 52 50 4f 58 53 58 5c 53 56 58 61 5e 50 57 55 54 57 58 56 54 5d 59 59 57 52 61 5c 57 60 5d 53 5e 5a 5d 5b 63 5b 56 5b 59 52 56 50 51 59 50 54 4e 4a 50 4f 4d 4d 4c 4f 49 49 45 36 38 20 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 03 19 1c 1f 26 35 45 41 41 49 4b 48 46 4c 4b 4b 50 4e 53 47 4c 4e 54 53 52 58 60 5d 5b 5b 57
 51 5d 55 5e 5e 63 66 69 68 6f 64 60 61 61 5e 5b 5c 57 64 61 58 59 59 51 4c 50 47 50 4a 50 49 4b 4c 49 49 4a 48 4f 4c 51 49 46 49 4a 44 4b 47 4a 48 45 4c 47 4b 4b 45 48 4b 4d 53 49 4c 4f 4d 40 41 2e 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 3b 4e 40 46 49 49 4c 43 3c 49 3f 49 47 4d 49 47 4c 4e 55 53 4e 56 57 51 50 4f 4d 52 53 52 56 52 47 57 4f 50 4d 54 52 53 56 54 50 50 59 50 53 54 58 58 54 55 51 64 53 50 54 56 4f 54 55 5b 60 5b 57 4f 55 51 5d 5a 58 5a 56 59 51 57 5b 5b 58 52 53 5d 54 53 4e 4b 49 51 43 4f 53 4b 55 4f 4e 46 47 46 38 42 3c 20 13 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 12 14 20 2b 31 3c 46 47 47 40 48 43 4d 44 49 4f 50 4f 56 4d 51 54 55 57 5e 61 53 57 59 52 5a 5e 59 61 62 64 6b 64 69 5e 60 5e 5b 60 60 5a 5d 5a 61 5e 5e 57 57 52 53 50 55 50 4e 50 53 48 51 50 4f 52 42 4c 4e 4d 4d 4b 52 4b 43 4a 52 4b 55 46 4e 4e 4e 4b 48 42 4a 55 50 51 51 4c 45 46 3c 2f 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 37 41 45 41 47 49 49 4b 4b 46 42 44 56 4b 4d 50 54 4e 53 4d 50 57 4f 50 51 50 4e 51 4b 51 4c 4e 54 45 51 4e 5a 59 4c 52 50 5a 4c 4f 54 50 56 51 5a 5a 5f 5b 57 56 55 52 52 53 55 60 5a 5f 58 51 5a 54 51 5c 56 54 5d 60 5a 5e 54 59 5d 5a 59 5e 55 5f 55 51 50 52 4c 57 47 5b 52 4b 4b 47 53 49 4f 4f 3d 38 34 1f 15 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 13 14 1a 31 33 38 48 49 44 41 45 48 46 57 4e 52 52 49 48 50 50 58 4f 50 5e 55 5f 60 57 5a 59 64 5e 6c 66 64 64 65 65 6d 59 5e 5c 5f 62 64 62 5e 5e 56 54 5e 53 52 56 52 58 4d 4d 48 4d 55 4b 4f 56 49 50 4a 47 47 49 53 49 51 45 47 4e 48 4b 51 49 4d 4e 54 4e 4c 4a 44 50 46 47 4b 44 4a 41 3c 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 30 3d 40 44 42 46 4a 50 49 44 43 4d 46 4b 4d 51 4e 49 43 54 4a 52 52 57 55 55 4f 53 4d 53 49 53 4e 4e 51 51 53 50 58 5b 52 56 57 57 5f 53 51 59 54 55 54 50 57 59 56 53 51 58 51 59 5d 59 55 52 58 55 58 5f 59 58 55 67 61 5e 5a 5a 56 58 55 57 52 56 5b 56 53 55 58 56 51 56 4a 58 51 50 49 4a 45 4c 3b 36 26 15 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 08 12 13 27 2a 37 4c 51 4a 4e 4c 53 4b 43 45 46 4f 44 4b 45 4a 50 4b 51 4b 54 4f 50 57 5a
 63 5d 69 64 67 68 5d 5f 5b 58 60 64 5c 5d 5a 5b 69 58 63 5b 5d 51 54 5a 52 56 54 4c 49 4a 49 49 4f 45 4b 4c 47 49 47 46 4a 51 51 4a 48 44 44 46 45 43 4d 49 49 52 48 45 45 47 3f 51 4a 46 3c 41 40 3a 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 32 42 42 42 44 43 46 47 4a 4c 4e 4e 49 4e 4d 4c 44 50 4f 47 51 4c 53 52 4a 4b 47 53 54 4c 50 52 4c 48 4d 50 52 59 4d 4c 58 58 55 4f 58 56 57 4c 56 54 4d 54 57 54 55 5f 52 55 57 58 4f 5c 52 5e 57 52 5a 5b 53 57 4d 58 5c 58 55 5c 5f 60 59 5d 4d 5d 5b 4f 5e 59 55 53 59 55 51 4d 4b 4d 4e 4e 45 3e 37 31 1a 0e 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 10 14 11 1d 2d 34 4d 4f 4d 4a 46 45 49 43 49 52 4c 4a 44 4d 4c 4f 49 4e 56 51 5b 59 56 56 5f 5c 65 64 5e 5f 61 5b 58 62 5c 54 5f 61 61 5e 5f 60 61 59 54 5f 58 57 57 4f 55 57 49 4d 55 4c 50 4b 4e 4e 4c 48 55 51 48 4a 4d 47 4b 4c 48 4d 47 4d 50 46 4d 51 47 4b 4d 4c 49 4e 47 48 49 40 43 39 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 26 41 47 3e 3d 44 41 49 43 40 3f 4d 4a 46 4a 47 4a 4e 52 55 49 52 52 4c 4f 4b 4f 55 4e 52 50 54 4e 4d 50 58 57 54 4c 59 56 51 59 52 5e 5a 57 59 4d 4e 53 4e 56 5a 59 5a 5c 55 5a 5e 59 5d 54 4f 5f 5d 5a 53 51 55 64 5b 58 54 5b 5c 5c 60 58 5d 5e 5f 58 53 58 63 56 53 56 4d 4f 4d 48 4f 4b 42 40 47 2f 29 21 0b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 00 0a 12 11 27 27 38 50 4e 4e 4e 47 45 44 41 45 4b 42 44 43 47 48 47 4f 4f 4b 4e 50 54 56 57 5d 61 60 66 5d 62 5a 5f 56 60 61 59 5f 61 5b 68 5b 5a 5c 67 50 53 61 56 59 60 4e 58 51 4f 47 4d 56 4c 56 50 49 4b 48 4a 50 4d 4d 48 45 49 46 52 49 4c 50 44 4d 50 49 45 4b 4a 4c 53 43 52 4a 40 3c 36 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 20 43 43 49 3f 4c 43 4b 43 45 44 47 50 4a 4c 49 4a 4b 4a 4e 51 54 4e 4d 4a 50 49 52 4f 52 51 51 51 4f 5a 5b 59 5f 57 57 5f 5a 52 4b 52 51 4f 51 4f 49 59 55 57 5b 56 55 5f 5f 4a 5f 58 58 5c 51 55 5a 53 54 57 59 5b 57 59 55 5d 59 5a 59 58 5f 65 61 62 5f 61 55 58 51 4d 4d 4b 49 49 4a 47 48 47 3c 2f 1f 17 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0d 11 14 23 31 40 4c 50 4d 3c 3d 3b 46 4e 40 4e 47 4d 46 42 4b 46 4b 44 45 45 50 56 55
 5e 59 5b 5c 64 60 5d 55 5c 5b 5d 5b 5b 60 63 61 60 5f 5c 5b 50 61 57 57 53 57 57 51 50 4d 56 4e 47 4f 4b 4c 54 4a 48 4f 4a 4e 4c 51 48 45 4e 50 4e 45 49 4b 46 49 4b 49 49 45 47 4a 46 4b 41 3f 3c 34 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 25 3b 3e 3f 49 46 46 47 45 46 44 47 53 45 46 50 44 4a 51 4d 56 4f 4c 50 50 51 44 4c 52 55 48 54 50 4f 54 51 55 58 56 57 58 59 58 4f 52 56 4f 5a 55 53 50 59 5d 58 60 59 5a 60 57 55 5b 5a 5a 52 59 50 50 5a 58 55 56 55 62 59 56 59 5b 55 5b 5f 5f 6d 63 52 53 59 49 4e 56 54 41 4d 49 49 4a 3a 3f 3c 28 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 05 00 0b 07 10 16 1e 30 3d 50 57 4b 44 3d 3c 43 46 4d 47 4a 41 46 45 47 48 4d 4d 4d 4d 4b 4b 53 5d 5f 5f 55 57 5d 5b 5d 58 58 5b 54 5b 58 61 62 5c 5d 53 62 55 5f 56 4e 4e 4f 49 51 4e 50 48 4f 4d 4a 4e 4b 50 4f 4f 4d 4c 42 52 45 4f 50 4e 4b 4c 4b 45 49 49 40 46 45 4d 4a 49 47 43 44 44 3b 3a 32 30 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 21 3c 3e 49 44 45 48 4e 42 47 3a 42 43 47 4b 49 48 53 4a 4a 47 4c 4e 4f 46 4f 4e 54 4c 51 4d 51 52 57 56 5a 59 60 56 55 62 58 59 4e 55 4e 4e 4f 50 54 4e 4d 55 55 62 59 5c 60 57 51 54 54 57 51 59 53 51 58 56 55 62 5f 5c 5c 5d 5a 5f 54 57 5f 5c 66 5b 5b 52 5a 4e 4d 49 48 48 45 48 45 49 3f 3c 2e 1f 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0c 08 12 16 1c 29 39 41 40 3f 42 40 44 45 43 42 48 47 44 46 47 45 48 4a 4f 49 48 4d 56 54 55 58 64 60 57 57 5a 5a 59 59 57 58 60 58 5a 5d 63 5a 5a 57 5a 56 59 54 50 55 4e 55 4c 4d 4e 4e 53 4b 4c 50 51 49 4a 4b 50 51 4c 46 52 47 41 4d 4d 4f 47 49 4a 47 3f 44 4b 48 49 48 40 49 40 3a 3d 3b 26 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 22 3b 3f 46 40 46 45 4c 3b 47 3c 42 3e 41 47 4f 47 4c 46 44 4e 52 57 4c 55 54 4b 4c 4b 57 58 56 58 53 53 57 5b 5c 57 55 5f 58 4f 52 4b 53 53 51 56 4f 4c 58 51 60 5a 5d 56 59 53 56 5b 5a 5c 5f 51 54 52 5a 58 5e 53 5f 5c 5d 5c 62 57 5d 5d 5e 5b 5c 59 52 51 50 4d 4e 4f 4c 4c 4b 47 45 41 42 35 2b 20 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 18 1c 2d 3d 42 3b 3e 43 43 44 49 3c 42 49 41 47 44 44 47 52 4e 46 51 4b 4c 56
 5b 55 5d 60 54 5a 5e 57 5c 5c 5b 58 5a 55 55 5b 61 5d 58 5f 5a 5d 51 4d 5e 53 55 4e 48 52 4d 4b 4f 50 48 4d 47 4e 49 4c 52 43 41 44 42 45 47 4d 41 4f 49 44 51 43 4a 52 48 4a 42 45 4a 47 42 3e 3c 3f 2c 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 3f 3e 3e 4b 3b 3e 40 3f 42 45 45 4e 48 43 4e 47 4e 43 49 4c 4d 52 4e 55 4c 4f 55 4f 51 50 5a 58 52 5b 51 58 57 52 52 4e 51 56 57 4d 53 4f 4d 51 4f 55 56 57 5b 56 5e 56 55 51 56 4e 58 52 4f 54 4d 53 53 58 53 57 58 59 58 55 50 5d 53 56 5e 5b 55 52 44 53 4b 40 48 4b 4b 47 46 4a 4a 44 3b 34 27 0b 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 10 27 2f 38 38 3c 41 38 3e 44 3d 43 48 44 42 42 43 49 4e 4b 44 52 3f 43 53 46 55 54 4f 51 59 51 5a 59 54 57 55 5b 4f 5c 5b 5d 53 5a 60 56 56 55 5b 54 56 51 48 4e 4b 4f 4d 4f 4e 4b 4d 4d 49 4c 4a 4a 4d 45 50 4a 49 51 47 4a 43 45 40 45 49 49 48 46 4b 43 49 48 41 3e 43 3c 42 33 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 18 3d 40 41 44 3f 40 41 3b 3b 3e 43 48 48 43 45 4c 45 4e 4e 58 4d 4c 4d 4a 4f 55 57 4c 4d 51 53 50 52 54 5e 58 51 58 53 5c 52 4f 4a 4f 56 51 51 5a 58 56 4e 55 53 51 5e 5a 59 57 56 51 5d 50 53 4f 50 52 57 53 54 59 60 5d 5f 4e 5b 4d 4e 4c 5d 56 52 4b 52 44 49 4f 4a 47 44 4d 4d 4d 44 41 3b 2b 22 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 06 0a 11 15 1c 27 37 3a 3f 3c 3f 3e 3d 44 40 46 43 44 42 4c 4a 46 4d 47 4e 4c 4e 4a 4e 4f 55 55 54 54 56 58 56 54 58 59 58 50 5f 55 5e 5a 51 5f 5a 52 59 55 52 5a 4f 51 58 44 4f 52 4b 51 51 4e 47 49 43 51 4a 4a 4b 4c 46 40 50 4f 49 4f 4c 45 4c 3b 48 4d 42 44 4b 4d 44 42 4a 45 42 40 42 33 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 15 3c 3b 45 4b 43 46 49 45 43 3a 46 46 44 4b 44 55 53 4f 4d 45 46 52 4b 53 54 4c 4f 48 4d 51 55 5a 53 54 54 55 56 57 52 53 4b 4d 50 59 54 58 4f 4e 51 53 59 5f 59 56 58 59 50 56 50 52 52 50 4f 51 55 53 59 56 53 58 62 60 60 55 57 55 4e 52 4f 4c 4c 49 4a 4a 51 4c 48 4e 45 45 46 51 3f 43 31 20 19 10 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 15 22 2b 3c 3b 35 3e 35 36 40 44 45 41 42 40 46 45 55 44 42 48 43 3e 44 51
 4a 52 43 4c 4e 54 4a 55 55 50 55 51 56 59 58 50 51 56 4e 50 56 55 59 52 51 4e 49 50 4f 4f 51 4f 45 50 4c 4c 45 4b 4d 46 4b 42 4d 44 47 4c 46 45 49 46 45 4a 46 4a 47 42 48 40 49 40 3b 45 40 41 41 3a 26 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 30 3c 41 40 49 3e 3f 3e 48 41 49 45 46 4e 48 4d 44 4e 4b 47 4e 4f 55 4a 47 49 50 4c 53 5a 47 52 52 5b 52 51 59 4d 58 53 49 4d 56 4f 55 50 4d 52 5d 55 58 5b 5f 58 59 50 55 50 49 52 4e 57 51 55 4a 51 58 54 4f 5a 55 58 56 5e 54 4c 59 4a 4d 49 4c 4d 4c 47 41 48 45 50 44 45 47 41 3b 3e 37 1e 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 1a 1a 29 3a 34 34 3c 3b 42 3b 42 3f 41 3e 47 40 47 50 47 42 45 41 4d 46 40 4b 4b 4f 4f 4b 56 4c 4f 53 4f 4f 4f 52 56 4e 4b 4a 4b 4b 55 54 54 57 45 50 4f 4f 4d 4b 4c 49 4f 4e 4b 51 4b 46 4b 50 48 49 4f 54 4b 49 47 4c 4b 42 47 47 4a 49 4e 4b 44 48 43 47 47 49 3b 40 3e 3f 38 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 3c 47 40 43 41 44 4a 41 44 44 4c 4d 48 41 4b 54 4a 4f 49 47 50 49 57 4a 50 4c 4c 55 53 51 55 45 4f 4f 4c 49 54 55 53 4d 4e 53 50 50 4a 4e 52 4c 57 54 54 5b 58 57 53 55 56 4e 4d 47 52 52 56 53 52 4e 4c 57 4f 52 5d 55 56 54 55 5a 47 50 4f 48 4b 44 45 49 43 4b 4f 3d 45 47 3b 43 39 3c 1a 1a 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0a 0c 1f 25 30 3d 39 39 38 3d 38 44 43 40 37 42 4a 43 46 4e 45 4c 42 44 49 45 51 4f 4c 4a 4b 52 52 53 4c 4f 4c 50 4d 56 51 4b 52 4a 54 50 4d 52 50 4f 55 5a 47 50 51 47 50 4b 47 49 47 4f 46 45 49 4a 4d 4b 43 44 52 49 4d 4f 52 4a 47 46 4a 4d 4b 41 46 3f 53 4a 48 40 3c 3e 38 3b 30 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 3c 33 4f 4d 3e 46 43 43 44 43 47 47 42 47 4d 4a 50 4b 4f 57 4b 50 52 48 50 4f 4b 56 4f 55 52 4f 52 58 55 5a 5b 55 4d 55 56 50 49 4b 4b 51 51 50 54 57 56 62 58 55 50 55 51 53 4b 4c 51 54 4d 54 51 52 57 53 50 59 5b 5d 50 52 52 46 46 47 44 4a 46 4c 45 46 40 42 41 47 48 42 47 48 39 30 22 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0a 0e 15 1f 21 31 33 33 3f 3a 44 43 3e 3a 42 3e 43 4a 48 4b 49 49 44 49 4a 40 50
 4a 50 43 45 45 53 4d 54 4d 53 43 4c 47 50 53 4a 50 50 4c 58 52 4a 4e 50 53 4c 50 4e 47 50 4a 53 55 4b 50 4e 46 57 4c 4e 4e 4d 45 4e 53 4d 41 43 4c 47 4c 4b 45 47 48 3b 4d 3e 41 44 45 4a 44 3e 34 3b 31 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 10 30 3c 4a 47 4c 4d 46 49 4e 44 4d 4b 50 51 4c 51 54 4b 4d 4b 4c 50 54 50 5b 4c 56 4c 4c 46 54 48 47 4e 4d 53 4d 4e 4e 56 51 50 4c 4c 51 45 4c 54 39 5c 5a 53 5d 4f 4c 4b 54 4e 52 50 52 4d 4f 53 52 4b 50 4c 4e 56 59 50 54 54 4e 4e 45 45 4e 4b 49 4a 46 46 43 47 4e 4b 44 40 42 3c 3e 2a 1a 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 0a 1b 16 25 2f 33 39 3f 33 3a 44 3c 3e 3d 3e 3f 42 3c 45 47 4a 46 41 41 43 4b 42 3f 47 45 4c 48 44 4b 4c 4b 50 4a 47 4f 49 52 50 4c 4e 53 4d 50 45 4e 4b 51 4f 47 4a 4b 46 4b 47 48 50 4c 47 42 48 49 4e 46 49 4d 47 45 4c 4e 4d 40 4a 42 47 44 3c 43 4d 48 4a 44 3d 3f 3d 3c 34 33 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 33 44 41 45 4b 4c 4c 50 44 42 49 4c 43 4c 4a 4f 51 4d 4f 4f 53 53 50 50 46 4a 4e 4e 4a 4d 4d 4d 50 41 4e 4d 51 47 4b 4e 46 4a 55 49 4a 52 4d 53 57 4a 50 55 51 46 4f 44 4e 52 4f 4c 54 51 4f 55 5a 4e 50 4f 4d 4d 54 49 54 49 4a 4a 45 49 48 4a 47 44 41 44 49 4c 43 41 41 43 48 44 2c 21 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 09 10 22 25 27 39 3f 43 3d 37 41 3b 38 3d 34 41 3f 4c 4a 45 44 49 43 48 45 40 43 48 44 43 52 47 4c 46 4f 4b 4a 44 4b 49 4c 51 53 4a 4b 4d 52 53 4e 49 4c 4c 44 4c 4e 52 46 48 49 48 4c 48 48 4d 49 47 4a 41 51 4e 46 45 47 4e 47 48 49 4b 4b 44 4a 3f 46 42 42 3c 45 41 40 3a 33 2e 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 29 3c 44 4d 4b 4d 51 51 4c 49 44 4e 45 55 4e 46 54 4d 50 52 4e 50 4b 51 50 4b 51 47 51 45 4f 42 47 48 4e 49 4f 52 4f 4f 4a 47 4c 4e 46 4c 46 53 4c 48 54 50 5b 53 49 53 4d 4c 55 4d 51 4d 4a 4a 4c 4f 46 48 4b 58 50 4d 4b 49 44 4a 47 43 47 44 4d 47 46 4c 3d 46 48 44 3f 43 40 35 31 1f 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0e 11 1a 23 28 35 35 3e 39 40 38 41 3e 3d 3f 42 49 45 4c 47 4d 51 46 4b 44
 42 45 45 42 42 4a 42 45 45 4b 47 4e 4c 45 45 47 4c 4b 48 4e 47 4e 51 4e 54 47 49 47 49 50 54 51 4a 4a 48 53 45 46 41 4b 46 44 48 4d 50 51 43 4b 4a 4a 42 4e 4f 45 4b 4c 46 43 50 40 46 46 44 3b 3c 3b 2c 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 25 49 47 4e 49 49 4d 4a 54 4c 48 4d 45 4b 50 4b 4d 51 50 4a 4e 4b 4b 4d 4e 4b 4b 47 4c 47 4b 4e 3e 4b 51 4e 4b 47 4a 4b 44 50 4c 46 44 46 4f 4b 53 4e 53 54 49 51 50 4b 4b 4d 50 4f 4d 55 48 4a 48 49 50 50 4e 4b 4b 4b 47 43 47 47 45 46 4f 4a 41 47 4f 4a 43 50 44 41 44 39 40 33 23 14 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 0f 11 18 21 33 39 3b 37 41 3d 3a 3e 3e 37 30 3b 40 3d 4d 43 44 45 41 40 46 41 49 3e 45 41 3b 48 4c 47 42 4c 3f 40 46 46 44 46 49 54 45 4c 51 44 49 45 47 42 46 40 45 4d 51 45 41 49 41 3e 47 45 46 3f 4e 46 47 4e 42 50 4b 4b 40 44 49 4b 47 48 4c 45 45 44 45 44 41 4a 3d 3c 2b 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 23 3f 41 3d 45 58 4f 4f 4a 45 4b 4d 4a 42 4e 4b 4a 4d 4c 4b 45 4f 4a 44 4b 4e 4b 4a 49 48 46 3f 45 41 42 47 40 4a 47 44 47 3f 41 4a 4b 4d 4b 49 4b 4c 46 4a 46 51 4b 4b 45 4a 47 41 48 4d 4f 55 53 4b 50 47 4e 55 51 42 47 45 41 3b 50 48 48 47 43 4a 46 41 44 40 41 48 42 3b 33 28 1f 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 12 17 1e 22 2b 2f 2f 3b 32 41 3d 3f 40 3c 40 3a 47 42 48 4f 3e 4e 4a 4b 48 49 45 43 4c 3f 44 3a 3b 53 4b 4b 48 45 47 47 47 44 4b 49 4f 3d 48 47 4a 42 4f 50 4d 42 48 45 47 43 48 4d 3b 44 40 3d 3e 47 43 4b 42 4b 44 4c 44 45 4f 47 45 4f 4d 49 46 40 4b 47 4a 44 3d 41 3b 36 37 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 28 3b 48 4d 4c 50 49 48 4c 45 4e 47 4f 46 4c 50 54 48 51 44 4a 50 47 4c 44 49 44 41 4f 4b 50 41 46 49 3e 45 4b 43 4b 3c 4a 43 42 4a 4a 52 40 4c 46 4a 4c 51 4a 48 52 4c 52 4d 4b 47 4f 4c 4e 4c 50 4d 48 44 4f 48 4e 4e 46 49 41 44 3d 47 44 4a 45 3e 42 49 49 4d 46 43 41 2e 30 22 12 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 0f 20 25 2b 35 30 38 2a 45 3e 37 37 39 3a 3b 42 40 3b 44 45 3e 45 48
 47 43 48 42 42 46 3e 46 3d 3c 44 45 3d 49 46 48 45 46 4d 4f 47 4c 4a 4a 42 4d 43 46 43 3d 49 45 48 47 4b 47 45 46 42 47 4e 4b 4c 45 49 4f 3e 49 4a 4a 45 4d 48 4c 4d 47 49 47 3c 46 42 43 44 48 42 39 38 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2b 44 4d 53 4a 47 4b 49 4d 47 50 41 4c 4c 49 4a 4b 48 4e 53 4b 52 46 4a 4e 45 4c 48 44 47 4a 3c 48 48 3f 46 43 44 44 44 49 46 44 44 43 47 46 4a 46 48 4e 44 46 4f 44 4c 54 4d 44 52 4f 4d 4a 4e 51 49 4d 4d 49 4a 4c 42 43 44 43 53 44 47 4f 41 4f 44 4c 44 45 4c 48 3b 44 36 23 23 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 16 12 1c 22 29 30 35 36 35 34 34 42 34 3c 40 38 44 3e 40 3c 41 48 44 41 43 3b 45 45 3b 3c 37 40 3b 3b 3a 3f 47 47 40 46 46 43 44 48 39 49 4b 50 4d 4a 4e 45 48 47 44 46 4e 4a 43 3e 45 44 48 49 3f 41 44 46 47 49 47 44 43 43 4b 4c 49 4c 45 41 4c 38 46 3f 41 40 41 3f 3b 3c 22 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 3e 43 4f 49 49 43 49 43 37 4f 49 42 3f 45 48 4c 42 3e 41 48 4b 49 42 4a 4b 4c 48 4d 3f 3d 43 3e 3f 39 42 4b 40 42 43 45 42 44 3d 46 4f 51 4d 46 47 45 4e 48 48 4b 4e 50 49 49 50 50 4f 5b 4b 50 4e 50 4f 47 47 49 3e 3d 41 46 3e 3e 43 4c 4e 48 43 44 40 3c 41 36 3e 36 24 21 09 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 06 0d 13 21 2e 2f 33 3a 3b 3a 38 32 3e 33 37 37 39 3d 43 3b 39 44 3e 41 44 3b 44 40 44 39 45 3d 46 44 48 3e 3f 44 43 42 44 4c 3b 41 42 35 45 44 45 44 44 45 4a 49 4d 45 4b 43 45 45 4d 44 46 4a 3f 45 4b 3e 44 49 42 46 3e 3d 44 44 48 42 45 47 48 4a 4c 3a 46 3a 41 40 38 32 25 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1b 46 4b 53 46 41 46 47 40 4b 49 45 3d 3c 3e 4b 45 47 42 49 41 42 45 43 43 42 4b 46 4c 47 3f 42 34 3b 3f 48 43 42 47 42 42 42 45 4f 4e 55 47 47 4a 40 42 44 52 44 46 52 4d 4e 4f 49 4a 4c 45 4d 4b 4c 4d 49 45 47 4c 44 37 42 4c 48 47 49 4c 43 49 4e 43 49 44 44 3b 39 36 23 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 07 0b 11 28 20 26 2b 32 32 37 34 3d 3b 36 48 45 36 3f 45 3e 3b 43 44
 3f 43 41 40 40 3d 44 44 40 44 3c 40 3e 47 45 42 4b 46 42 45 49 3e 3e 45 41 44 4e 46 44 47 44 41 45 45 49 4a 45 48 46 44 4c 48 45 46 39 4a 3b 43 4d 44 45 4b 4d 45 40 48 3f 49 41 40 3d 3e 45 41 4b 3e 3c 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 39 44 44 45 42 4b 43 48 4c 49 45 3d 48 48 4a 43 42 46 45 45 43 4d 3f 45 40 3b 37 3f 42 3d 43 3c 3d 4b 42 43 4d 40 4a 47 40 4b 43 46 50 4f 48 4f 49 4a 48 4f 4d 51 53 48 4a 44 49 52 50 4f 52 53 4b 4f 49 49 49 45 44 52 4e 4f 55 4c 4f 51 56 4d 4c 48 4a 46 3d 3c 31 28 1d 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 11 17 24 28 28 33 3d 3a 35 34 34 42 3d 41 42 3b 3f 3a 40 41 44 39 3f 43 3f 48 44 3e 3f 40 3f 3d 3e 3b 47 42 3d 44 42 45 43 3a 41 3d 41 3d 47 3e 43 48 4d 47 44 43 48 45 3f 43 45 4b 49 4d 43 45 42 3f 48 3b 3d 45 3f 3e 48 3b 43 4d 3f 45 45 43 45 3b 46 41 3e 41 3c 34 2c 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 30 3e 45 3b 46 3e 3c 44 40 41 49 47 48 44 42 2d 40 40 41 46 3e 45 40 3c 47 4a 3f 4d 40 41 3e 3e 47 44 48 46 46 44 3d 45 4b 4e 4e 44 47 48 50 4a 49 49 50 49 4e 4d 4d 48 47 4d 47 4c 4f 4c 41 51 44 52 54 4d 50 47 4e 50 55 5f 57 5a 5c 58 56 59 53 57 51 48 3e 2d 28 1b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 13 12 22 27 33 2c 38 3b 38 35 37 3a 35 39 36 3b 3f 3c 3b 3d 3c 3d 44 3e 3b 41 3e 3e 3c 48 3a 3f 47 40 3f 3d 41 44 40 45 44 3f 3a 45 43 42 38 3e 42 41 44 41 3f 42 40 3f 47 45 45 44 45 47 41 42 43 41 45 39 40 3b 39 3a 3a 3e 3f 41 40 47 3b 44 49 3e 41 45 38 38 36 39 29 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 27 3d 42 43 44 45 3f 45 44 49 41 45 36 3a 36 40 3c 3c 43 41 44 3f 3a 44 46 40 42 41 38 3d 42 3b 3e 48 43 3d 44 47 4a 45 49 4b 42 4d 51 4f 4b 47 4a 4c 4d 4e 4e 49 48 43 47 47 48 52 4e 50 57 4e 4a 4d 4a 50 57 51 59 54 4c 5d 68 62 60 67 62 65 5b 4c 47 3c 2f 33 22 0e 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 12 10 1c 29 25 28 30 37 36 34 35 3e 3e 3c 3c 38 3f 3c 3a 3b 43
 3b 3f 40 38 39 3e 3f 3b 41 44 4b 4b 3e 47 3e 3c 4b 41 47 44 3f 43 3e 3a 47 45 49 44 43 41 44 4a 4b 49 4e 45 4b 46 45 4b 41 42 47 41 48 41 3b 40 45 44 44 44 3f 3e 38 42 37 42 44 44 3c 43 45 42 39 3b 3f 28 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 2a 3b 47 44 47 3f 3a 40 39 3e 49 40 40 41 47 44 3e 3f 3e 43 3d 42 44 44 3f 3f 3a 48 41 39 37 39 45 3c 42 45 4a 49 44 46 52 45 4e 50 47 41 4d 4f 4b 50 4a 49 52 49 44 47 45 44 51 49 48 50 54 54 53 51 54 5c 64 58 5e 63 60 67 6d 70 65 69 68 62 57 4d 47 3f 3c 1f 17 12 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 1c 20 26 31 2e 3a 39 39 34 36 3b 3e 3a 41 41 37 44 3a 3b 38 3b 39 3e 3b 41 42 44 42 45 40 46 40 44 40 44 3b 3c 3d 43 3b 3a 4b 3d 47 44 40 3f 3e 49 44 45 49 3f 3f 4b 44 47 47 45 47 41 4b 43 43 41 44 47 42 47 43 3a 42 42 45 38 3e 3e 3d 44 3d 45 3c 3b 3d 3b 39 28 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 28 41 4b 41 44 3a 3e 41 37 3b 3a 3d 42 45 3b 41 41 3b 3d 44 31 3c 40 3f 43 37 40 44 41 43 43 3b 48 41 45 46 46 46 47 51 49 39 50 4b 52 4b 44 4b 51 44 56 48 4f 50 43 4b 48 4c 44 4e 59 4b 57 57 50 55 5a 5a 65 69 77 6e 71 73 6d 6e 6f 6a 68 61 56 5c 41 39 2c 15 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 15 15 21 2f 26 2b 31 37 32 39 3d 35 37 38 39 40 3d 3f 3c 3d 3d 3a 36 3d 3d 36 35 42 3c 48 43 3e 3c 41 49 41 3d 37 40 43 45 44 40 3d 3b 3b 45 47 40 43 42 44 44 48 4b 48 45 4d 4d 45 4a 48 44 48 3f 3c 3c 46 3e 3a 38 33 38 3d 40 3f 37 3a 39 39 40 3b 43 3c 34 30 2b 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 25 3a 47 41 3c 3d 3e 42 3c 44 3b 37 40 3e 35 40 3e 42 3e 42 40 3e 40 3f 38 3a 3d 42 46 43 38 45 3b 46 43 3f 4c 42 48 3d 44 43 46 45 4a 4e 52 4f 40 49 48 43 49 46 49 45 44 4d 4d 52 53 53 4f 55 56 62 6f 76 73 72 68 80 6e 6c 77 61 6e 65 66 64 57 53 39 31 22 14 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 14 22 21 31 2f 2d 33 31 37 3c 37 43 43 3d 3b 3b 35 35
 3a 41 3d 3e 39 42 39 40 3a 3f 41 41 3e 3e 3a 43 3f 42 41 41 42 45 3d 44 3f 40 48 46 41 47 44 46 45 42 4c 56 4f 54 56 4e 55 42 4b 44 3d 3d 39 41 47 42 40 3b 39 3c 3a 40 3c 37 3b 3c 36 46 38 3a 33 2d 35 2c 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 26 43 44 3d 46 3d 3c 47 37 3a 41 42 3c 3d 3e 3d 41 3a 37 3f 3d 47 3e 41 3f 3a 44 40 41 45 3e 44 44 4a 46 48 4a 47 43 43 43 45 47 44 4f 4c 50 4d 4d 4e 4a 4e 45 43 49 4b 44 4a 51 4d 52 5a 57 64 66 68 6f 76 7e 7a 75 73 6c 71 6b 6a 6b 62 5f 50 2a 36 32 2d 19 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 18 1d 2f 26 2c 35 34 32 38 37 3d 3f 2e 3c 3a 32 42 3a 3d 3d 45 3d 36 3f 3f 3d 3a 45 3b 3a 3d 36 45 3e 3a 43 3a 42 3e 47 44 41 3c 45 4a 4d 47 4c 44 43 49 4a 49 57 5e 5d 5c 5b 50 4a 47 3a 3d 41 3d 3d 3c 3a 3f 3e 37 3d 37 38 3f 43 34 35 3b 3e 31 34 38 35 30 25 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2f 3c 3f 41 44 3f 44 43 37 37 42 3e 40 47 3d 42 35 3c 3b 40 43 42 44 36 3c 3d 3e 3f 3b 44 45 43 45 3d 44 41 45 3e 43 44 49 4b 4b 43 49 49 45 4e 45 44 4c 4b 46 49 48 45 46 54 49 5f 57 66 62 72 71 7d 81 80 8b 75 70 79 6f 6d 69 66 5d 63 59 54 45 36 22 1f 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0d 11 1c 25 26 25 2a 36 35 32 3a 37 3c 43 3d 3a 3f 3f 43 41 44 3e 41 41 40 39 3d 36 36 3c 38 3f 43 36 3c 38 47 43 44 3d 35 43 45 4c 47 44 51 48 47 41 45 49 4e 50 60 5f 5b 5a 53 50 45 48 42 35 3a 39 3e 35 36 36 33 36 3a 37 2d 35 3b 3e 31 3c 3e 33 33 34 32 2f 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 1a 37 4a 46 42 3a 3e 3f 3b 45 3f 3f 33 3e 41 3e 3e 3b 3f 3c 37 42 3e 41 3f 3f 43 47 40 44 42 44 3d 46 41 42 42 41 46 44 48 3e 3a 40 43 47 4d 4e 4a 4f 42 48 52 4d 4b 44 44 4d 50 5c 63 6f 7f 7d 79 7f 7e 84 7f 7d 77 75 69 67 66 63 65 56 58 4a 38 30 16 0b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 11 1a 25 29 2e 32 27 2c 3a 34 41 39 37 38 38 40 3f
 44 46 38 41 42 43 39 37 3d 42 3f 3b 3b 3e 3b 3b 39 3d 45 41 3e 3e 3e 42 49 44 49 49 43 4e 45 45 49 43 4d 54 5d 5e 5d 63 49 47 43 40 37 34 32 35 3d 3a 40 35 3b 3a 37 3d 36 33 3e 37 38 3b 37 3a 35 38 33 28 15 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 3b 40 40 41 3e 35 47 40 46 42 42 42 3e 49 41 46 41 41 44 46 46 44 3d 44 45 3b 48 45 45 43 45 41 44 42 45 46 3c 40 37 39 3f 3f 45 45 42 49 41 49 40 42 47 4f 4a 4e 56 4d 60 5d 6a 72 77 7f 82 81 7f 7c 78 75 79 7a 6d 66 6c 62 64 62 51 52 43 30 21 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 14 1f 22 21 24 30 30 39 38 39 3a 40 38 3b 3c 37 3a 39 3b 43 45 3e 3e 40 35 3b 39 3a 35 38 35 38 32 3f 37 3c 39 3d 41 43 43 3f 4a 46 4f 4a 46 44 42 43 4c 55 4a 59 58 51 47 48 42 40 37 44 35 3b 36 35 3e 3d 33 3d 33 37 3b 35 3a 3a 3b 35 32 40 30 38 35 35 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1c 3f 42 48 43 3d 3b 41 3e 3d 43 3d 41 48 42 46 44 49 48 49 49 4b 48 4b 49 43 40 41 43 4b 45 42 3c 3e 3e 4b 3e 3a 38 3d 41 3f 45 42 3f 46 41 44 43 45 49 4b 48 4e 4b 4a 4b 5e 6c 80 7e 7d 85 7f 7d 81 7b 7a 75 70 66 6d 61 69 5d 5e 52 53 4e 34 22 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0e 1b 25 26 28 28 30 2f 31 34 39 3d 39 3d 42 37 42 41 3f 41 44 3f 3b 3a 3a 3e 30 37 38 35 3e 33 30 39 3b 3e 3a 44 3e 37 47 42 46 44 44 44 39 42 3d 47 3e 4a 51 46 47 4d 43 3f 3e 3c 3e 3d 3a 3c 39 35 38 35 39 32 36 35 35 31 3d 3c 38 3b 36 36 37 33 38 30 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 3a 3f 48 40 3e 41 46 3f 44 3f 42 4a 4c 47 46 43 47 44 43 49 46 47 4b 45 4a 43 43 45 42 43 3a 3e 3d 35 41 3d 36 37 36 3c 3a 3b 42 44 41 44 45 40 3f 48 46 4c 3f 4d 53 5f 68 75 77 81 7d 83 80 7b 74 7a 74 6e 6c 61 65 5e 62 67 55 52 46 3b 2c 1a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 11 19 1b 2a 2a 31 2e 32 3b 3c 3f 4a 44 3d 3b
 43 3c 45 49 37 48 3e 43 40 47 39 3b 3a 3a 36 3d 37 34 38 3d 36 39 35 3b 3e 42 3e 3c 3a 3f 3c 40 36 38 40 47 3f 44 47 45 48 3a 3e 3b 37 40 39 3c 41 35 3d 36 31 33 36 3a 36 30 3d 42 45 38 37 36 35 39 33 2f 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 32 3c 4a 48 41 42 47 3a 40 45 44 3d 46 40 44 42 49 49 4c 42 4d 45 44 4c 4b 3c 44 3a 45 3e 3e 3c 38 3b 41 3d 3d 3d 39 3b 44 3d 3d 47 45 43 43 43 48 45 42 4d 4c 59 63 6e 78 7b 88 89 83 80 75 76 7c 78 6a 70 6d 64 69 5b 58 59 53 49 40 32 1d 07 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0d 1e 25 2a 30 2c 34 36 3b 44 3e 42 38 3b 3a 44 43 40 42 45 44 43 41 43 3c 39 3d 3d 34 44 36 37 39 37 35 38 3c 3c 44 3a 3e 36 39 3c 37 3f 40 40 3e 3b 3e 3f 41 39 3d 39 3a 3e 3f 41 38 35 3c 3a 31 37 3c 32 37 32 39 37 36 3f 3d 41 38 35 38 34 30 30 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 35 3c 46 43 44 3a 48 3e 3b 39 40 40 39 4c 44 38 40 4a 42 46 48 47 4e 4d 43 41 44 40 3d 41 37 3b 44 35 37 39 3f 34 3e 3f 3d 43 4c 48 45 3c 46 47 46 4b 4b 58 5f 67 77 7d 7d 7f 83 86 81 81 76 7b 78 6d 6d 6c 6c 6a 5e 51 5c 51 43 41 34 22 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 19 14 26 2d 2c 2f 32 37 39 3d 3b 35 37 3d 4a 3a 44 3d 4a 4b 42 44 44 3c 3b 37 3f 32 35 2d 37 33 38 3a 34 3a 3c 3a 40 33 3a 38 31 36 39 39 39 36 3a 3e 3d 35 3f 39 31 31 3f 39 3c 3d 3e 36 31 2e 33 35 3e 32 2f 3b 2f 30 30 38 3a 37 35 33 30 2c 30 1e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 36 35 33 3f 46 42 4b 3e 41 3d 3b 3d 41 41 41 3c 38 40 44 43 45 3c 46 44 43 3d 3f 41 41 37 35 33 3d 3b 3e 39 3d 35 42 3a 39 3e 40 43 40 48 4a 4d 4c 52 55 63 6c 74 84 81 7f 7e 7d 7b 71 77 7b 6e 6c 6e 64 68 71 65 5e 54 52 4d 42 33 23 11 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 19 20 24 2c 30 3a 38 3c 3c 36 43 3d
 3b 3f 40 44 41 46 43 49 44 45 3a 35 36 3b 3b 3b 35 36 41 35 3c 3a 35 37 3e 38 30 32 2e 37 3d 3b 37 34 36 39 3d 40 35 33 37 38 39 42 3c 3b 2b 35 39 36 3b 3e 31 39 31 33 35 36 2e 2e 31 33 36 35 33 31 2f 36 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 2e 3f 35 39 3f 3e 4e 4a 47 4a 42 3f 35 3c 35 40 42 41 3c 43 3b 37 3c 48 47 3d 3c 34 41 3a 37 38 3f 3e 40 3f 40 46 42 38 39 42 45 40 40 55 48 47 55 62 6d 72 79 83 88 80 7f 7f 78 7d 72 79 68 6a 69 5d 5e 5b 5f 62 57 4b 4d 42 3a 2a 12 08 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 12 18 29 1f 30 2b 2d 3d 38 38 40 3a 40 47 45 43 44 46 3d 4b 47 4c 40 34 37 38 31 33 3b 33 32 3a 34 38 33 3c 39 33 35 33 3a 3a 37 36 32 3d 39 3d 35 3e 39 39 42 3a 3f 3b 39 42 3f 36 3d 33 33 36 33 32 38 34 31 37 3a 3b 37 38 37 2a 33 2f 2f 2c 22 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 26 38 38 3e 3f 3e 4a 48 45 4a 46 37 45 39 40 40 3c 3f 42 3c 3f 40 3e 3c 3b 42 42 36 34 37 3e 3b 3b 41 3c 35 39 37 31 46 43 42 45 45 46 55 53 5e 69 72 7a 7c 86 82 80 82 79 80 74 79 72 71 4f 64 63 62 62 66 58 5a 58 4c 3f 34 2d 1b 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 1c 1b 24 25 2d 2f 2f 34 2f 35 31 46 45 43 4b 47 47 47 3b 3e 43 3b 42 38 3b 34 3e 33 41 36 35 31 30 35 32 35 40 37 3a 32 31 32 37 32 37 37 30 25 3a 32 39 34 32 3a 3f 3e 36 3c 33 36 33 34 3b 33 34 39 2b 33 2d 2b 33 36 31 26 2b 33 30 39 2c 25 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 2b 2b 39 36 3a 36 49 3c 53 4b 38 39 38 39 45 48 40 3d 3f 3d 3d 3b 40 44 3a 3a 41 36 3b 42 38 41 3f 39 3b 3a 35 43 37 3d 3c 42 41 48 49 56 6a 72 78 80 7f 7c 81 76 78 78 71 70 75 65 6a 6e 64 6a 65 5a 59 5b 55 4d 50 3a 31 22 16 0a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0e 17 28 23 23 25 34 2e 35 35 3c
 3b 47 4c 48 45 41 3f 3f 3f 3b 40 39 3c 37 38 32 2e 38 35 3a 3e 3c 39 34 30 30 36 39 35 38 32 36 33 37 3a 3c 32 2b 2e 35 35 3f 35 31 35 30 39 38 34 2e 37 32 36 37 35 2a 30 35 37 3e 31 2e 34 2f 2f 30 2f 2a 1b 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 23 34 39 3a 39 35 3f 47 40 35 3c 32 32 3c 34 37 41 36 36 3e 35 41 43 3b 3b 35 3c 32 3e 37 37 38 3c 3a 38 42 38 40 45 44 48 40 53 5e 64 71 73 78 7d 80 81 7a 81 79 78 6e 6f 72 6a 68 5e 6b 5b 5f 60 56 51 56 4f 47 3a 33 28 1b 16 05 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0f 20 20 2d 24 2e 2d 30 35 30 40 39 46 44 45 48 41 3f 47 40 39 38 3b 37 3c 3f 33 33 37 40 37 3c 39 39 3a 3b 3c 35 2f 32 32 40 37 35 37 37 35 30 36 33 34 2c 38 38 36 3a 38 32 32 2f 34 33 33 35 30 25 31 31 39 37 2d 33 2c 32 2f 31 2c 2a 27 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 30 35 3b 43 40 3f 41 42 39 35 37 38 39 39 38 33 3d 3a 3d 2a 3b 39 3a 3c 3e 37 44 3a 2a 3f 38 43 38 3b 3d 3e 41 44 48 51 4d 5c 6d 6a 85 7e 7a 7f 7e 7e 7c 76 79 75 76 6f 64 6e 62 63 61 5d 5a 62 5c 53 53 4a 42 39 2b 20 16 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 17 1a 23 22 24 2c 2e 2f 32 3a 42 48 44 43 4c 3f 44 3b 38 3d 39 3b 3a 3e 3f 37 3c 3c 3f 35 3b 2f 37 3c 34 3a 33 33 2f 35 36 38 39 3c 36 2b 31 30 35 3a 32 31 39 33 2f 31 31 35 38 31 31 33 30 37 32 30 2e 35 32 2a 38 2e 2d 33 2c 27 2c 19 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1c 2c 30 3b 38 3d 44 38 39 36 2d 34 39 33 35 33 33 30 36 37 36 36 38 30 36 3e 37 38 35 37 39 37 3c 3c 40 3e 3d 41 44 4c 57 61 6c 75 75 7f 7e 7a 7b 7c 75 6c 70 6c 66 66 63 5f 64 61 5d 56 60 4c 4b 4f 47 54 3e 3b 2e 1f 14 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 1f 20 26 22 22 2a 2e
 37 39 37 43 3d 3b 39 3b 43 44 3b 3b 3a 36 33 3c 37 42 37 3b 3a 3e 3e 32 39 32 31 37 38 2c 2d 40 36 36 35 3b 37 34 2b 30 34 30 2f 34 34 3a 2a 33 2a 2e 2b 26 2e 30 2f 2e 33 30 2b 31 31 34 2b 34 28 28 2a 29 27 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 2a 33 32 3c 3d 3b 2e 36 31 24 33 34 2b 38 30 29 2b 2e 32 2d 35 3f 27 33 37 37 2c 34 2c 2c 34 30 3b 3d 36 3e 4a 57 60 60 75 76 79 71 74 7c 70 73 72 6d 68 65 5f 5d 61 5d 58 5e 5e 4e 4f 4a 53 54 4d 44 3a 31 23 1f 06 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 11 14 1d 26 28 2e 2d 31 2e 33 3a 3d 3c 45 3c 3b 41 3e 41 3b 36 42 39 34 3b 3b 37 3d 31 3a 3e 3b 38 39 36 3b 40 3c 3e 30 32 31 3c 38 30 2d 35 39 33 31 36 2f 28 31 2f 36 30 2c 29 2a 2e 2f 2e 2a 34 27 34 30 27 2f 2c 32 28 2c 29 2c 27 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 21 2e 33 35 41 39 33 31 32 2e 2a 33 35 37 2a 31 25 2b 2e 31 35 30 2f 31 2f 2e 33 32 31 33 34 39 3e 3e 44 50 52 57 73 69 72 68 71 70 6c 63 65 6c 6a 66 5f 5f 5b 5e 53 58 56 55 4a 4b 4b 4f 45 4e 46 32 33 25 15 0c 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 10 1a 1f 23 1f 25 29 2e 33 2f 38 3d 3d 31 34 3c 47 3a 39 3d 3f 3d 3b 38 39 3e 3e 34 3c 38 38 3b 37 31 3c 38 31 3c 40 43 35 35 35 34 35 33 2e 2e 2a 2f 2f 2e 2a 21 25 2e 2b 23 2c 28 2f 2b 2f 31 32 24 30 2a 2d 2d 26 27 24 2c 27 1b 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 17 25 30 2a 26 2a 2a 28 23 1e 24 22 2f 24 22 26 2b 23 1f 24 29 2b 28 2e 25 2e 2c 2d 2b 28 2b 34 47 43 4c 51 5a 60 62 5b 60 5a 5c 5a 59 56 51 50 50 4e 4c 4e 54 47 46 50 4f 47 4a 49 45 4b 39 31 2f 28 22 17 0e 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0e 17 19 24 23 24
 32 31 2a 2c 2f 35 39 34 34 38 35 37 33 36 39 37 33 35 38 3b 38 38 36 2c 35 3a 36 34 3c 31 3b 44 4a 39 37 3b 28 2b 2b 2a 30 2a 29 2a 20 1e 12 1f 1c 1e 21 24 26 2b 2d 28 2a 21 26 2a 1c 25 27 28 22 1e 1e 22 17 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 25 1d 1e 1a 16 22 1d 1d 19 1a 1d 15 15 17 15 14 11 24 1e 18 22 1e 1e 14 24 22 1f 20 1c 2f 30 36 40 3f 44 3f 42 3e 40 42 44 41 45 40 48 3a 3b 3c 3a 3e 39 36 3b 34 33 33 3f 35 37 35 2e 29 29 21 14 09 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 16 0e 23 25 25 26 2a 29 2e 39 38 30 35 33 37 3a 36 2c 34 39 3d 37 31 3d 37 39 34 3a 35 37 3d 35 35 38 35 3d 4d 49 41 49 39 3e 32 29 2d 2f 28 26 25 15 11 09 14 18 18 1b 23 28 20 26 29 1f 27 22 24 1f 21 25 21 18 18 16 12 14 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 11 0e 0c 0b 0d 15 10 0e 0a 0f 17 0d 16 11 14 0e 11 0f 0a 15 10 14 15 0b 12 1d 18 21 25 2d 2d 31 32 31 30 28 2c 2f 2a 2f 2c 2f 2a 32 29 22 31 27 2c 27 27 30 26 23 1f 24 27 1f 17 19 0d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 17 16 1b 2b 2c 26 26 2b 31 2b 2d 33 36 34 35 38 34 36 35 30 32 3a 39 32 32 38 34 42 3e 35 35 38 3b 41 42 47 41 47 42 3a 32 33 2d 28 27 22 1c 17 08 06 05 0e 0b 15 0d 19 1d 1f 20 16 16 1a 14 0b 14 0d 0b 14 0f 0e 0b 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 0f 0c 05 03 05 06 05 03 00 0d 08 03 04 0b 08 0d 0d 08 18 12 12 0c 15 15 15 16 1e 1d 19 1b 1e 15 15 18 1c 1f 21 14 18 1e 13 10 1b 17 1b 15 1b 1d 1a 14 12 19 0b 10 08 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 17 13 23
 20 24 21 27 25 1f 28 2e 30 2e 28 31 31 30 2c 33 36 30 38 34 30 38 2f 34 32 2f 2d 2f 39 2b 42 3b 3a 36 3c 41 30 2a 21 21 22 1f 12 0b 05 00 06 05 03 00 09 08 0a 0b 06 0d 0b 04 06 0b 06 0d 06 05 07 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 0d 09 01 06 06 03 07 08 06 0c 04 07 05 0e 04 06 05 03 0c 07 0a 0b 09 06 08 03 06 06 0b 05 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 1e 1b 26 23 20 24 23 2d 2d 2f 2f 2e 32 2c 2f 33 2b 28 27 29 2a 2a 2f 27 25 2c 23 18 1b 26 2b 2b 2f 32 3a 33 32 26 2a 21 21 17 14 11 08 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 1d 1d 1d 1c 23 1b 20 28 2a 25 26 1e 2e 22 27 21 21 20 25 2b 26 22 26 23 1b 16 15 0e 09 12 15 1c 19 1f 1f 20 17 0f 16 0a 0b 0d 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 08 07 0e 15 15 1b 1b 1f 18 23 14 21 1e 1f 1a 1d 13 12 19 11 13 19 21 10 14 0a 09 06 03 01 06 0d 06 00 0d 06 0f 05 06 09 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 09 1b 14 0b 17 11 16 16 0c 10 0a 08 08 06 06 09 04 06 0c 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 03 0f 06 05 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
