 ff ff 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 49 52 52 52 5b 5b 52 52 49 52 00 49 49 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 9b a4 f7 07 f7 07 07 07 f7 a4 a4 f7 f7 f7 a4 5b 52 49 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 52 5b a4 a4 a4 a4 f7 07 f6 ff ff f6 07 f7 f7 a4 9b a4 a4 9b 9b 5b 5b 5b 5b 52 49 49 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 52 a4 a4 9b 9b a4 f7 f7 07 07 ff ff ff ff ff ff ff 08 07 f7 f7 a4 a4 f7 a4 a4 a4 5b 5b 5b 5b 5b 52 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 52 5b 9b 9b a4 a4 f7 07 07 08 f6 ff ff ff ff ff ff ff ff ff f6 07 07 f7 07 07 f7 f7 a4 a4 a4 9b 9b 5b 52 9b 52 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 49 9b 5b 9b a4 f7 f7 07 07 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 08 07 08 07 f7 f7 f7 a4 9b 9b 9b 9b 5b 5b 52 49 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 52 a4 5b a4 a4 f7 07 07 08 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 08 07 07 f7 f7 a4 a4 a4 a4 5b 9b 9b 9b 49 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 49 52 a4 5b a4 f7 07 07 08 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 f6 f6 f6 f6 07 07 07 07 f7 f7 a4 9b a4 9b a4 52 00 00 00 00 00
 00 00 00 00 00 00 00 00 49 52 f7 a4 9b a4 f7 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ff f6 f6 f6 08 f6 f6 f6 f6 f6 f6 f6 ff f6 08 08 07 07 f7 a4 a4 a4 a4 a4 9b 00 00 00 00 00
 00 00 00 00 00 00 00 52 a4 a4 a4 a4 a4 f7 07 08 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 08 f6 f6 f6 f6 f6 f6 f6 f6 f6 08 07 07 f7 a4 a4 a4 a4 a4 f7 49 00 00 00 00
 00 00 00 00 00 00 52 a4 f7 a4 a4 f7 f7 07 07 08 08 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 08 f6 f6 f6 f6 f6 f6 f6 08 07 f7 f7 a4 a4 a4 a4 9b 9b f7 49 00 00 00 00
 00 00 00 00 00 00 52 07 a4 a4 a4 a4 f7 07 07 08 08 f6 f6 ff ff ff ff f6 ff f6 ff ff ff ff ff ff ff ff ff ff f6 f6 f6 f6 f6 f6 f6 f6 08 07 07 f7 a4 a4 a4 a4 9b 9b f7 49 00 00 00 00
 00 00 00 00 00 00 9b f7 a4 a4 a4 a4 f7 07 07 08 f6 f6 f6 ff ff f6 f6 f6 f6 ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 f6 f6 f6 f6 f6 08 07 07 f7 a4 f7 a4 a4 a4 9b a4 49 00 00 00 00
 00 00 00 00 00 49 a4 5b 9b a4 a4 f7 f7 07 07 07 08 f6 f6 f6 f6 f6 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff 08 08 f6 f6 f6 08 08 08 07 07 07 f7 f7 f7 f7 a4 a4 a4 a4 52 00 00 00 00
 00 00 00 00 00 49 f7 5b 9b a4 f7 f7 f7 07 07 08 f6 f6 f6 f6 f6 f6 f6 f6 ff ff ff ff ff ff 07 07 ff 07 ff ff 08 08 08 f6 08 08 08 07 07 07 f7 f7 f7 a4 f7 a4 a4 5b f7 5b 00 00 00 00
 00 00 00 00 00 49 f7 9b 9b a4 a4 f7 07 07 08 f6 f6 f6 ff f6 f6 ff ff ff ff ff ff ff ff 9b 5b 52 52 5b f7 f6 07 08 07 07 07 07 07 07 f7 f7 f7 f7 f7 a4 a4 a4 9b 5b f7 5b 00 00 00 00
 00 00 00 00 00 49 f7 9b 9b 9b a4 f7 07 07 08 08 f6 f6 f6 f6 f6 f6 ff ff ff f6 f6 ff f7 52 49 49 49 52 52 08 07 07 07 07 07 f7 f7 f7 f7 f7 a4 a4 a4 a4 a4 a4 9b 5b f7 5b 00 00 00 00
 00 00 00 00 00 49 a4 a4 a4 a4 a4 f7 07 07 07 07 07 08 08 f6 f6 f6 f6 f6 f6 f6 f6 08 5b 49 00 00 00 49 49 07 07 07 07 07 f7 f7 f7 f7 f7 a4 a4 a4 a4 a4 a4 a4 9b 5b f7 9b 00 00 00 00
 00 00 00 00 00 49 a4 a4 a4 a4 f7 f7 f7 07 07 07 07 07 07 07 07 08 08 08 08 08 08 07 52 00 00 00 00 00 00 07 07 07 07 f7 a4 a4 a4 a4 a4 a4 a4 f7 a4 a4 a4 a4 9b 5b a4 5b 00 00 00 00
 00 00 00 00 00 49 a4 a4 a4 a4 f7 f7 f7 f7 f7 f7 f7 f7 07 07 07 07 07 07 07 07 07 f7 5b 00 00 00 00 00 00 f7 f7 f7 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 9b 9b 5b a4 5b 00 00 00 00
 00 00 00 00 00 49 a4 9b a4 a4 f7 f7 f7 f7 f7 07 07 f7 f7 f7 f7 f7 f7 f7 f7 f7 f7 a4 9b 00 00 00 00 00 00 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 9b 9b a4 a4 a4 9b 9b 5b 00 00 00 00
 00 00 00 00 00 49 a4 9b 9b 9b a4 a4 f7 f7 f7 f7 f7 f7 f7 f7 f7 a4 f7 a4 a4 a4 a4 a4 9b 00 00 00 00 00 00 a4 a4 a4 9b 9b a4 9b a4 a4 a4 a4 9b 9b 9b 9b 9b a4 9b 9b 9b 9b 00 00 00 00
 00 00 00 00 00 49 a4 9b 9b 9b a4 a4 a4 f7 f7 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 5b 00 00 00 00 00 00 9b 9b 9b 9b 5b 9b a4 a4 a4 a4 9b 9b 9b 9b 5b 9b 9b 9b 9b 5b 9b 00 00 00 00
 00 00 00 00 00 49 9b 9b 9b 9b a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 a4 9b a4 9b a4 9b 9b 5b 00 00 00 00 00 00 5b 5b 5b 5b 5b 9b 9b 9b 9b 5b 9b 9b 9b 5b 5b 9b 9b 5b 9b 5b a4 00 00 00 00
 00 00 00 00 00 52 9b 9b 9b 9b a4 a4 a4 a4 a4 a4 a4 a4 a4 9b 9b 9b 9b 9b a4 9b 5b 5b 5b 00 00 00 00 00 00 5b 5b 9b 5b 5b 9b 9b 5b 5b 5b 9b 5b 5b 5b 5b 9b 5b 9b 5b 5b 5b 00 00 00 00
 00 00 00 00 00 52 5b 5b 9b 5b 5b 9b 9b 9b a4 a4 a4 9b 9b 9b 5b 5b 9b 9b 9b 9b 5b 5b 52 00 00 00 00 00 00 52 5b 5b 5b 5b 9b 5b 5b 5b 5b 5b 5b 5b 5b 9b 5b 5b 5b 5b 5b 52 00 00 00 00
 00 00 00 00 00 52 5b 9b 9b 9b 9b 9b 9b 9b 9b a4 9b 9b 9b 5b 9b 9b 9b 9b 5b 52 5b 52 52 00 00 00 00 00 00 52 5b 5b 5b 5b 5b 5b 5b 5b 5b 5b 52 5b 5b 5b 5b 5b 5b 5b 5b 52 00 00 00 00
 00 00 00 00 00 52 9b 5b 5b 5b 5b 9b 9b 9b 5b 9b 9b 9b 9b 5b 5b 5b a4 5b 5b 5b 52 5b 52 00 00 00 00 00 00 52 52 5b 9b 5b 5b 5b 5b 5b 52 5b 52 52 5b 5b 5b 52 5b 5b 5b 49 00 00 00 00
 00 00 00 00 00 52 a4 5b 9b 5b 9b 5b 5b 5b 5b 5b 5b 5b 9b 9b 5b a4 9b 9b 5b 5b 52 52 52 00 00 00 00 00 00 52 52 52 5b 5b 5b 5b 5b 5b 5b 5b 52 5b 52 5b 52 5b 5b 5b 5b 49 00 00 00 00
 00 00 00 00 00 49 9b 5b 5b 5b 5b 5b 9b 9b 5b 5b 5b 5b 9b 5b 5b 9b 9b 52 5b 5b 52 52 52 00 00 00 00 00 00 49 52 5b 52 5b 5b 5b 5b 5b 52 5b 52 52 52 5b 52 5b 5b 5b 5b 00 00 00 00 00
 00 00 00 00 00 00 52 5b 5b 5b 5b 5b 52 5b 5b 5b 5b 5b 5b 52 5b 9b 9b 5b 5b 5b 52 5b 52 00 00 00 00 00 00 00 5b 52 52 5b 5b 5b 5b 52 5b 5b 5b 52 52 5b 52 5b 5b 52 52 00 00 00 00 00
 00 00 00 00 00 00 52 9b 5b 52 5b 5b 5b 5b 52 5b 5b 52 52 5b 5b 5b 52 52 5b 5b 9b 5b 52 00 00 00 00 00 00 00 52 5b 5b 9b 5b 5b 52 52 5b 5b 52 52 52 5b 5b 5b 5b 5b 49 00 00 00 00 00
 00 00 00 00 00 00 49 52 5b 5b 5b 52 52 52 52 52 5b 5b 5b 52 52 5b 52 52 52 5b 5b 5b 9b 00 00 00 00 00 00 00 5b 5b 5b 5b 5b 5b 52 5b 5b 5b 5b 52 52 52 52 5b 5b 52 00 00 00 00 00 00
 00 00 00 00 00 00 00 52 52 52 52 5b 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 5b 5b 00 00 00 00 00 00 00 5b 5b 5b 5b 5b 5b 5b 52 9b 5b 52 5b 52 52 5b 5b 5b 49 00 00 00 00 00 00
 00 00 00 00 00 00 00 49 5b 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 5b 00 00 00 00 00 00 00 5b 52 5b 5b 5b 5b 5b 5b 5b 5b 52 52 52 52 5b 5b 52 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 5b 5b 52 52 00 00 00 00 00 00 00 52 52 5b 5b 5b 5b 5b 52 52 52 52 5b 5b 52 5b 5b 52 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 5b 5b 52 52 52 52 52 52 52 5b 5b 52 49 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 5b 5b 5b 5b 52 52 52 52 52 52 52 52 52 5b 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 5b 52 49 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 5b 52 52 00 00 00 00 00 00 00 52 5b 52 52 52 52 52 52 52 52 52 5b 5b 9b 52 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 52 5b a4 f7 a4 a4 52 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 52 52 5b 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 52 52 52 52 a4 f7 f7 a4 a4 a4 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 5b 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 52 52 52 f7 f7 a4 a4 a4 9b 5b 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 52 52 52 52 52 5b f7 a4 a4 a4 a4 9b 9b 49 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 52 49 52 52 52 00 00 00 00 00 00 00 49 52 52 52 9b a4 a4 a4 9b 9b 9b 9b 5b 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 49 52 52 49 00 00 00 00 00 00 00 52 52 5b a4 a4 a4 a4 9b 9b 9b 5b 5b 49 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 52 52 49 00 00 00 00 00 00 00 52 5b a4 a4 a4 a4 9b 9b 9b 5b 52 52 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 52 52 52 52 52 52 52 52 00 00 00 00 00 00 00 5b a4 a4 a4 a4 9b 5b 9b 5b 5b 52 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 52 52 52 49 52 52 52 5b 52 52 00 00 00 00 00 00 00 52 9b 5b 5b 9b 52 52 52 52 49 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 49 49 49 49 49 52 5b 52 52 00 00 00 00 00 00 00 00 00 49 00 49 49 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
