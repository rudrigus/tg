-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "11/18/2015 21:55:21"
                                                            
-- Vhdl Test Bench template for design  :  ProcessadorImagemGMAW
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;
--use work.imagensteste.all;

ENTITY ProcessadorImagemGMAW_TB IS
END ProcessadorImagemGMAW_TB;
ARCHITECTURE ProcessadorImagemGMAW_arch OF ProcessadorImagemGMAW_TB IS
-- constants                                                 
  -- usando Img332 a Img335 de "Resultados 2 Livre com valores de trigger muito baixos 70 150"
  constant imagem_teste0 : MatrizImagem :=  ((X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"13", X"20", X"22", X"1a", X"13", X"0b", X"0f", X"10", X"13", X"06", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"1b", X"30", X"41", X"3a", X"38", X"34", X"31", X"3b", X"3d", X"3b", X"24", X"1b", X"19", X"15", X"0f", X"04", X"03", X"03", X"02", X"03", X"03", X"05", X"09", X"0b", X"0a", X"0b", X"0c", X"0e", X"1a", X"22", X"25", X"21", X"22", X"22", X"16", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"17", X"2e", X"4b", X"4d", X"3e", X"3b", X"38", X"3b", X"4f", X"56", X"55", X"4f", X"30", X"2d", X"29", X"24", X"05", X"03", X"03", X"02", X"03", X"03", X"0e", X"2a", X"27", X"27", X"28", X"2a", X"2a", X"2f", X"42", X"5d", X"67", X"62", X"5f", X"5a", X"34", X"07", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0e", X"28", X"3a", X"48", X"3f", X"3c", X"38", X"39", X"3c", X"4f", X"5b", X"5a", X"5c", X"3b", X"31", X"2c", X"26", X"05", X"03", X"03", X"02", X"03", X"03", X"14", X"31", X"2f", X"2f", X"2e", X"2f", X"32", X"34", X"36", X"3e", X"5a", X"71", X"75", X"72", X"65", X"2c", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"1f", X"31", X"3e", X"3d", X"3c", X"3b", X"38", X"3f", X"3f", X"4a", X"52", X"51", X"55", X"3b", X"32", X"2f", X"26", X"04", X"03", X"03", X"02", X"03", X"03", X"18", X"31", X"32", X"32", X"32", X"31", X"31", X"34", X"36", X"37", X"3a", X"45", X"60", X"70", X"6c", X"46", X"19", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"13", X"2a", X"3a", X"3e", X"3e", X"3c", X"3b", X"3b", X"3d", X"3e", X"48", X"49", X"42", X"44", X"37", X"31", X"31", X"26", X"04", X"03", X"03", X"02", X"03", X"03", X"1b", X"33", X"34", X"32", X"32", X"32", X"35", X"38", X"38", X"3b", X"3a", X"3a", X"3d", X"41", X"42", X"41", X"34", X"0c", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"22", X"34", X"3e", X"40", X"43", X"3a", X"3d", X"3e", X"3f", X"40", X"42", X"3e", X"3b", X"39", X"35", X"34", X"33", X"22", X"04", X"03", X"03", X"02", X"03", X"03", X"21", X"35", X"35", X"35", X"34", X"35", X"35", X"37", X"38", X"3a", X"3b", X"3a", X"3c", X"3a", X"39", X"3e", X"42", X"24", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"11", X"2a", X"3b", X"43", X"40", X"40", X"3a", X"3d", X"40", X"3f", X"41", X"40", X"3e", X"3b", X"38", X"38", X"35", X"32", X"1e", X"03", X"03", X"03", X"02", X"03", X"03", X"25", X"37", X"37", X"36", X"37", X"38", X"36", X"3b", X"3c", X"3d", X"3e", X"3f", X"3d", X"3b", X"3a", X"3f", X"43", X"3a", X"0b", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"05", X"1d", X"37", X"40", X"46", X"41", X"3f", X"3e", X"3e", X"40", X"3f", X"3f", X"3f", X"3a", X"3a", X"37", X"38", X"34", X"30", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"26", X"36", X"38", X"39", X"39", X"39", X"38", X"3e", X"3e", X"3e", X"42", X"41", X"3f", X"3c", X"3e", X"41", X"45", X"44", X"23", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0a", X"29", X"41", X"40", X"42", X"41", X"46", X"3e", X"41", X"42", X"40", X"3f", X"3f", X"3c", X"3b", X"38", X"36", X"34", X"2f", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"2c", X"38", X"3c", X"3d", X"3d", X"3d", X"3d", X"41", X"42", X"44", X"44", X"43", X"44", X"40", X"41", X"43", X"46", X"45", X"39", X"08", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"11", X"35", X"46", X"41", X"46", X"45", X"4a", X"44", X"46", X"44", X"42", X"3e", X"3f", X"3d", X"3b", X"39", X"36", X"35", X"31", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"31", X"39", X"3d", X"3f", X"40", X"40", X"41", X"40", X"46", X"47", X"48", X"46", X"46", X"44", X"44", X"45", X"49", X"48", X"42", X"18", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"05", X"1e", X"42", X"49", X"40", X"41", X"41", X"41", X"40", X"43", X"43", X"44", X"41", X"40", X"3f", X"3d", X"3b", X"37", X"37", X"32", X"18", X"03", X"03", X"03", X"02", X"03", X"04", X"36", X"3e", X"3f", X"40", X"3e", X"40", X"41", X"40", X"45", X"47", X"48", X"47", X"49", X"47", X"48", X"49", X"4a", X"49", X"45", X"2a", X"05", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"09", X"2f", X"44", X"46", X"3f", X"42", X"41", X"40", X"42", X"43", X"44", X"42", X"41", X"41", X"3d", X"3b", X"39", X"38", X"37", X"33", X"16", X"03", X"03", X"03", X"02", X"03", X"06", X"3a", X"42", X"42", X"41", X"42", X"3f", X"40", X"40", X"42", X"47", X"47", X"47", X"48", X"48", X"4a", X"4b", X"4f", X"4f", X"4a", X"39", X"0d", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"11", X"37", X"46", X"44", X"41", X"45", X"43", X"43", X"42", X"42", X"41", X"44", X"42", X"40", X"3d", X"3a", X"39", X"3b", X"38", X"35", X"14", X"03", X"03", X"03", X"02", X"03", X"08", X"49", X"4a", X"46", X"45", X"48", X"48", X"46", X"45", X"44", X"46", X"48", X"47", X"49", X"49", X"4b", X"4c", X"51", X"51", X"4f", X"3f", X"1e", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"17", X"43", X"46", X"41", X"41", X"43", X"43", X"42", X"43", X"42", X"42", X"42", X"41", X"41", X"3d", X"3b", X"39", X"3b", X"39", X"36", X"12", X"03", X"03", X"03", X"02", X"03", X"0c", X"4d", X"57", X"54", X"55", X"53", X"54", X"4c", X"4c", X"46", X"47", X"48", X"49", X"49", X"4a", X"4c", X"4d", X"52", X"58", X"4d", X"45", X"2a", X"06", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"07", X"1f", X"4a", X"46", X"44", X"43", X"46", X"45", X"44", X"44", X"43", X"42", X"45", X"43", X"40", X"3d", X"3c", X"3b", X"3e", X"3f", X"3c", X"13", X"03", X"03", X"03", X"02", X"03", X"11", X"4d", X"4e", X"4f", X"52", X"51", X"57", X"58", X"53", X"4f", X"4e", X"4d", X"4b", X"4c", X"4b", X"4f", X"53", X"5c", X"59", X"53", X"4b", X"38", X"0d", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"29", X"4f", X"49", X"47", X"47", X"47", X"45", X"46", X"44", X"44", X"44", X"45", X"43", X"43", X"41", X"43", X"47", X"47", X"45", X"46", X"15", X"03", X"03", X"03", X"02", X"03", X"17", X"50", X"4f", X"53", X"59", X"5e", X"5a", X"56", X"53", X"53", X"53", X"53", X"4e", X"4c", X"4c", X"58", X"77", X"7d", X"64", X"5a", X"4d", X"46", X"1b", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"3d", X"55", X"49", X"49", X"4a", X"4c", X"4a", X"48", X"45", X"45", X"47", X"46", X"44", X"46", X"4c", X"51", X"4b", X"49", X"49", X"46", X"12", X"03", X"03", X"03", X"02", X"03", X"1f", X"54", X"56", X"5a", X"62", X"6b", X"5d", X"56", X"56", X"58", X"5d", X"5c", X"56", X"50", X"4d", X"67", X"8f", X"85", X"6b", X"5f", X"4f", X"47", X"2d", X"07", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"12", X"65", X"56", X"4d", X"4c", X"4f", X"4f", X"51", X"51", X"50", X"52", X"52", X"4f", X"4e", X"52", X"53", X"54", X"54", X"52", X"51", X"4d", X"10", X"03", X"03", X"03", X"02", X"03", X"25", X"5b", X"5d", X"5d", X"60", X"60", X"5d", X"5b", X"59", X"57", X"56", X"57", X"5f", X"57", X"57", X"62", X"71", X"67", X"61", X"5e", X"4f", X"49", X"39", X"12", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"2b", X"78", X"55", X"51", X"52", X"53", X"5c", X"63", X"61", X"60", X"60", X"5d", X"5c", X"59", X"5a", X"59", X"59", X"5b", X"5a", X"59", X"53", X"0e", X"03", X"03", X"03", X"02", X"03", X"2e", X"63", X"60", X"62", X"62", X"62", X"61", X"5e", X"5c", X"5b", X"58", X"53", X"5b", X"5c", X"60", X"63", X"60", X"5c", X"5d", X"52", X"4a", X"46", X"40", X"2b", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"06", X"43", X"7a", X"54", X"53", X"58", X"63", X"67", X"67", X"69", X"6d", X"72", X"74", X"74", X"6f", X"6f", X"6d", X"6d", X"6a", X"6c", X"6a", X"63", X"0d", X"03", X"03", X"03", X"02", X"03", X"44", X"7a", X"77", X"7b", X"7d", X"77", X"68", X"64", X"61", X"5e", X"5a", X"55", X"53", X"58", X"5d", X"63", X"63", X"57", X"5c", X"5d", X"4d", X"44", X"45", X"4b", X"09", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0b", X"4f", X"7f", X"58", X"5a", X"68", X"65", X"6a", X"79", X"84", X"86", X"86", X"8a", X"8f", X"91", X"8e", X"8e", X"8c", X"8c", X"8f", X"8c", X"7e", X"0b", X"03", X"03", X"03", X"02", X"03", X"56", X"84", X"7b", X"7d", X"7b", X"7b", X"72", X"6d", X"66", X"62", X"5f", X"5d", X"56", X"54", X"5d", X"69", X"70", X"62", X"5b", X"66", X"50", X"45", X"4c", X"52", X"12", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0e", X"4f", X"87", X"65", X"66", X"67", X"6c", X"84", X"8b", X"84", X"83", X"83", X"88", X"8a", X"8d", X"95", X"95", X"8f", X"8a", X"86", X"83", X"72", X"08", X"03", X"03", X"03", X"03", X"04", X"57", X"73", X"73", X"76", X"75", X"77", X"76", X"72", X"6d", X"68", X"64", X"60", X"5e", X"5d", X"57", X"5a", X"65", X"62", X"59", X"59", X"51", X"44", X"5a", X"56", X"14", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0e", X"4e", X"92", X"76", X"6b", X"70", X"7b", X"84", X"83", X"80", X"82", X"84", X"86", X"8d", X"92", X"9c", X"9d", X"96", X"8c", X"8b", X"89", X"78", X"07", X"03", X"03", X"03", X"03", X"07", X"63", X"78", X"79", X"7b", X"7e", X"7f", X"7e", X"7c", X"76", X"6d", X"6a", X"66", X"61", X"63", X"60", X"5c", X"63", X"64", X"5b", X"58", X"50", X"4a", X"6c", X"53", X"11", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0d", X"4b", X"95", X"76", X"72", X"7f", X"85", X"88", X"87", X"88", X"8a", X"8c", X"92", X"99", X"a1", X"ab", X"a7", X"a1", X"9a", X"9f", X"a2", X"80", X"05", X"04", X"03", X"03", X"04", X"0a", X"71", X"80", X"81", X"82", X"85", X"87", X"85", X"81", X"7a", X"76", X"72", X"6b", X"66", X"65", X"67", X"61", X"62", X"67", X"62", X"5d", X"53", X"50", X"70", X"52", X"11", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0a", X"44", X"93", X"76", X"7d", X"89", X"88", X"8d", X"91", X"92", X"93", X"96", X"99", X"9f", X"ac", X"b6", X"b3", X"b0", X"ac", X"b7", X"bf", X"84", X"06", X"04", X"03", X"03", X"06", X"11", X"7b", X"8e", X"89", X"8b", X"8b", X"8e", X"8b", X"83", X"7e", X"79", X"76", X"6f", X"6b", X"68", X"67", X"6c", X"63", X"65", X"6d", X"65", X"59", X"57", X"72", X"4a", X"0c", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"09", X"3b", X"91", X"7b", X"83", X"8a", X"89", X"92", X"98", X"9c", X"9f", X"a0", X"a3", X"a3", X"ab", X"b6", X"b9", X"b6", X"b4", X"bc", X"c8", X"84", X"0a", X"06", X"04", X"03", X"08", X"1d", X"7d", X"95", X"98", X"95", X"96", X"98", X"90", X"89", X"83", X"7f", X"7d", X"77", X"71", X"6d", X"6b", X"70", X"70", X"69", X"6b", X"6d", X"6b", X"61", X"70", X"3f", X"09", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"06", X"2d", X"85", X"81", X"86", X"8c", X"90", X"9a", X"a0", X"a3", X"a5", X"a7", X"a8", X"ac", X"aa", X"b0", X"b3", X"b6", X"b3", X"b3", X"c2", X"85", X"17", X"0f", X"0a", X"0c", X"16", X"34", X"a5", X"ab", X"98", X"98", X"9f", X"9d", X"95", X"8e", X"88", X"87", X"85", X"81", X"7b", X"77", X"75", X"74", X"79", X"77", X"6f", X"6a", X"70", X"69", X"67", X"2d", X"05", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"1d", X"75", X"7f", X"81", X"91", X"93", X"97", X"9f", X"a3", X"a7", X"a8", X"ab", X"ab", X"a6", X"ad", X"b1", X"b1", X"af", X"ad", X"b3", X"9d", X"3a", X"24", X"1f", X"23", X"30", X"58", X"c9", X"e1", X"a5", X"96", X"a7", X"a3", X"9a", X"96", X"91", X"90", X"8e", X"8a", X"89", X"85", X"80", X"7e", X"7c", X"7b", X"79", X"71", X"6d", X"70", X"5a", X"16", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0f", X"62", X"78", X"7f", X"8a", X"86", X"8c", X"94", X"9a", X"a0", X"a4", X"a9", X"ab", X"a8", X"a8", X"aa", X"b7", X"a8", X"a6", X"ab", X"bc", X"71", X"52", X"41", X"49", X"6b", X"81", X"d5", X"ea", X"b3", X"97", X"a7", X"aa", X"a2", X"9a", X"9a", X"97", X"96", X"97", X"97", X"93", X"8a", X"87", X"82", X"7b", X"7b", X"77", X"6e", X"69", X"49", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0a", X"59", X"77", X"7b", X"78", X"73", X"7d", X"86", X"8b", X"92", X"a2", X"aa", X"ad", X"ac", X"aa", X"a8", X"b2", X"ae", X"a8", X"ac", X"c9", X"c3", X"8f", X"7a", X"75", X"9b", X"d2", X"fc", X"df", X"ae", X"9f", X"a9", X"ad", X"a7", X"a2", X"a2", X"a1", X"a1", X"a2", X"a4", X"a3", X"99", X"92", X"87", X"7f", X"78", X"76", X"6f", X"63", X"34", X"05", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0a", X"5f", X"7d", X"6f", X"69", X"6b", X"74", X"79", X"7e", X"88", X"9c", X"ae", X"b2", X"b1", X"b0", X"b0", X"bf", X"c2", X"be", X"c2", X"dc", X"f9", X"ec", X"de", X"da", X"f5", X"fe", X"fb", X"dc", X"bb", X"b8", X"b2", X"b3", X"b2", X"b0", X"ad", X"aa", X"ad", X"ad", X"b1", X"b1", X"a6", X"9d", X"90", X"83", X"7c", X"70", X"6d", X"6a", X"3b", X"03", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"64", X"88", X"69", X"68", X"6d", X"72", X"77", X"7b", X"88", X"a1", X"b5", X"bb", X"b9", X"b7", X"c0", X"d4", X"d1", X"d5", X"dd", X"e6", X"f1", X"fb", X"ff", X"ff", X"ff", X"ff", X"fb", X"e7", X"e7", X"e8", X"df", X"d5", X"cd", X"c4", X"b9", X"b9", X"ba", X"b8", X"bc", X"b3", X"a8", X"9e", X"91", X"7e", X"7a", X"73", X"6a", X"73", X"52", X"04", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"07", X"47", X"93", X"6c", X"70", X"74", X"75", X"7d", X"84", X"99", X"b3", X"c6", X"d1", X"cd", X"c8", X"cd", X"d8", X"de", X"de", X"dc", X"dc", X"dd", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fd", X"fe", X"fd", X"fa", X"f1", X"dc", X"c9", X"c6", X"c5", X"c2", X"bd", X"b6", X"a7", X"99", X"8f", X"83", X"73", X"6e", X"6a", X"7b", X"5c", X"07", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"26", X"7f", X"89", X"76", X"79", X"7b", X"7c", X"84", X"92", X"aa", X"ca", X"d6", X"cf", X"ca", X"cf", X"da", X"de", X"e3", X"e2", X"dd", X"da", X"eb", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f7", X"f5", X"ef", X"eb", X"e3", X"da", X"d1", X"ce", X"cb", X"c8", X"c4", X"b5", X"a7", X"98", X"8d", X"7f", X"70", X"72", X"97", X"60", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"0b", X"49", X"7d", X"72", X"78", X"7d", X"7b", X"7a", X"81", X"94", X"ab", X"ac", X"a0", X"a5", X"bb", X"d2", X"e4", X"ee", X"ea", X"de", X"db", X"ea", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fc", X"fa", X"fa", X"f5", X"f1", X"e8", X"e4", X"e0", X"dd", X"de", X"dc", X"d3", X"c5", X"b4", X"9f", X"92", X"87", X"7d", X"9e", X"49", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"1c", X"5b", X"61", X"77", X"86", X"8d", X"87", X"8e", X"94", X"90", X"90", X"8c", X"94", X"a5", X"bf", X"d6", X"ee", X"e8", X"dc", X"de", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fa", X"f5", X"ea", X"ea", X"ea", X"e9", X"e5", X"e7", X"eb", X"ee", X"e6", X"dc", X"ce", X"b6", X"a3", X"95", X"86", X"84", X"2c", X"04", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"31", X"58", X"6b", X"84", X"92", X"96", X"96", X"9a", X"92", X"98", X"8e", X"91", X"9d", X"b2", X"ce", X"e3", X"e3", X"e1", X"ea", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"ea", X"da", X"d2", X"d5", X"db", X"d9", X"df", X"e3", X"ec", X"ed", X"ee", X"ef", X"e0", X"c7", X"a2", X"9e", X"70", X"1b", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"10", X"44", X"76", X"7d", X"87", X"8a", X"91", X"9d", X"9e", X"9f", X"9a", X"92", X"9b", X"b3", X"cd", X"df", X"e7", X"ee", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fc", X"fe", X"ff", X"fa", X"e8", X"d7", X"c9", X"c7", X"d0", X"e7", X"f4", X"f1", X"f7", X"ef", X"e8", X"f0", X"d6", X"ba", X"bf", X"af", X"3a", X"07", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"22", X"67", X"7b", X"6d", X"6b", X"79", X"97", X"a0", X"a5", X"a3", X"9e", X"a2", X"b6", X"ce", X"e1", X"eb", X"f7", X"fc", X"fe", X"ff", X"ff", X"fe", X"f5", X"dd", X"e0", X"f3", X"fe", X"fe", X"ec", X"d5", X"cd", X"d2", X"f5", X"fc", X"f2", X"df", X"f0", X"d8", X"d7", X"c5", X"a2", X"a2", X"ae", X"3f", X"0f", X"04", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"14", X"35", X"57", X"59", X"5e", X"6a", X"6d", X"85", X"98", X"a8", X"a7", X"b3", X"bf", X"c7", X"d2", X"e6", X"ca", X"c2", X"d9", X"e7", X"de", X"c0", X"b8", X"b1", X"cb", X"e7", X"e4", X"e4", X"d1", X"c7", X"ea", X"fe", X"f9", X"e9", X"e9", X"cd", X"b3", X"ae", X"9f", X"82", X"90", X"48", X"0c", X"04", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"08", X"19", X"2d", X"3c", X"49", X"5d", X"66", X"7a", X"94", X"93", X"92", X"98", X"9a", X"ad", X"b3", X"9c", X"8f", X"93", X"a4", X"9f", X"9c", X"aa", X"a2", X"9c", X"a6", X"a1", X"a2", X"9f", X"a6", X"c6", X"f9", X"f6", X"ef", X"ce", X"a2", X"8f", X"87", X"69", X"4e", X"34", X"0a", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"18", X"2a", X"46", X"53", X"6f", X"76", X"75", X"7c", X"7f", X"77", X"79", X"78", X"76", X"7d", X"8a", X"98", X"99", X"a0", X"96", X"8f", X"85", X"7a", X"78", X"83", X"87", X"96", X"a8", X"c5", X"d0", X"cb", X"ba", X"87", X"6f", X"52", X"31", X"14", X"04", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"0f", X"23", X"25", X"23", X"3a", X"48", X"56", X"64", X"67", X"6d", X"6e", X"6d", X"71", X"79", X"7a", X"7c", X"83", X"81", X"78", X"6e", X"68", X"5d", X"6b", X"72", X"8a", X"a7", X"93", X"a8", X"bc", X"9b", X"6d", X"2a", X"10", X"06", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"04", X"06", X"05", X"0a", X"13", X"16", X"1f", X"2c", X"3b", X"48", X"4b", X"4d", X"57", X"5f", X"62", X"64", X"64", X"5c", X"52", X"4a", X"43", X"48", X"3e", X"41", X"45", X"3b", X"31", X"23", X"18", X"0d", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"0a", X"0c", X"12", X"21", X"30", X"2b", X"37", X"42", X"39", X"2c", X"27", X"1f", X"1c", X"16", X"14", X"0f", X"0e", X"0b", X"07", X"07", X"07", X"05", X"05", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"03", X"05", X"07", X"0d", X"10", X"0d", X"0e", X"0c", X"0a", X"06", X"04", X"06", X"03", X"03", X"03", X"05", X"03", X"03", X"04", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"));
  

  constant imagem_teste1 : MatrizImagem := ((X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"08", X"1b", X"27", X"20", X"17", X"12", X"09", X"0a", X"07", X"04", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"08", X"25", X"34", X"34", X"31", X"33", X"2d", X"27", X"25", X"22", X"19", X"0b", X"18", X"18", X"14", X"0e", X"03", X"03", X"03", X"02", X"03", X"03", X"06", X"11", X"1d", X"23", X"27", X"28", X"23", X"23", X"21", X"22", X"1f", X"1e", X"1d", X"12", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"05", X"22", X"34", X"3a", X"36", X"34", X"33", X"31", X"2e", X"2f", X"2b", X"29", X"26", X"27", X"27", X"26", X"20", X"03", X"03", X"03", X"02", X"03", X"03", X"13", X"2c", X"30", X"42", X"59", X"6c", X"6f", X"6e", X"69", X"63", X"5d", X"54", X"51", X"4e", X"35", X"0b", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"18", X"35", X"35", X"37", X"33", X"33", X"33", X"32", X"2f", X"2f", X"2e", X"2e", X"2d", X"2e", X"2d", X"2d", X"29", X"04", X"03", X"03", X"02", X"03", X"03", X"1b", X"33", X"34", X"36", X"3a", X"4b", X"69", X"7b", X"7e", X"79", X"72", X"6a", X"62", X"5d", X"5c", X"39", X"07", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0b", X"3b", X"36", X"35", X"36", X"35", X"37", X"35", X"37", X"32", X"32", X"31", X"31", X"31", X"31", X"33", X"36", X"2d", X"03", X"03", X"03", X"02", X"03", X"03", X"24", X"39", X"39", X"3a", X"3e", X"3d", X"41", X"51", X"65", X"70", X"76", X"75", X"73", X"6c", X"67", X"5e", X"23", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"25", X"46", X"39", X"36", X"37", X"39", X"3a", X"37", X"35", X"33", X"35", X"35", X"37", X"35", X"33", X"33", X"34", X"26", X"03", X"03", X"03", X"02", X"03", X"03", X"2b", X"42", X"45", X"4a", X"49", X"4a", X"4f", X"53", X"4d", X"4b", X"4c", X"57", X"65", X"6d", X"6d", X"66", X"3c", X"0c", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0a", X"35", X"3d", X"3d", X"38", X"37", X"38", X"3a", X"39", X"38", X"37", X"3a", X"3d", X"48", X"39", X"35", X"35", X"35", X"24", X"03", X"03", X"03", X"02", X"03", X"03", X"35", X"4a", X"4a", X"4f", X"54", X"58", X"50", X"4d", X"4a", X"47", X"41", X"41", X"44", X"47", X"4c", X"4f", X"41", X"22", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"18", X"36", X"3b", X"3b", X"37", X"38", X"37", X"3a", X"3c", X"40", X"3e", X"40", X"43", X"46", X"3d", X"3c", X"37", X"36", X"23", X"03", X"03", X"03", X"02", X"03", X"04", X"3d", X"4d", X"4d", X"51", X"52", X"55", X"4b", X"4e", X"48", X"43", X"43", X"45", X"44", X"42", X"40", X"44", X"44", X"39", X"0d", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"25", X"3e", X"3c", X"3b", X"38", X"3a", X"3c", X"3e", X"41", X"3f", X"40", X"47", X"42", X"3f", X"3d", X"3e", X"3c", X"3b", X"23", X"03", X"03", X"03", X"02", X"03", X"04", X"41", X"4e", X"50", X"57", X"52", X"4e", X"4b", X"4e", X"51", X"43", X"45", X"46", X"45", X"44", X"45", X"47", X"49", X"45", X"26", X"04", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0c", X"31", X"44", X"3a", X"3c", X"3b", X"3e", X"41", X"42", X"41", X"42", X"46", X"4a", X"42", X"40", X"40", X"43", X"42", X"43", X"24", X"03", X"03", X"03", X"02", X"03", X"06", X"4d", X"54", X"54", X"59", X"58", X"53", X"4e", X"4d", X"52", X"4f", X"44", X"44", X"48", X"47", X"48", X"49", X"4f", X"48", X"3d", X"0b", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"14", X"38", X"3e", X"3b", X"42", X"42", X"3f", X"40", X"43", X"45", X"46", X"48", X"46", X"42", X"42", X"46", X"46", X"48", X"47", X"23", X"03", X"03", X"03", X"02", X"03", X"08", X"59", X"58", X"55", X"58", X"5a", X"57", X"53", X"4c", X"50", X"59", X"55", X"47", X"46", X"49", X"4a", X"4a", X"5a", X"52", X"48", X"20", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"06", X"20", X"41", X"3e", X"3d", X"41", X"41", X"3f", X"40", X"44", X"46", X"49", X"49", X"46", X"46", X"47", X"49", X"46", X"48", X"45", X"1e", X"03", X"03", X"03", X"02", X"03", X"0a", X"62", X"5b", X"5a", X"5d", X"5a", X"54", X"52", X"4c", X"4d", X"4d", X"4f", X"4d", X"53", X"4e", X"4d", X"4e", X"57", X"60", X"4e", X"3c", X"0b", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"09", X"2e", X"41", X"41", X"44", X"42", X"40", X"40", X"43", X"46", X"48", X"48", X"48", X"48", X"47", X"4a", X"47", X"47", X"4a", X"4b", X"1e", X"03", X"03", X"03", X"02", X"03", X"10", X"63", X"5e", X"61", X"61", X"58", X"50", X"50", X"4d", X"4b", X"4e", X"4a", X"49", X"4e", X"4d", X"4b", X"4d", X"50", X"58", X"58", X"5b", X"27", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"12", X"36", X"44", X"45", X"42", X"43", X"42", X"43", X"43", X"46", X"47", X"4a", X"4a", X"4c", X"4e", X"4c", X"4b", X"50", X"54", X"57", X"1f", X"03", X"03", X"03", X"02", X"03", X"15", X"68", X"65", X"65", X"5e", X"57", X"53", X"52", X"54", X"4e", X"4d", X"4d", X"4b", X"4c", X"4d", X"51", X"50", X"52", X"54", X"5c", X"64", X"45", X"08", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"19", X"3d", X"44", X"42", X"3e", X"41", X"41", X"42", X"45", X"48", X"4b", X"4b", X"4f", X"54", X"53", X"54", X"54", X"5c", X"61", X"5a", X"1c", X"03", X"03", X"03", X"02", X"03", X"1e", X"72", X"6a", X"65", X"64", X"5b", X"57", X"57", X"56", X"50", X"4e", X"4e", X"52", X"4f", X"4d", X"57", X"53", X"53", X"52", X"54", X"58", X"55", X"19", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"08", X"1f", X"41", X"43", X"42", X"3f", X"43", X"42", X"43", X"49", X"4e", X"4e", X"55", X"5b", X"5a", X"5d", X"62", X"65", X"69", X"61", X"64", X"1b", X"03", X"03", X"03", X"02", X"03", X"26", X"77", X"71", X"6e", X"72", X"67", X"63", X"5c", X"57", X"53", X"50", X"50", X"52", X"53", X"4f", X"4f", X"51", X"4f", X"50", X"56", X"59", X"56", X"29", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"26", X"47", X"4a", X"47", X"45", X"44", X"45", X"4d", X"50", X"51", X"58", X"60", X"65", X"68", X"70", X"75", X"70", X"68", X"68", X"68", X"17", X"03", X"03", X"03", X"02", X"03", X"31", X"80", X"78", X"7d", X"78", X"72", X"69", X"60", X"5a", X"5a", X"56", X"52", X"4f", X"51", X"50", X"52", X"53", X"52", X"55", X"55", X"59", X"57", X"3a", X"06", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0c", X"41", X"5e", X"54", X"50", X"4d", X"50", X"52", X"52", X"52", X"5a", X"64", X"6a", X"6c", X"74", X"81", X"82", X"73", X"6a", X"6a", X"68", X"10", X"03", X"03", X"03", X"02", X"04", X"3c", X"82", X"7c", X"81", X"7a", X"7d", X"6d", X"61", X"5f", X"5d", X"5d", X"5b", X"58", X"53", X"4f", X"4e", X"4f", X"50", X"54", X"54", X"56", X"57", X"46", X"0c", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"15", X"6a", X"61", X"5a", X"53", X"54", X"55", X"59", X"58", X"5d", X"69", X"71", X"75", X"76", X"7f", X"85", X"81", X"76", X"6f", X"6e", X"67", X"0e", X"03", X"03", X"03", X"03", X"04", X"43", X"82", X"7d", X"7e", X"86", X"88", X"75", X"6c", X"68", X"64", X"60", X"5d", X"5a", X"54", X"50", X"50", X"51", X"51", X"51", X"54", X"54", X"57", X"4c", X"18", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"2e", X"78", X"58", X"5c", X"56", X"56", X"5e", X"65", X"65", X"6b", X"75", X"7d", X"85", X"88", X"8a", X"84", X"7e", X"78", X"71", X"6d", X"63", X"0b", X"03", X"03", X"03", X"02", X"04", X"4c", X"86", X"82", X"85", X"8c", X"8a", X"7d", X"73", X"6b", X"66", X"60", X"5a", X"58", X"55", X"54", X"55", X"54", X"54", X"51", X"57", X"52", X"52", X"4d", X"32", X"04", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"07", X"45", X"7a", X"57", X"5d", X"5c", X"60", X"6b", X"75", X"76", X"77", X"82", X"8c", X"92", X"92", X"8d", X"86", X"82", X"7e", X"7b", X"75", X"66", X"09", X"03", X"03", X"03", X"03", X"05", X"59", X"86", X"88", X"8b", X"8e", X"8e", X"87", X"86", X"7a", X"6b", X"63", X"5d", X"5a", X"5a", X"59", X"58", X"5a", X"56", X"53", X"57", X"58", X"52", X"50", X"4c", X"0a", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0c", X"4f", X"81", X"64", X"5e", X"61", X"6a", X"7d", X"86", X"83", X"83", X"8b", X"94", X"97", X"98", X"93", X"8f", X"8c", X"8a", X"88", X"83", X"6a", X"06", X"03", X"03", X"03", X"03", X"09", X"63", X"85", X"8c", X"90", X"90", X"94", X"90", X"94", X"8e", X"79", X"6c", X"65", X"5e", X"60", X"5f", X"5f", X"5d", X"5b", X"57", X"55", X"59", X"56", X"52", X"54", X"10", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"10", X"50", X"88", X"74", X"60", X"68", X"72", X"7e", X"8a", X"93", X"8e", X"8f", X"98", X"9d", X"9f", X"9e", X"9a", X"9c", X"9c", X"95", X"8b", X"6a", X"05", X"04", X"03", X"03", X"05", X"0d", X"6e", X"88", X"90", X"90", X"8c", X"8f", X"91", X"98", X"98", X"84", X"75", X"6d", X"69", X"67", X"64", X"61", X"60", X"5d", X"5a", X"58", X"59", X"53", X"53", X"57", X"12", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"10", X"51", X"91", X"80", X"69", X"74", X"78", X"81", X"8c", X"96", X"94", X"96", X"9c", X"a6", X"a9", X"ab", X"ab", X"b1", X"ad", X"a3", X"93", X"6a", X"05", X"04", X"04", X"03", X"06", X"13", X"7c", X"8e", X"92", X"8e", X"91", X"95", X"92", X"93", X"9d", X"95", X"87", X"7b", X"73", X"6f", X"6a", X"6a", X"69", X"61", X"5f", X"5b", X"59", X"56", X"58", X"54", X"0d", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0f", X"4c", X"95", X"7a", X"73", X"78", X"7d", X"8c", X"95", X"9d", X"a1", X"a1", X"a8", X"b2", X"b9", X"bd", X"bd", X"c3", X"bc", X"ab", X"96", X"64", X"06", X"06", X"05", X"05", X"0b", X"1c", X"85", X"91", X"94", X"8f", X"8c", X"8d", X"8b", X"90", X"93", X"98", X"8e", X"84", X"7f", X"78", X"72", X"75", X"76", X"6c", X"67", X"62", X"5c", X"56", X"5a", X"53", X"0d", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0b", X"45", X"92", X"7d", X"76", X"74", X"78", X"8b", X"9c", X"a6", X"ae", X"b8", X"b5", X"be", X"c6", X"cb", X"ca", X"cb", X"c6", X"ae", X"98", X"5d", X"09", X"08", X"07", X"08", X"13", X"2e", X"90", X"9c", X"9e", X"9b", X"93", X"91", X"8c", X"8b", X"96", X"92", X"8f", X"8a", X"85", X"7f", X"7a", X"7d", X"7a", X"76", X"73", X"69", X"5d", X"54", X"60", X"4b", X"09", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0a", X"3c", X"91", X"83", X"70", X"76", X"78", X"87", X"98", X"a4", X"b0", X"c1", X"cb", X"c8", X"cf", X"d1", X"d1", X"d3", X"ca", X"b2", X"9e", X"5e", X"10", X"0f", X"11", X"14", X"1d", X"3f", X"9e", X"aa", X"b3", X"b3", X"aa", X"a2", X"96", X"92", X"a1", X"9e", X"9d", X"95", X"8d", X"84", X"7f", X"7f", X"7e", X"7c", X"7a", X"74", X"68", X"5c", X"69", X"3d", X"08", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"07", X"2f", X"83", X"a9", X"8e", X"81", X"7a", X"88", X"93", X"9d", X"b1", X"c5", X"ce", X"d2", X"cf", X"d6", X"d6", X"da", X"d1", X"b5", X"a6", X"72", X"23", X"1f", X"21", X"2a", X"37", X"5a", X"cb", X"c3", X"cc", X"cd", X"c4", X"b4", X"a8", X"a8", X"aa", X"a9", X"a9", X"9e", X"90", X"8b", X"8a", X"7f", X"7c", X"7b", X"7a", X"76", X"75", X"68", X"6a", X"2a", X"05", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"20", X"77", X"b7", X"a4", X"a8", X"86", X"96", X"a6", X"b1", X"bc", X"c7", X"d3", X"da", X"d7", X"dc", X"dc", X"df", X"d9", X"bd", X"ac", X"93", X"48", X"46", X"52", X"66", X"87", X"c2", X"fd", X"ea", X"f0", X"ef", X"df", X"cc", X"c1", X"bc", X"b6", X"b5", X"b1", X"a6", X"a2", X"99", X"99", X"8e", X"85", X"80", X"7c", X"78", X"74", X"77", X"5d", X"16", X"04", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"12", X"65", X"b5", X"ae", X"be", X"b0", X"b6", X"bf", X"c8", X"cb", X"d1", X"db", X"e6", X"eb", X"e8", X"e6", X"e5", X"e0", X"c9", X"bd", X"df", X"b3", X"d3", X"e7", X"f4", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ee", X"de", X"ce", X"c5", X"bd", X"b9", X"b5", X"b4", X"ab", X"a6", X"a0", X"98", X"8d", X"87", X"80", X"77", X"71", X"49", X"09", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0d", X"5e", X"b6", X"b8", X"d2", X"dd", X"c9", X"cf", X"d8", X"e1", X"e3", X"e7", X"f2", X"f7", X"fa", X"f6", X"f4", X"f3", X"e2", X"d8", X"fe", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f0", X"db", X"ce", X"c2", X"bc", X"bf", X"be", X"b8", X"b3", X"b7", X"a6", X"9e", X"8e", X"89", X"7c", X"6e", X"35", X"06", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0e", X"6a", X"c0", X"be", X"d7", X"d7", X"d3", X"df", X"eb", X"f7", X"fd", X"fb", X"fc", X"fc", X"fe", X"fe", X"fe", X"fe", X"fe", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"eb", X"d9", X"cb", X"c3", X"c2", X"c2", X"c3", X"bb", X"b4", X"ab", X"9b", X"98", X"8b", X"80", X"78", X"47", X"04", X"03", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"12", X"79", X"b3", X"ac", X"da", X"f6", X"e4", X"f1", X"f7", X"fd", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f5", X"e6", X"d8", X"d0", X"d4", X"d2", X"cc", X"c5", X"b6", X"9f", X"99", X"90", X"82", X"7f", X"69", X"07", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0d", X"6a", X"a2", X"8a", X"b4", X"f3", X"f2", X"fa", X"fb", X"fd", X"fd", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"ee", X"e4", X"df", X"dd", X"d6", X"df", X"c1", X"aa", X"a3", X"99", X"8f", X"92", X"83", X"0a", X"03", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"06", X"46", X"7b", X"73", X"8a", X"d6", X"eb", X"f1", X"fe", X"fb", X"f3", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fa", X"ee", X"e5", X"e5", X"e4", X"df", X"be", X"b1", X"a6", X"99", X"94", X"98", X"90", X"0c", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"18", X"5e", X"63", X"6f", X"be", X"e2", X"ed", X"fb", X"f6", X"ed", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f3", X"e7", X"ee", X"fe", X"fc", X"d3", X"b2", X"ac", X"a2", X"99", X"b6", X"72", X"0a", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"09", X"3d", X"64", X"64", X"b0", X"c7", X"e6", X"f3", X"f1", X"f3", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f0", X"e4", X"f6", X"ff", X"fe", X"e3", X"ae", X"9d", X"94", X"93", X"c1", X"47", X"04", X"03", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"05", X"1c", X"50", X"6e", X"9f", X"ba", X"cf", X"e4", X"e7", X"f7", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f0", X"e0", X"ea", X"fd", X"ff", X"e8", X"ae", X"8b", X"83", X"9b", X"9f", X"2a", X"04", X"03", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"08", X"2e", X"6e", X"90", X"b9", X"c0", X"cd", X"d9", X"f6", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"da", X"d0", X"ee", X"fe", X"f5", X"b3", X"87", X"8b", X"8f", X"4b", X"0b", X"03", X"02", X"04", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"0a", X"39", X"75", X"b4", X"d9", X"cb", X"d3", X"dd", X"f6", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"d3", X"b9", X"c0", X"dc", X"d7", X"a2", X"86", X"88", X"49", X"14", X"05", X"03", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"09", X"2b", X"82", X"f3", X"f6", X"e4", X"d9", X"ec", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"e7", X"b8", X"9a", X"8b", X"9a", X"9a", X"78", X"66", X"44", X"16", X"05", X"03", X"03", X"03", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"08", X"1f", X"48", X"79", X"8a", X"c3", X"c7", X"e8", X"fc", X"fe", X"fa", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fe", X"fe", X"ff", X"fe", X"fd", X"fa", X"f9", X"df", X"bf", X"96", X"95", X"9f", X"70", X"5c", X"42", X"23", X"0a", X"05", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"0a", X"17", X"37", X"63", X"96", X"c4", X"d2", X"e6", X"f7", X"fa", X"fe", X"ff", X"ff", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f5", X"ea", X"e4", X"f5", X"f6", X"db", X"c9", X"c2", X"b3", X"a7", X"9c", X"a9", X"94", X"47", X"2e", X"17", X"06", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"04", X"09", X"13", X"24", X"41", X"5d", X"82", X"a2", X"cd", X"f6", X"ff", X"ff", X"fe", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"df", X"d8", X"d5", X"e8", X"ed", X"db", X"c3", X"a6", X"93", X"84", X"65", X"48", X"2f", X"13", X"0a", X"06", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"08", X"0f", X"14", X"1f", X"37", X"5d", X"bd", X"c9", X"e3", X"fa", X"fd", X"fe", X"ff", X"ff", X"ff", X"ff", X"fe", X"f9", X"d5", X"c0", X"ba", X"af", X"8f", X"6b", X"5b", X"49", X"37", X"26", X"18", X"0f", X"08", X"04", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"03", X"04", X"06", X"07", X"0c", X"18", X"20", X"2a", X"4b", X"56", X"8f", X"cd", X"e7", X"e5", X"f8", X"f0", X"d6", X"b7", X"94", X"6f", X"6d", X"62", X"40", X"29", X"25", X"17", X"13", X"11", X"10", X"09", X"09", X"04", X"03", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"06", X"09", X"0b", X"0e", X"1c", X"21", X"42", X"4c", X"60", X"68", X"b1", X"ba", X"59", X"47", X"35", X"2f", X"2b", X"1e", X"11", X"0f", X"14", X"08", X"09", X"09", X"05", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"04", X"04", X"05", X"07", X"09", X"0e", X"17", X"1a", X"21", X"25", X"24", X"27", X"21", X"14", X"0d", X"0e", X"0d", X"07", X"06", X"06", X"04", X"04", X"03", X"04", X"03", X"04", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"05", X"06", X"0b", X"0a", X"11", X"13", X"1b", X"15", X"0e", X"0c", X"06", X"05", X"04", X"04", X"04", X"03", X"03", X"04", X"03", X"03", X"02", X"04", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"04", X"05", X"06", X"09", X"07", X"05", X"06", X"04", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"03", X"04", X"03", X"04", X"04", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", x"03"));
  
  constant imagem_teste2 : MatrizImagem := ((X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"15", X"1d", X"1d", X"17", X"16", X"0d", X"14", X"0f", X"06", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"1e", X"2c", X"32", X"34", X"35", X"35", X"35", X"40", X"2e", X"1e", X"10", X"1b", X"1b", X"17", X"0f", X"03", X"03", X"03", X"02", X"03", X"03", X"08", X"0f", X"0e", X"0e", X"0f", X"13", X"19", X"27", X"27", X"28", X"23", X"21", X"1d", X"0e", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"05", X"1b", X"2d", X"3e", X"3d", X"3a", X"39", X"38", X"35", X"37", X"32", X"31", X"2f", X"2e", X"2f", X"2d", X"21", X"03", X"03", X"03", X"02", X"03", X"03", X"1d", X"38", X"30", X"30", X"31", X"33", X"34", X"42", X"5f", X"6f", X"6b", X"5f", X"56", X"47", X"21", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"12", X"2d", X"38", X"44", X"41", X"38", X"37", X"36", X"35", X"36", X"35", X"39", X"36", X"35", X"32", X"31", X"21", X"03", X"03", X"03", X"02", X"03", X"03", X"27", X"41", X"3d", X"3d", X"3d", X"3c", X"3a", X"3c", X"41", X"59", X"76", X"7a", X"6c", X"5f", X"4b", X"1a", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"08", X"24", X"36", X"3c", X"41", X"3e", X"39", X"37", X"3c", X"3d", X"3e", X"44", X"3c", X"39", X"35", X"37", X"37", X"22", X"03", X"03", X"03", X"02", X"03", X"03", X"31", X"41", X"41", X"43", X"46", X"43", X"3d", X"3b", X"3e", X"44", X"4c", X"6b", X"7e", X"73", X"63", X"47", X"0e", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"18", X"2f", X"3a", X"3b", X"3f", X"3c", X"3c", X"3e", X"41", X"47", X"48", X"58", X"43", X"3b", X"39", X"39", X"37", X"1f", X"03", X"03", X"03", X"02", X"03", X"04", X"37", X"3e", X"3f", X"3f", X"41", X"40", X"43", X"42", X"42", X"48", X"48", X"4d", X"69", X"7a", X"71", X"61", X"31", X"07", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"09", X"28", X"36", X"3b", X"3c", X"3d", X"3f", X"41", X"40", X"40", X"42", X"44", X"47", X"44", X"40", X"3d", X"3f", X"3e", X"1e", X"03", X"03", X"03", X"02", X"03", X"04", X"39", X"3f", X"3f", X"3e", X"3f", X"3f", X"3f", X"45", X"48", X"4b", X"4b", X"47", X"50", X"58", X"63", X"67", X"51", X"1c", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"15", X"31", X"38", X"3e", X"40", X"41", X"3f", X"42", X"45", X"43", X"46", X"46", X"46", X"45", X"44", X"46", X"44", X"40", X"1c", X"03", X"03", X"03", X"02", X"03", X"06", X"42", X"45", X"45", X"45", X"45", X"44", X"40", X"44", X"46", X"4a", X"49", X"4c", X"4e", X"4b", X"47", X"4b", X"49", X"37", X"0b", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"22", X"3a", X"3c", X"45", X"45", X"45", X"46", X"47", X"4a", X"4a", X"49", X"49", X"45", X"48", X"48", X"48", X"45", X"40", X"18", X"03", X"03", X"03", X"02", X"03", X"09", X"45", X"4b", X"4a", X"4d", X"4b", X"49", X"46", X"48", X"47", X"4b", X"4e", X"4c", X"4d", X"4c", X"49", X"46", X"46", X"43", X"24", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0b", X"2e", X"3d", X"40", X"47", X"46", X"4b", X"4e", X"4f", X"4f", X"50", X"4c", X"4c", X"4a", X"4a", X"49", X"47", X"45", X"3f", X"16", X"03", X"03", X"03", X"02", X"03", X"0c", X"43", X"46", X"4a", X"4d", X"4f", X"4f", X"4e", X"51", X"4e", X"50", X"55", X"4f", X"51", X"50", X"54", X"4a", X"46", X"45", X"39", X"09", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"14", X"3a", X"40", X"44", X"49", X"4d", X"56", X"57", X"58", X"59", X"55", X"4e", X"4d", X"4a", X"48", X"49", X"47", X"47", X"41", X"15", X"03", X"03", X"03", X"02", X"03", X"0f", X"41", X"41", X"47", X"4b", X"4f", X"50", X"55", X"55", X"51", X"52", X"58", X"54", X"53", X"55", X"5a", X"55", X"4e", X"49", X"45", X"1b", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"06", X"22", X"4a", X"45", X"47", X"4b", X"55", X"5f", X"5b", X"5d", X"5c", X"56", X"50", X"4d", X"4c", X"4a", X"4a", X"49", X"49", X"42", X"11", X"03", X"03", X"03", X"02", X"03", X"12", X"43", X"45", X"49", X"4d", X"4d", X"4f", X"52", X"57", X"54", X"51", X"57", X"58", X"56", X"56", X"59", X"5b", X"5c", X"50", X"48", X"30", X"06", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"09", X"2d", X"46", X"4b", X"4e", X"56", X"59", X"60", X"64", X"5f", X"5d", X"54", X"4f", X"4d", X"4a", X"4a", X"4a", X"4b", X"4b", X"45", X"0f", X"03", X"03", X"03", X"02", X"03", X"19", X"45", X"47", X"4b", X"4e", X"51", X"50", X"4f", X"53", X"53", X"55", X"56", X"55", X"57", X"57", X"5a", X"59", X"55", X"51", X"4d", X"41", X"12", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"12", X"35", X"4d", X"50", X"55", X"5b", X"58", X"59", X"5e", X"5e", X"5b", X"57", X"4f", X"4d", X"4c", X"4b", X"4c", X"50", X"4e", X"4a", X"0c", X"03", X"03", X"03", X"02", X"03", X"1e", X"49", X"4b", X"4e", X"52", X"55", X"54", X"52", X"55", X"54", X"54", X"59", X"54", X"58", X"58", X"5b", X"5b", X"57", X"51", X"51", X"49", X"24", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"18", X"3b", X"4e", X"52", X"56", X"58", X"58", X"58", X"5c", X"5d", X"5b", X"56", X"4f", X"4e", X"4c", X"4e", X"4e", X"52", X"52", X"4b", X"0a", X"04", X"03", X"03", X"02", X"03", X"24", X"49", X"4b", X"4f", X"54", X"55", X"57", X"57", X"55", X"52", X"55", X"56", X"57", X"5b", X"57", X"5c", X"5c", X"59", X"55", X"50", X"4d", X"35", X"06", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"08", X"1f", X"46", X"52", X"55", X"55", X"5b", X"5a", X"57", X"58", X"5b", X"5d", X"59", X"53", X"4e", X"4e", X"50", X"51", X"56", X"57", X"4f", X"08", X"03", X"03", X"03", X"02", X"03", X"2b", X"4e", X"4f", X"53", X"58", X"58", X"5e", X"5d", X"5a", X"57", X"58", X"59", X"59", X"61", X"58", X"5a", X"5d", X"5a", X"56", X"56", X"4f", X"47", X"11", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"0d", X"2b", X"54", X"56", X"56", X"59", X"5d", X"5b", X"59", X"57", X"58", X"5d", X"5f", X"55", X"53", X"53", X"55", X"5b", X"5e", X"60", X"52", X"06", X"03", X"03", X"03", X"02", X"03", X"34", X"55", X"56", X"58", X"5d", X"5f", X"62", X"63", X"60", X"5e", X"5d", X"5c", X"5c", X"62", X"58", X"5a", X"5c", X"5c", X"59", X"58", X"52", X"52", X"29", X"04", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"0d", X"44", X"5b", X"56", X"58", X"5e", X"62", X"5e", X"5a", X"58", X"59", X"5a", X"5e", X"5b", X"56", X"5b", X"62", X"63", X"65", X"68", X"57", X"04", X"03", X"03", X"03", X"02", X"04", X"42", X"5f", X"62", X"64", X"64", X"68", X"68", X"66", X"66", X"63", X"62", X"61", X"65", X"62", X"58", X"58", X"5a", X"5a", X"58", X"56", X"54", X"56", X"41", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"16", X"6a", X"5c", X"5a", X"5d", X"64", X"64", X"62", X"5e", X"5c", X"5e", X"5d", X"5b", X"6c", X"6a", X"6a", X"6a", X"6d", X"69", X"72", X"5c", X"04", X"04", X"03", X"03", X"03", X"04", X"4a", X"65", X"6c", X"6f", X"71", X"6f", X"6d", X"6d", X"70", X"6c", X"64", X"66", X"69", X"5c", X"57", X"59", X"5b", X"5b", X"57", X"54", X"55", X"5b", X"4e", X"16", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"05", X"2f", X"7a", X"5d", X"60", X"67", X"69", X"69", X"66", X"61", X"61", X"62", X"5f", X"61", X"77", X"75", X"67", X"6a", X"72", X"73", X"7c", X"5c", X"04", X"03", X"04", X"03", X"03", X"05", X"57", X"6e", X"6f", X"76", X"7d", X"79", X"75", X"71", X"72", X"6f", X"6e", X"69", X"5e", X"57", X"5a", X"5c", X"5c", X"5a", X"55", X"54", X"50", X"59", X"55", X"32", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"07", X"47", X"81", X"60", X"66", X"6e", X"70", X"6f", X"6d", X"6b", X"69", X"67", X"66", X"69", X"6f", X"6e", X"6d", X"72", X"75", X"7f", X"8f", X"5c", X"04", X"04", X"05", X"03", X"03", X"08", X"63", X"75", X"74", X"77", X"79", X"6e", X"66", X"67", X"6b", X"69", X"68", X"61", X"5c", X"59", X"5a", X"5c", X"5f", X"58", X"53", X"54", X"53", X"58", X"5a", X"4f", X"08", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0d", X"55", X"8c", X"69", X"6a", X"70", X"70", X"76", X"76", X"73", X"72", X"6e", X"6d", X"73", X"75", X"71", X"77", X"7c", X"81", X"87", X"8e", X"58", X"05", X"06", X"0d", X"05", X"05", X"0e", X"68", X"74", X"76", X"7c", X"74", X"6b", X"66", X"66", X"64", X"68", X"6a", X"60", X"5a", X"5a", X"5a", X"5e", X"5f", X"59", X"56", X"59", X"58", X"5c", X"5c", X"5b", X"0e", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"12", X"56", X"98", X"77", X"6d", X"6f", X"74", X"7f", X"7e", X"7b", X"79", X"75", X"74", X"7f", X"79", X"7e", X"83", X"89", X"92", X"91", X"90", X"53", X"08", X"0b", X"1d", X"06", X"07", X"15", X"70", X"77", X"7c", X"80", X"6f", X"6c", X"68", X"65", X"61", X"61", X"6a", X"62", X"5d", X"5c", X"5a", X"5a", X"5c", X"5a", X"5a", X"5d", X"5e", X"5d", X"5f", X"61", X"10", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"13", X"57", X"a6", X"82", X"72", X"76", X"7c", X"86", X"88", X"83", X"82", X"7f", X"7c", X"8e", X"83", X"91", X"97", X"9f", X"a5", X"a0", X"9d", X"56", X"0c", X"16", X"2e", X"0b", X"0a", X"21", X"7c", X"80", X"83", X"83", X"75", X"6f", X"6b", X"67", X"63", X"5f", X"61", X"68", X"5e", X"5c", X"5c", X"5e", X"5f", X"5e", X"5f", X"60", X"60", X"63", X"6b", X"61", X"0c", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"13", X"55", X"af", X"83", X"79", X"7e", X"86", X"8f", X"8f", X"8e", X"8c", X"88", X"88", X"9c", X"96", X"a4", X"a9", X"b1", X"be", X"b5", X"b0", X"55", X"15", X"25", X"40", X"15", X"13", X"30", X"8d", X"8a", X"8b", X"8a", X"7f", X"75", X"6f", X"69", X"62", X"60", X"62", X"65", X"65", X"60", X"5f", X"60", X"65", X"65", X"64", X"67", X"65", X"66", X"77", X"5f", X"0c", X"03", X"03"),
  (X"03", X"02", X"03", X"04", X"03", X"0f", X"4f", X"b2", X"86", X"7e", X"82", X"86", X"91", X"98", X"99", X"96", X"93", X"95", X"a9", X"a6", X"ac", X"b4", X"bd", X"d6", X"d4", X"c5", X"52", X"1f", X"35", X"58", X"22", X"1c", X"45", X"a1", X"9a", X"94", X"94", X"87", X"7d", X"74", X"6b", X"65", X"60", X"61", X"64", X"6a", X"65", X"62", X"66", X"6a", X"6b", X"6c", X"6d", X"6a", X"68", X"83", X"52", X"09", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"04", X"0e", X"45", X"b0", X"8b", X"86", X"8a", X"8a", X"93", X"9d", X"a3", X"a2", X"a0", X"ab", X"b6", X"b4", X"bc", X"c3", X"d2", X"ed", X"f1", X"de", X"60", X"2e", X"4c", X"73", X"38", X"26", X"5c", X"b4", X"ab", X"a4", X"a1", X"94", X"8a", X"7f", X"75", X"6c", X"67", X"66", X"69", X"6f", X"6c", X"6a", X"6d", X"70", X"73", X"73", X"73", X"6f", X"70", X"8b", X"41", X"08", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"0b", X"38", X"a6", X"90", X"8f", X"91", X"92", X"9a", X"a3", X"aa", X"ab", X"b1", X"c3", X"bf", X"be", X"cb", X"d5", X"ed", X"fe", X"fe", X"fa", X"76", X"4b", X"68", X"8a", X"52", X"3b", X"7c", X"c9", X"be", X"b4", X"ab", X"a2", X"98", X"8d", X"82", X"76", X"71", X"6e", X"6f", X"7a", X"75", X"74", X"74", X"76", X"78", X"77", X"72", X"71", X"7c", X"83", X"2a", X"05", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"06", X"27", X"9d", X"95", X"90", X"96", X"98", X"9e", X"a7", X"af", X"b8", X"c1", X"c8", X"c5", X"cb", X"dc", X"ea", X"fc", X"ff", X"ff", X"fe", X"e2", X"af", X"b7", X"b0", X"94", X"7f", X"b5", X"e5", X"d6", X"c8", X"bb", X"b3", X"a8", X"9e", X"93", X"87", X"7e", X"7a", X"7f", X"8d", X"81", X"80", X"83", X"81", X"7d", X"80", X"77", X"6f", X"90", X"6a", X"15", X"04", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"05", X"19", X"8e", X"9a", X"8b", X"94", X"9c", X"a7", X"ac", X"b8", X"c4", X"c8", X"cb", X"d3", X"dc", X"ed", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"fd", X"fd", X"f2", X"de", X"d0", X"c4", X"bc", X"b2", X"a5", X"9b", X"95", X"97", X"99", X"97", X"8d", X"8c", X"8f", X"8a", X"83", X"85", X"80", X"6e", X"92", X"50", X"08", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"14", X"85", X"9b", X"88", X"94", X"9d", X"a9", X"b7", X"c2", X"ca", X"d3", X"da", X"e3", X"ed", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f2", X"e4", X"d4", X"ca", X"c5", X"bd", X"b5", X"af", X"aa", X"a5", X"9e", X"99", X"95", X"94", X"8a", X"82", X"80", X"7e", X"70", X"8c", X"39", X"05", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"14", X"83", X"a3", X"80", X"90", X"9e", X"ad", X"be", X"c5", X"cf", X"dd", X"ea", X"f4", X"fa", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f6", X"e7", X"db", X"d2", X"cb", X"c5", X"bd", X"ba", X"b1", X"aa", X"a3", X"9a", X"96", X"8c", X"7e", X"79", X"75", X"6c", X"83", X"3b", X"04", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"05", X"17", X"78", X"a5", X"71", X"84", X"99", X"aa", X"b6", X"bf", X"d0", X"e2", X"f5", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"f2", X"e7", X"e2", X"dc", X"d4", X"c9", X"bc", X"b8", X"af", X"a8", X"a3", X"96", X"84", X"7a", X"77", X"69", X"79", X"4a", X"05", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"04", X"10", X"61", X"9c", X"74", X"75", X"8c", X"a1", X"b3", X"c0", X"d2", X"e9", X"fa", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f9", X"ef", X"ed", X"e9", X"d8", X"cc", X"bf", X"ad", X"9d", X"96", X"90", X"88", X"81", X"75", X"64", X"70", X"4e", X"08", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"08", X"3e", X"7e", X"80", X"6b", X"7d", X"90", X"a3", X"b9", X"cf", X"ec", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fa", X"fc", X"f2", X"e6", X"d8", X"c6", X"b5", X"a4", X"92", X"84", X"7e", X"7d", X"72", X"61", X"73", X"51", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"06", X"16", X"3e", X"61", X"73", X"74", X"83", X"90", X"a5", X"c1", X"e0", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"ef", X"db", X"c8", X"b8", X"ab", X"9d", X"8c", X"76", X"6f", X"70", X"6e", X"82", X"43", X"09", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"0a", X"22", X"58", X"7c", X"68", X"73", X"82", X"92", X"ab", X"cd", X"ed", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fd", X"fa", X"ec", X"d7", X"c4", X"b7", X"a4", X"91", X"87", X"7c", X"6e", X"70", X"9b", X"77", X"2d", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"05", X"11", X"38", X"72", X"6c", X"72", X"80", X"8c", X"9d", X"b8", X"d8", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f2", X"ea", X"db", X"c4", X"af", X"a7", X"9b", X"90", X"7d", X"72", X"79", X"82", X"96", X"53", X"1c", X"03", X"03", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"07", X"18", X"39", X"68", X"87", X"99", X"b1", X"bb", X"bb", X"d2", X"f7", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ed", X"da", X"c4", X"b0", X"a1", X"99", X"8f", X"82", X"78", X"71", X"9c", X"8c", X"4f", X"23", X"07", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"06", X"16", X"35", X"6f", X"a3", X"cf", X"cf", X"d7", X"de", X"e1", X"f1", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"da", X"c5", X"b3", X"a4", X"96", X"86", X"7c", X"72", X"6b", X"78", X"43", X"1c", X"0b", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"14", X"31", X"5f", X"b2", X"c6", X"9b", X"ac", X"c4", X"df", X"fa", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fe", X"fd", X"fc", X"f5", X"e5", X"ca", X"ad", X"98", X"83", X"76", X"73", X"70", X"5e", X"3d", X"15", X"08", X"04", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"0c", X"1b", X"3d", X"73", X"9c", X"a3", X"b2", X"c4", X"d5", X"e1", X"ef", X"fc", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f8", X"ee", X"e0", X"d7", X"d0", X"c9", X"bc", X"9f", X"83", X"76", X"6b", X"6c", X"52", X"2a", X"0e", X"04", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"04", X"08", X"10", X"25", X"44", X"73", X"9e", X"b4", X"b7", X"c0", X"cf", X"e4", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fe", X"f8", X"ec", X"dc", X"d1", X"bb", X"ab", X"9e", X"92", X"87", X"79", X"73", X"67", X"4e", X"2f", X"16", X"09", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"05", X"0a", X"15", X"21", X"33", X"52", X"97", X"ac", X"ad", X"c5", X"da", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f4", X"d5", X"c6", X"b6", X"ac", X"a2", X"90", X"7e", X"75", X"6f", X"6c", X"69", X"45", X"24", X"14", X"09", X"05", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"06", X"0c", X"11", X"18", X"2e", X"66", X"5e", X"80", X"a5", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f2", X"a9", X"97", X"8b", X"81", X"7a", X"68", X"57", X"4c", X"3e", X"35", X"1b", X"0b", X"07", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"03", X"04", X"07", X"09", X"10", X"16", X"28", X"32", X"79", X"a6", X"e1", X"f2", X"fe", X"fe", X"ff", X"fe", X"de", X"b2", X"79", X"44", X"45", X"3f", X"2e", X"23", X"17", X"0f", X"09", X"09", X"07", X"05", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"07", X"0d", X"10", X"12", X"22", X"2d", X"46", X"5b", X"87", X"87", X"b4", X"ad", X"66", X"39", X"28", X"1e", X"18", X"10", X"0c", X"08", X"07", X"04", X"04", X"05", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"04", X"05", X"06", X"09", X"0d", X"12", X"1a", X"1c", X"23", X"27", X"27", X"27", X"1e", X"14", X"0b", X"09", X"07", X"04", X"04", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"07", X"09", X"0d", X"0c", X"0f", X"0f", X"15", X"11", X"0c", X"0b", X"05", X"04", X"03", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"05", X"05", X"06", X"06", X"06", X"05", X"04", X"05", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
  (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"04", X"04", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"));

  constant imagem_teste3 : MatrizImagem :=  ((X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"04", X"04", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0a", X"1e", X"25", X"27", X"26", X"1e", X"0d", X"0b", X"07", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0b", X"2d", X"38", X"37", X"39", X"3f", X"3f", X"2d", X"2a", X"24", X"17", X"0a", X"16", X"16", X"13", X"0b", X"03", X"03", X"03", X"02", X"03", X"03", X"06", X"09", X"0c", X"16", X"24", X"25", X"1f", X"20", X"1f", X"22", X"1f", X"1f", X"1e", X"15", X"06", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"2b", X"3c", X"3d", X"3e", X"3e", X"40", X"41", X"35", X"37", X"2e", X"2a", X"26", X"29", X"2c", X"29", X"1a", X"03", X"03", X"03", X"02", X"03", X"03", X"18", X"27", X"27", X"2b", X"41", X"61", X"68", X"66", X"62", X"5f", X"5b", X"54", X"4f", X"49", X"35", X"0e", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"1b", X"3c", X"3e", X"41", X"40", X"42", X"46", X"42", X"3e", X"3a", X"34", X"35", X"35", X"33", X"2e", X"2a", X"1b", X"03", X"03", X"03", X"02", X"03", X"03", X"21", X"2d", X"2f", X"31", X"34", X"41", X"5e", X"72", X"78", X"78", X"74", X"6e", X"66", X"5e", X"55", X"3b", X"0a", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0c", X"33", X"3c", X"41", X"44", X"45", X"51", X"52", X"43", X"3f", X"3c", X"36", X"37", X"3b", X"3a", X"32", X"2d", X"19", X"03", X"03", X"03", X"02", X"03", X"03", X"2a", X"31", X"34", X"35", X"39", X"3a", X"3e", X"48", X"54", X"5c", X"66", X"71", X"78", X"77", X"71", X"64", X"36", X"06", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"20", X"3c", X"42", X"43", X"42", X"42", X"47", X"3d", X"35", X"34", X"38", X"39", X"39", X"39", X"3d", X"3b", X"30", X"16", X"03", X"03", X"03", X"02", X"03", X"04", X"32", X"36", X"38", X"3a", X"3d", X"3f", X"42", X"44", X"43", X"44", X"43", X"47", X"50", X"5e", X"6d", X"77", X"60", X"24", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"0b", X"31", X"42", X"44", X"43", X"3f", X"40", X"3d", X"39", X"36", X"36", X"38", X"37", X"3a", X"38", X"38", X"3c", X"38", X"17", X"03", X"03", X"03", X"02", X"03", X"05", X"34", X"3e", X"3f", X"46", X"46", X"4a", X"48", X"49", X"4c", X"4a", X"48", X"44", X"42", X"41", X"43", X"52", X"60", X"4d", X"09", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"1b", X"3d", X"43", X"45", X"40", X"3e", X"3d", X"39", X"38", X"36", X"38", X"38", X"39", X"3a", X"38", X"39", X"34", X"32", X"15", X"03", X"03", X"03", X"02", X"03", X"08", X"37", X"3a", X"3e", X"41", X"44", X"46", X"46", X"4a", X"4b", X"4d", X"4f", X"58", X"47", X"47", X"46", X"51", X"4d", X"48", X"1c", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"2a", X"44", X"42", X"45", X"41", X"3f", X"3c", X"38", X"38", X"37", X"38", X"3a", X"37", X"37", X"35", X"35", X"34", X"32", X"10", X"03", X"03", X"03", X"02", X"03", X"0b", X"3b", X"3c", X"3c", X"3f", X"41", X"44", X"48", X"4e", X"4b", X"49", X"4d", X"5e", X"57", X"51", X"55", X"4f", X"4b", X"48", X"35", X"07", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0c", X"35", X"45", X"41", X"42", X"40", X"3e", X"3a", X"39", X"3a", X"39", X"39", X"3b", X"38", X"38", X"35", X"35", X"36", X"33", X"0f", X"03", X"03", X"03", X"02", X"03", X"10", X"44", X"41", X"45", X"47", X"49", X"4a", X"48", X"4a", X"49", X"4b", X"4b", X"4c", X"4f", X"4b", X"4a", X"4a", X"4a", X"45", X"46", X"16", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"15", X"3f", X"45", X"42", X"44", X"3f", X"3d", X"3b", X"3d", X"3e", X"3c", X"3a", X"3c", X"3a", X"39", X"3a", X"38", X"3a", X"35", X"0e", X"03", X"03", X"03", X"02", X"03", X"14", X"43", X"46", X"4a", X"4d", X"4d", X"4a", X"4a", X"47", X"49", X"4b", X"4b", X"4a", X"4b", X"4c", X"4c", X"4c", X"4a", X"47", X"47", X"2b", X"04", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"06", X"23", X"48", X"45", X"43", X"42", X"40", X"3d", X"3b", X"3e", X"3f", X"40", X"3e", X"3f", X"40", X"40", X"40", X"3c", X"3c", X"36", X"0a", X"03", X"03", X"03", X"02", X"03", X"18", X"44", X"52", X"5b", X"50", X"4c", X"4a", X"4a", X"47", X"49", X"49", X"4b", X"49", X"4b", X"4c", X"4e", X"4f", X"4d", X"49", X"47", X"3a", X"0d", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"09", X"31", X"46", X"46", X"43", X"45", X"44", X"3f", X"40", X"42", X"43", X"40", X"41", X"43", X"43", X"46", X"44", X"41", X"40", X"39", X"08", X"03", X"03", X"03", X"02", X"03", X"1e", X"45", X"4c", X"58", X"51", X"50", X"4a", X"48", X"46", X"47", X"4a", X"4a", X"49", X"49", X"4a", X"4e", X"51", X"51", X"4e", X"4a", X"46", X"1f", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"12", X"3b", X"47", X"47", X"46", X"4a", X"45", X"4b", X"47", X"45", X"43", X"46", X"46", X"49", X"4b", X"4d", X"4a", X"4a", X"4b", X"46", X"08", X"03", X"03", X"03", X"02", X"03", X"24", X"4a", X"4e", X"51", X"52", X"52", X"4e", X"4a", X"4a", X"48", X"49", X"4b", X"48", X"49", X"49", X"4e", X"52", X"57", X"53", X"50", X"4b", X"39", X"04", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"19", X"42", X"48", X"46", X"47", X"49", X"47", X"4d", X"49", X"49", X"48", X"49", X"4b", X"4e", X"50", X"51", X"51", X"54", X"5b", X"49", X"06", X"03", X"03", X"03", X"02", X"03", X"2f", X"52", X"55", X"56", X"54", X"52", X"52", X"51", X"4a", X"47", X"49", X"4b", X"4a", X"49", X"48", X"4e", X"52", X"57", X"59", X"52", X"4f", X"48", X"0f", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"08", X"21", X"50", X"4d", X"4a", X"49", X"4c", X"49", X"47", X"47", X"48", X"49", X"4d", X"4c", X"4c", X"4e", X"51", X"50", X"56", X"55", X"41", X"04", X"03", X"03", X"03", X"02", X"03", X"3c", X"5f", X"5d", X"5a", X"58", X"54", X"57", X"54", X"4d", X"4a", X"4b", X"4c", X"49", X"4c", X"49", X"4c", X"52", X"55", X"57", X"59", X"53", X"4f", X"1e", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"0b", X"31", X"5b", X"5e", X"4e", X"4b", X"4a", X"48", X"48", X"47", X"47", X"47", X"48", X"49", X"4b", X"4d", X"4f", X"52", X"56", X"50", X"3e", X"03", X"03", X"03", X"03", X"02", X"03", X"49", X"6b", X"63", X"5e", X"5c", X"5b", X"5c", X"60", X"50", X"4d", X"4d", X"4b", X"47", X"49", X"49", X"4c", X"51", X"54", X"57", X"56", X"53", X"54", X"30", X"04", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"04", X"0d", X"4d", X"62", X"67", X"5a", X"4f", X"50", X"4f", X"4d", X"4a", X"49", X"4b", X"4b", X"49", X"4c", X"4f", X"54", X"55", X"59", X"56", X"42", X"03", X"03", X"03", X"03", X"02", X"04", X"5e", X"72", X"69", X"66", X"63", X"63", X"62", X"5c", X"53", X"4e", X"50", X"50", X"4e", X"4b", X"4b", X"4d", X"52", X"54", X"56", X"56", X"56", X"54", X"3b", X"08", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"05", X"1c", X"72", X"61", X"66", X"6a", X"5f", X"54", X"57", X"55", X"52", X"52", X"54", X"53", X"4f", X"51", X"52", X"59", X"5b", X"61", X"60", X"45", X"03", X"03", X"03", X"03", X"03", X"06", X"73", X"7a", X"70", X"6d", X"6e", X"73", X"6a", X"5d", X"58", X"57", X"57", X"55", X"53", X"50", X"4e", X"51", X"55", X"57", X"57", X"57", X"5c", X"5c", X"43", X"12", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"06", X"3a", X"81", X"69", X"6d", X"7f", X"62", X"56", X"5a", X"56", X"54", X"54", X"54", X"56", X"52", X"51", X"55", X"5a", X"61", X"64", X"60", X"3f", X"03", X"03", X"03", X"03", X"02", X"09", X"77", X"7f", X"74", X"75", X"76", X"74", X"6b", X"61", X"59", X"58", X"59", X"54", X"52", X"50", X"51", X"54", X"56", X"58", X"56", X"55", X"55", X"58", X"54", X"27", X"04", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"08", X"51", X"83", X"75", X"81", X"7a", X"60", X"5a", X"5c", X"5c", X"59", X"57", X"59", X"57", X"54", X"54", X"5a", X"63", X"74", X"64", X"63", X"3b", X"03", X"03", X"03", X"03", X"02", X"0e", X"79", X"7d", X"75", X"74", X"70", X"70", X"6e", X"6d", X"63", X"5b", X"59", X"56", X"53", X"53", X"53", X"54", X"58", X"57", X"56", X"55", X"55", X"54", X"65", X"48", X"07", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"0f", X"5e", X"8e", X"90", X"86", X"61", X"5f", X"5e", X"5d", X"5c", X"5d", X"5c", X"5d", X"5a", X"5a", X"5c", X"64", X"66", X"6d", X"66", X"6a", X"3a", X"03", X"03", X"03", X"03", X"03", X"16", X"83", X"70", X"70", X"74", X"73", X"76", X"74", X"76", X"70", X"62", X"5b", X"5a", X"53", X"54", X"54", X"57", X"58", X"5a", X"58", X"56", X"58", X"55", X"63", X"58", X"0c", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"13", X"62", X"92", X"79", X"6a", X"61", X"61", X"61", X"5d", X"5c", X"5e", X"5f", X"61", X"5d", X"64", X"6f", X"70", X"6a", X"70", X"68", X"6e", X"35", X"03", X"03", X"03", X"03", X"03", X"1e", X"80", X"73", X"75", X"79", X"77", X"78", X"79", X"78", X"75", X"6e", X"5e", X"5a", X"57", X"57", X"56", X"54", X"56", X"59", X"59", X"59", X"59", X"55", X"62", X"5b", X"0e", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"13", X"61", X"90", X"79", X"6e", X"63", X"61", X"61", X"62", X"5e", X"60", X"63", X"62", X"61", X"70", X"76", X"6e", X"6f", X"76", X"73", X"76", X"32", X"03", X"03", X"03", X"03", X"04", X"2a", X"89", X"7f", X"7e", X"7e", X"7f", X"7b", X"7a", X"7c", X"7a", X"75", X"64", X"5d", X"59", X"58", X"59", X"56", X"57", X"58", X"5a", X"59", X"58", X"5d", X"69", X"53", X"0b", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"12", X"58", X"95", X"7c", X"6d", X"63", X"63", X"66", X"65", X"66", X"65", X"66", X"67", X"68", X"76", X"7d", X"76", X"78", X"7b", X"83", X"81", X"2b", X"03", X"04", X"03", X"03", X"06", X"39", X"94", X"8a", X"88", X"87", X"86", X"7f", X"7d", X"7f", X"7b", X"78", X"6c", X"60", X"5d", X"5c", X"5a", X"59", X"5b", X"59", X"59", X"5a", X"5b", X"62", X"6d", X"4f", X"0b", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"0d", X"4b", X"92", X"73", X"6b", X"62", X"5f", X"64", X"67", X"68", X"68", X"6a", X"6c", X"74", X"77", X"7f", X"85", X"81", X"89", X"8b", X"88", X"26", X"03", X"03", X"03", X"03", X"08", X"4f", X"a3", X"98", X"92", X"91", X"89", X"84", X"80", X"7f", X"7e", X"77", X"6f", X"63", X"62", X"61", X"5d", X"5f", X"5f", X"5e", X"5d", X"5a", X"5f", X"64", X"6e", X"45", X"08", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"0c", X"3e", X"8f", X"78", X"66", X"65", X"5b", X"5f", X"64", X"68", X"6b", X"6e", X"75", X"7c", X"7e", X"84", X"91", X"91", X"96", X"9d", X"aa", X"27", X"04", X"04", X"03", X"04", X"0b", X"62", X"b4", X"a4", X"9e", X"99", X"90", X"8b", X"85", X"84", X"82", X"7c", X"77", X"68", X"65", X"64", X"62", X"65", X"66", X"65", X"63", X"62", X"69", X"6f", X"71", X"38", X"06", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"08", X"30", X"80", X"a2", X"64", X"67", X"61", X"5e", X"63", X"66", X"6a", X"74", X"7d", X"81", X"84", X"90", X"9b", X"a3", X"a5", X"af", X"c1", X"1d", X"07", X"06", X"05", X"06", X"11", X"6d", X"b6", X"af", X"a5", X"9e", X"97", X"91", X"8b", X"8a", X"87", X"84", X"7f", X"71", X"69", X"68", X"67", X"66", X"69", X"6a", X"69", X"69", X"72", X"87", X"6c", X"25", X"04", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"04", X"1e", X"6f", X"a5", X"6f", X"61", X"64", X"69", X"6c", X"6c", X"73", X"77", X"7d", X"86", X"8e", X"9f", X"a7", X"ab", X"b0", X"cd", X"aa", X"27", X"10", X"0c", X"0b", X"0e", X"1e", X"7b", X"bb", X"b3", X"af", X"a8", X"a2", X"9b", X"95", X"94", X"91", X"8e", X"88", X"7a", X"72", X"6f", X"6b", X"6b", X"6b", X"6b", X"70", X"76", X"7a", X"9a", X"5b", X"11", X"04", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"11", X"5f", X"9c", X"72", X"63", X"65", X"6c", X"74", X"78", X"73", X"78", X"86", X"93", X"9f", X"ad", X"b5", X"b7", X"b5", X"dd", X"d7", X"4c", X"2a", X"20", X"1e", X"26", X"3a", X"99", X"c7", X"bb", X"b6", X"b2", X"b1", X"ae", X"a7", X"a0", X"9e", X"9a", X"94", X"88", X"7e", X"79", X"71", X"70", X"71", X"71", X"7a", X"81", X"80", X"9b", X"47", X"07", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"0c", X"58", X"87", X"62", X"66", X"6d", X"72", X"78", X"89", X"78", X"83", X"91", X"9f", X"a9", X"b6", X"bf", X"bf", X"ba", X"dd", X"fb", X"98", X"5a", X"49", X"46", X"52", X"7f", X"e2", X"d6", X"cb", X"c4", X"c3", X"c1", X"bf", X"b8", X"b2", X"af", X"a9", X"a4", X"99", X"8f", X"89", X"80", X"7e", X"7c", X"80", X"86", X"8c", X"86", X"97", X"34", X"05", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"0c", X"56", X"67", X"58", X"62", X"6a", X"74", X"81", X"8e", X"8c", X"8d", X"97", X"a0", X"ab", X"b9", X"c6", X"c4", X"bd", X"d1", X"ff", X"f4", X"dc", X"be", X"c1", X"d9", X"f5", X"fe", X"f5", X"ed", X"e6", X"e1", X"dc", X"d6", X"ce", X"c5", X"bb", X"b0", X"aa", X"a1", X"99", X"92", X"87", X"84", X"86", X"87", X"8c", X"8b", X"88", X"98", X"3a", X"03", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"0e", X"4d", X"6b", X"6f", X"5f", X"69", X"73", X"7f", X"8e", X"9b", X"99", X"a0", X"a9", X"b3", X"c3", X"d0", X"d0", X"c9", X"d5", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fd", X"fb", X"ee", X"dc", X"cf", X"c1", X"b6", X"ab", X"a1", X"9d", X"8d", X"82", X"7b", X"7b", X"81", X"84", X"86", X"84", X"99", X"4f", X"04", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"09", X"47", X"7a", X"7c", X"69", X"75", X"73", X"7d", X"90", X"a5", X"b0", X"b7", X"bd", X"c6", X"d6", X"e0", X"e7", X"ee", X"f6", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"ea", X"d9", X"c8", X"ba", X"b0", X"aa", X"a5", X"a1", X"8e", X"7d", X"74", X"76", X"78", X"7a", X"7a", X"92", X"56", X"07", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"05", X"2d", X"5f", X"73", X"69", X"85", X"8f", X"8b", X"99", X"ab", X"be", X"cd", X"d7", X"de", X"ec", X"f9", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f9", X"e8", X"d3", X"bd", X"af", X"a5", X"9f", X"a0", X"9a", X"8c", X"80", X"78", X"6f", X"6f", X"73", X"91", X"58", X"07", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"04", X"0f", X"3a", X"62", X"77", X"7a", X"9f", X"aa", X"b0", X"bb", X"c9", X"da", X"ed", X"f7", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"e5", X"d0", X"bc", X"ad", X"a4", X"9c", X"94", X"91", X"8b", X"82", X"78", X"6c", X"6c", X"90", X"46", X"07", X"03", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"06", X"1d", X"41", X"65", X"71", X"80", X"9e", X"b3", X"c6", X"df", X"f3", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"e2", X"c8", X"b6", X"aa", X"a4", X"98", X"8f", X"88", X"7f", X"75", X"6f", X"7a", X"7d", X"32", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"0b", X"20", X"49", X"77", X"84", X"8f", X"a0", X"bb", X"dc", X"f8", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"f1", X"db", X"c3", X"ab", X"9d", X"93", X"8f", X"85", X"79", X"6a", X"66", X"81", X"57", X"1c", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"07", X"12", X"29", X"5f", X"8d", X"93", X"a4", X"bd", X"d4", X"e3", X"ee", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f3", X"dd", X"df", X"d7", X"c6", X"aa", X"8e", X"7f", X"77", X"72", X"6a", X"62", X"6d", X"4b", X"24", X"06", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"0e", X"1c", X"58", X"a2", X"98", X"a8", X"be", X"db", X"f5", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f9", X"d6", X"be", X"b4", X"a9", X"9c", X"87", X"73", X"66", X"5c", X"63", X"68", X"4c", X"1c", X"07", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"0e", X"1d", X"54", X"99", X"a4", X"c1", X"ee", X"fe", X"fc", X"fe", X"ff", X"ff", X"ff", X"fe", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"ff", X"fa", X"ee", X"d9", X"c0", X"a8", X"96", X"8d", X"85", X"79", X"6c", X"6e", X"5b", X"28", X"21", X"07", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"13", X"14", X"16", X"5d", X"9c", X"bb", X"d0", X"d4", X"cf", X"df", X"e8", X"e4", X"ec", X"e6", X"eb", X"ef", X"e6", X"e8", X"f1", X"f9", X"f4", X"f6", X"fb", X"ff", X"fd", X"fc", X"fc", X"f8", X"ec", X"df", X"cd", X"bc", X"b0", X"a0", X"96", X"8f", X"96", X"97", X"5a", X"1f", X"0f", X"05", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"04", X"05", X"0d", X"2f", X"60", X"8d", X"9f", X"a8", X"a0", X"7a", X"74", X"87", X"8c", X"97", X"a7", X"a5", X"ae", X"b3", X"cd", X"f8", X"f8", X"e3", X"f1", X"ec", X"e4", X"e3", X"e2", X"da", X"d3", X"c9", X"b8", X"b2", X"ab", X"a0", X"a0", X"7e", X"48", X"24", X"07", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"06", X"0a", X"16", X"31", X"4f", X"48", X"5f", X"6d", X"78", X"7e", X"89", X"8e", X"8b", X"84", X"8e", X"89", X"98", X"d1", X"bb", X"b5", X"be", X"bc", X"b5", X"ac", X"ad", X"ab", X"ad", X"b6", X"c8", X"a0", X"5d", X"39", X"1d", X"0c", X"06", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"04", X"04", X"05", X"08", X"0e", X"24", X"45", X"4a", X"78", X"83", X"79", X"7b", X"7d", X"84", X"88", X"70", X"5e", X"70", X"7b", X"8a", X"93", X"90", X"7e", X"6b", X"68", X"6d", X"52", X"30", X"17", X"0b", X"07", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"05", X"0c", X"10", X"26", X"42", X"5f", X"6c", X"5d", X"5d", X"47", X"48", X"3d", X"38", X"3d", X"43", X"46", X"3f", X"2c", X"22", X"15", X"0d", X"08", X"07", X"05", X"05", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"04", X"03", X"03", X"07", X"07", X"18", X"26", X"19", X"15", X"22", X"1a", X"0b", X"09", X"08", X"0a", X"09", X"05", X"05", X"04", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"04", X"03", X"04", X"04", X"04", X"04", X"04", X"03", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"04", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"),
 (X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"02", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"03", X"02", X"03", X"03"));

-- signals                                                   
SIGNAL ENDSIM : STD_LOGIC := '0';
SIGNAL clk_count : natural := 0;
SIGNAL brilho_maximo : UNSIGNED(24 DOWNTO 0);
SIGNAL threshold1    : std_logic_vector(7 downto 0);
SIGNAL meioVert      : unsigned(7 downto 0);
SIGNAL meioImagem    : unsigned(7 downto 0);
SIGNAL in_clock : STD_LOGIC;
SIGNAL in_janela : STD_LOGIC;
SIGNAL RX : STD_LOGIC_VECTOR(3 DOWNTO 0) := (others => '0');
SIGNAL pixel_entrada : STD_LOGIC_VECTOR(7 DOWNTO 0) := (others => '0');
SIGNAL bloco_atual : natural range qtd_imagens downto 0 := 0;
SIGNAL linha : integer range 0 to numcols - 1 := 0;
SIGNAL coluna : integer range 0 to numlin - 1 := 0;
SIGNAL reset : STD_LOGIC;
SIGNAL start_stop :  STD_LOGIC;
SIGNAL contador12b : STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL qtd_imagens : UNSIGNED(1 DOWNTO 0) := "11";
--SIGNAL fim_imagem : STD_LOGIC := '0';
SIGNAL frequencia_camera : real := 85.000E6;


COMPONENT ProcessadorImagemGMAW
	PORT (
	in_clock      : in std_logic;                                       -- clock gerado pela camera
  FVAL_teste    : in std_logic;                                       -- para simulacao
  RX            : in std_logic_vector(3 downto 0);                    -- canais de dados
  brilho_maximo : in unsigned(24 downto 0) := to_unsigned(720000,25);
  threshold1    : in std_logic_vector(7 downto 0);
  meioVert      : in unsigned(7 downto 0);
  meioImagem    : in unsigned(7 downto 0);
  pixel_entrada : in std_logic_vector(7 downto 0) := "00000000";      -- para simulacao
  limEsqPoca    : out natural range numcols downto 0;
  limDirPoca    : out natural range numcols downto 0);	
END COMPONENT;


-- Procedure for clock generation
  procedure clk_gen(signal clk : out std_logic; constant FREQ : real) is
    constant PERIOD    : time := 1 sec / FREQ;        -- Full period
    constant HIGH_TIME : time := PERIOD / 2;          -- High time
    constant LOW_TIME  : time := PERIOD - HIGH_TIME;  -- Low time; always >= HIGH_TIME
  begin
    -- Check the arguments
    assert (HIGH_TIME /= 0 fs) report "clk_plain: High time is zero; time resolution to large for frequency" severity FAILURE;
    -- Generate a clock cycle
    loop
      if (ENDSIM = '0') then
        clk <= '1';
        wait for HIGH_TIME;
        clk <= '0';
        wait for LOW_TIME;
      else
        wait;
      end if;
    end loop;
  end procedure;



BEGIN
  -- Clock generation with concurrent procedure call
  clk_gen(in_clock, frequencia_camera);  -- 166.667 MHz clock

  -- Time resolution show
  assert FALSE report "Time resolution: " & time'image(time'succ(0 fs)) severity NOTE;



	i1 : ProcessadorImagemGMAW
	PORT MAP (
-- list connections between master ports and signals
	brilho_maximo => brilho_maximo,
  threshold1 => threshold1,
  meioVert => meioVert,
  meioImagem => meioImagem,
  in_clock => in_clock,
	RX => RX,
	FVAL_teste => in_janela,
	pixel_entrada => pixel_entrada
	);

brilho_maximo <= to_unsigned(720000,25) after 0 ns;
threshold1    <= "00001010" after 0 ns;
meioVert      <= to_unsigned(30,8) after 0 ns;
meioImagem    <= to_unsigned(31,8) after 0 ns;

in_janela <= '1' after 0 ns,
             '0' after 5 ns,
             '1' after (1 sec / frequencia_camera) * (numcols * numlin)- 1 ns,
             '0' after (1 sec / frequencia_camera) * (numcols * numlin + 1) - 1 ns,
             '1' after (1 sec / frequencia_camera) * 2 * (numcols * numlin) - 1 ns,
             '0' after (1 sec / frequencia_camera) * (2 *(numcols * numlin) + 1) - 1 ns,
             '1' after (1 sec / frequencia_camera) * 3 * (numcols * numlin) - 1 ns,
             '0' after (1 sec / frequencia_camera) * (3 *(numcols * numlin) + 1) - 1 ns;

IN_process: process (in_clock) begin
  if(rising_edge(in_clock)) then
    clk_count <= clk_count + 1;

    -- avanca as imagens
    case bloco_atual is
      when 0 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste0(linha, coluna));
      when 1 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste1(linha, coluna));
      when 2 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste2(linha, coluna));
      when 3 => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste3(linha, coluna));
      when others => pixel_entrada <= STD_LOGIC_VECTOR(imagem_teste0(linha, coluna));
    end case;

    -- marcacao de linhas, colunas e parada na simulacao
    if (coluna = numcols - 1) then
      coluna <= 0;
      if (linha = numlin -1) then
        linha <= 0;
        --fim_imagem <= '1';
        bloco_atual <= bloco_atual + 1;
      else
        linha <= linha + 1;
      end if;    
    else
      coluna <= coluna + 1;
    end if;

    if (clk_count = 4 * (numlin * numcols)) then
      ENDSIM <= '1';
    end if;
  end if;
  

--when -label end_of_simulation {end_of_sim == '1'} {echo "End of simulation" ; stop ;}
end process;


END ProcessadorImagemGMAW_arch;