 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 04 06 05 0a 04 06 05 03 09 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 05 0a 02 06 0f 11 08 0d 08 05 0d 0d 17 12 11 0d 06 0a 05 09 05 08 06 06 09 0c 0b 0b 05 08 00 06 0f 04 09 07 05 03 04 06 07 04 08 06 06 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 03 06 06 03 00 06 05 03 04 06 05 03 01 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 02 06 05 0b 00 0e 08 0c 0d 11 18 12 17 11 15 16 19 16 15 18 14 13 0a 15 09 12 0f 0c 13 0b 14 16 15 13 10 10 0f 08 0b 04 0a 0a 05 03 07 06 05 03 00 06 05 04 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 05 07 09 0a 05 0b 19 10 05 05 02 13 1b 11 13 1a 14 17 15 1a 24 1e 23 21 12 0c 22 1e 24 1f 1f 13 13 1b 1a 1f 24 15 0d 09 0b 08 14 13 09 03 04 06 05 03 08 0a 0c 15 0b 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 15 10 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 07 06 08 03 00 08 05 0a 03 0a 05 06 11 11 08 0d 13 15 18 17 17 18 12 17 16 1e 25 28 27 23 18 1e 2f 2b 31 29 38 28 23 2a 27 29 27 13 0f 11 0e 0e 20 1f 19 12 0e 06 08 06 12 13 19 08 0e 0f 0a 05 04 0d 07 03 0a 06 05 03 02 08 05 03 04 06 08 17 0a 06 05 03 02 06 05 03 00 06 05 03 07 06 05 03 09 07 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 12 0b 07 0b 06 0d 0a 08 0a 06 0d 0e 12 16 1c 22 26 31 40 31 29 21 10 1c 1b 2b 2e 3b 33 2a 2c 30 41 3e 42 4a 3b 30 31 38 3e 36 2e 20 20 17 17 14 17 24 23 1e 14 13 1b 10 17 12 14 13 10 13 19 0b 0e 09 08 0a 11 14 0a 03 07 07 07 07 05 06 05 03 0f 0d 06 0b 00 06 05 03 00 07 05 07 02 06 07 04 0a 08 0c 03 04 06 05 0a 00 06 06 0b 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 08 05 03 0a 10 0a 0c 0f 0e 0c 0f 0f 0b 12 11 1f 25 22 2e 2a 34 39 4f 45 2f 25 28 2f 2e 3e 3f 3e 35 3b 3a 49 52 47 51 59 3c 3c 35 3c 40 2a 2f 26 2c 27 1d 29 27 34 22 2b 23 22 17 1e 1d 0f 1a 1c 14 12 19 10 0f 1a 16 1a 0b 0b 12 0f 13 12 07 0b 06 05 0d 0c 10 05 03 07 06 05 03 09 0a 05 0c 0e 06 06 03 04 12 0a 05 02 06 05 03 01 09 05 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0a 06 04 03 06 05 03 0f 14 0c 0b 12 13 0b 10 14 10 15 12 18 21 24 29 39 2a 28 27 2b 2f 3a 40 3f 38 37 33 3b 3c 43 41 49 40 42 41 45 43 48 4a 48 49 3e 3a 47 4c 41 3a 41 3b 36 30 36 3f 38 32 36 2f 2a 2a 2e 37 27 2c 27 28 24 1f 2b 22 22 22 23 24 23 24 1f 16 1b 16 16 0e 17 1a 11 1a 1a 0d 14 0e 0b 08 0b 0c 10 07 0b 07 0a 06 06 08 09 0a 0c 06 05 09 0f 06 05 09 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 03 06 07 04 00 06 0b 0f 0b 0a 06 0b 0f 06 0d 14 15 0d 14 07 14 1c 11 20 18 1a 18 18 21 2f 31 2b 3b 32 31 33 2f 35 2f 3c 44 3d 43 3b 46 4a 51 58 54 50 47 4f 54 59 55 4b 49 4e 48 41 46 4e 48 4c 57 54 51 42 3f 44 3d 48 41 3d 41 35 35 33 35 32 2f 36 32 2f 2b 26 2e 32 2c 31 2b 2c 25 26 25 22 1e 1b 1e 23 29 27 25 20 24 21 17 10 20 0f 0e 1a 0d 15 0f 0a 05 0b 07 0f 12 09 0b 0d 03 06 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 10 0f 0d 13 0a 0a 0e 08 0f 0d 10 16 1b 11 16 21 25 22 24 24 27 33 2d 38 3a 3e 3d 45 40 36 3e 3e 3a 3d 3b 4b 47 4c 4f 4a 57 53 55 54 60 5d 5b 56 51 51 5a 55 57 55 50 53 55 57 53 58 56 52 4f 54 50 44 4e 43 49 33 45 3f 36 37 3b 3a 3a 30 33 35 3c 3b 39 3b 32 2e 2f 2c 37 31 33 35 34 31 34 3d 39 33 2e 2c 2f 22 22 25 15 1e 1f 1e 22 18 16 0d 16 0d 0d 06 09 04 06 06 0e 03 06 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 0c 06 05 0b 0b 0c 0f 06 16 24 14 1a 11 17 15 18 12 11 1d 21 25 22 2c 2b 2f 35 3b 42 41 49 3c 39 41 44 44 4e 46 4b 4a 4b 58 54 4b 4c 4f 52 51 57 58 54 5d 5d 63 59 5e 60 62 65 68 62 63 6d 6a 66 69 61 6a 67 67 71 63 65 5d 60 62 5b 58 54 55 4e 4e 49 4b 4b 4c 4c 46 3e 3e 43 45 44 4c 4a 44 38 34 2e 35 34 38 32 36 33 35 3f 3b 3d 3c 3b 35 34 2f 32 34 2a 27 2e 30 2a 23 20 1d 24 20 17 14 14 11 11 05 0d 0a 06 0d 03 02 08 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0a 0c 05 11 05 06 0a 05 02 09 13 0e 0e 16 12 1b 25 25 1c 10 17 17 17 1e 20 1e 2b 30 35 3a 39 32 31 4e 46 48 4f 4b 45 4b 52 5f 63 63 54 57 5b 55 53 5d 59 51 58 57 5a 60 61 66 68 66 67 6a 69 69 72 6d 6a 6f 6f 72 71 70 71 78 73 6f 6f 7b 72 63 6d 66 6b 61 67 64 59 56 5a 56 55 55 5d 51 54 57 50 4f 5b 60 5a 56 55 4a 4f 3d 4f 47 4b 4d 4b 49 51 57 53 48 47 4b 42 4a 4c 47 44 3c 41 3b 44 36 31 27 2b 27 2f 31 28 1d 1a 16 20 12 0d 09 05 07 00 07 07 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 10 03 0e 0c 16 12 06 05 08 08 0c 14 10 11 0f 16 11 1c 22 20 20 2a 2a 25 32 30 31 39 40 38 41 3e 36 46 54 56 60 5b 5a 53 59 63 6a 71 67 65 60 5e 5b 5f 68 5a 5a 64 64 64 5c 69 5d 75 71 6e 68 6e 6a 6b 70 6a 6e 77 73 78 75 78 78 6a 73 70 6f 78 69 70 6a 76 6a 6c 64 64 57 5e 61 5b 5e 5c 55 55 4c 56 4e 59 5e 59 60 5f 5b 61 61 6b 6b 65 69 6a 6a 71 6d 7e 7b 77 82 7c 7b 7b 6f 69 60 57 6a 5e 55 54 54 3e 3b 36 35 39 30 3e 34 37 28 1e 11 0b 0b 07 06 09 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 13 17 08 12 13 18 1c 20 18 09 14 0c 11 16 1c 20 1f 22 25 25 29 2e 26 30 32 41 3a 35 3b 3d 4e 51 45 46 49 4d 5a 61 60 6a 70 6b 64 5c 6d 73 7a 73 69 6c 5e 61 66 6d 66 5f 60 65 63 66 6f 71 75 76 76 75 6e 6b 6d 6e 6a 74 77 78 80 75 74 80 7a 79 7b 82 75 77 77 73 6a 69 67 6a 66 5b 62 6d 62 5d 5f 59 5a 59 52 61 63 67 6e 5d 64 63 65 71 70 7b 73 6d 80 8a 8a 8e 92 9b 9e a4 a7 9f 93 8e 73 74 81 96 9e 92 94 8b 7c 6a 54 4e 4c 4d 5c 56 55 54 3a 34 32 1c 16 0d 0c 11 09 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 10 0d 1a 1a 1a 14 14 21 20 24 25 1d 1b 19 19 14 1e 1e 2d 34 2a 30 35 33 3c 37 3d 49 4b 52 4e 54 59 5e 5a 6a 6d 66 64 62 64 69 6e 6c 6b 75 6e 6c 70 75 75 71 6f 6e 6b 71 77 7a 6f 6d 68 6e 6f 6e 7b 78 78 79 78 7d 77 7a 7b 76 7c 7a 7f 81 83 7b 81 82 83 7d 81 84 7b 73 7e 77 78 73 6f 6b 71 66 73 70 70 66 68 61 5d 58 59 5f 6a 6e 67 6b 6f 6e 73 71 7a 72 7a 82 89 96 9b a8 ad af b7 bb af a4 90 8a 88 86 8c b1 c3 c4 c1 ba bf a6 9b 8a 86 80 7a 81 81 6f 64 59 41 28 24 1e 0d 13 11 06 05 03 02 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 05 06 0b 0f 0b 1f 1e 24 2d 32 28 27 2a 2e 2f 2a 1d 26 1c 27 28 2a 29 3a 3d 43 45 4c 5e 52 60 5a 5e 61 64 60 67 67 73 76 6e 70 6c 69 70 76 74 6f 72 7b 6f 71 71 75 75 66 62 79 6b 79 7a 78 75 72 73 73 72 76 7d 7b 7e 7a 81 7b 84 79 70 7b 84 7f 8b 7f 88 84 82 83 86 7f 86 84 84 7e 7d 74 7a 7b 75 67 73 70 70 77 71 67 6a 5d 57 57 5d 60 68 70 68 64 6d 72 6f 73 72 72 7b 87 94 9a a0 b5 b3 ae b5 b5 ab 9e 94 83 89 8a 9d b7 c9 d3 dc e8 e4 de e0 cf c5 ba b6 a6 a5 96 81 6d 55 39 33 33 25 26 1e 15 05 06 09 06 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 14 1c 1c 1c 24 36 3c 37 40 35 38 31 27 2e 2c 2c 33 33 3e 4a 4c 57 5e 62 6a 6b 63 62 60 6e 65 68 7c 7a 72 7b 80 80 6e 76 77 71 7e 7a 74 73 73 70 67 65 6d 6d 72 6b 6d 6d 6e 75 79 7a 84 82 80 77 7f 88 8d 87 84 83 87 83 7b 81 84 81 89 8c 94 8e 8e 8d 8b 85 8a 86 89 86 85 7c 83 7d 80 75 76 77 75 7a 7a 73 69 6a 5f 5f 63 65 60 61 70 6f 71 74 71 6d 6f 76 75 78 76 7e 8c a0 9e a6 aa a9 a9 a7 9f 9b 8f 88 93 a4 b3 c2 c4 c8 d4 ed f4 fb f9 f8 ed de cc bd b3 a3 90 7e 66 4d 47 3d 3c 33 34 2d 16 0d 03 06 11 0a 0b 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 08 06 0e 0b 0d 1d 1c 25 31 38 3c 48 47 3d 37 3d 33 3a 3d 4e 55 62 61 6b 6c 73 75 79 75 6e 6e 6a 70 72 71 77 84 85 81 82 84 86 7e 7d 7a 76 72 79 75 6e 74 75 79 71 6d 6c 68 6e 6b 6f 6c 72 70 76 7c 77 84 84 81 8f 96 99 96 85 90 84 85 81 81 8c 92 99 9a a0 94 8e 9c 95 8e 87 80 87 88 88 84 86 82 7c 80 81 75 7d 82 79 71 73 71 67 6b 62 61 6d 79 82 79 76 72 6c 74 76 83 83 84 82 85 9c 9a 9d a2 ae ad a5 94 9c 99 9e ad c4 d4 cc c1 b5 c5 dd e8 f0 f4 f6 ea d9 be af a8 9f 89 7b 6b 61 64 56 57 4d 49 44 37 23 20 0e 15 07 0f 0e 06 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 0e 0c 0d 13 12 13 15 2a 27 3a 3e 42 49 47 46 4b 4d 47 59 56 62 6a 76 6f 7c 77 74 73 7a 7a 75 77 71 7b 7d 7d 80 91 7c 81 7e 7b 80 74 74 75 6c 71 72 6d 6b 67 70 6f 74 72 74 74 6d 6d 6b 73 69 73 79 7a 7c 83 89 89 8b 90 9b 98 90 95 8e 92 88 91 8c 98 9c aa a6 a2 9c 9a 92 92 90 96 90 93 8d 87 81 8d 8c 82 76 81 7e 7d 80 6e 6d 74 74 71 6e 6f 77 80 87 7b 77 6d 6d 75 7f 83 87 89 87 92 91 9a 9f a8 aa a4 a2 a5 a8 a9 b7 cd e1 dd cf c5 b7 bd c7 cf dc d8 d9 cc c9 b0 a6 9c 8f 7a 71 72 78 81 7c 6e 60 50 4a 4a 38 38 21 23 15 16 15 14 05 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 0f 0c 16 1c 15 20 23 22 34 37 41 46 4c 4d 4d 4d 53 5a 67 68 77 79 7e 85 80 76 71 74 71 77 72 79 75 73 78 7c 79 75 6a 69 7e 7b 75 7d 74 6f 73 70 6f 68 77 74 76 7c 74 80 7c 75 70 75 77 71 78 6f 83 7e 75 70 7e 79 84 8d 96 9c a4 a5 9e 9e 92 96 96 a0 a2 a5 a7 aa a6 a2 9e 94 92 93 93 96 90 8f 93 91 90 89 85 87 83 7b 7b 71 7d 76 6a 6f 69 7a 7c 7f 89 87 7e 7e 81 84 86 8e 8a 8f 98 93 9a 95 a0 a4 a5 a7 a5 b4 b2 be d4 ee fb db cd c5 ba bd c1 c0 c5 c6 c1 bb b3 ad 9c 94 80 7a 7e 79 78 7f 69 6b 62 5a 5a 53 55 4d 39 31 37 31 1f 1e 11 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 05 08 07 0d 19 1a 1c 1f 2d 2a 2b 30 35 32 43 40 46 4a 44 48 4e 55 65 66 6f 75 7c 75 73 78 72 7a 75 79 7a 74 76 7b 76 77 7c 7c 81 7c 82 7d 86 86 84 80 83 72 74 78 82 79 81 80 86 7e 81 81 72 83 78 7b 80 7c 7f 85 7d 7f 79 77 76 7b 85 87 94 a9 9e a5 9f a3 99 95 9e a1 9c a2 ab a6 a4 9a a3 a0 a4 9b 98 99 8e 9c 91 99 98 91 8b 8d 82 7e 80 7c 84 75 7e 7b 86 89 86 8e 90 85 91 92 99 96 94 8b 92 99 99 9e a8 9f 9f a9 ac b5 c0 ca da ed f8 ec e0 c9 c2 cb cc c4 b3 b8 bd c3 b6 a5 a3 95 96 7f 80 85 83 7b 79 74 6b 68 63 5d 60 5e 5e 58 4d 4a 47 3a 2d 1f 17 10 07 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 0e 0f 13 0c 1a 1d 24 2e 35 39 37 36 38 3a 3c 44 48 49 5e 65 54 5f 5e 64 6b 67 68 6f 6c 70 76 74 7e 7e 81 7d 78 7f 7a 76 7d 75 7f 89 80 82 87 7f 8d 8c 85 84 8a 89 86 84 88 93 95 98 90 91 85 8d 80 84 89 7d 85 80 86 8d 84 7e 85 7b 7d 7d 86 8e 9e a7 a4 a0 a0 a0 9f 97 9e 9d 99 a3 a3 a3 a6 a6 af ad a5 a6 9b 9e 9a 9b 92 96 90 91 83 85 82 8c 8d 87 8e 93 8b 87 8e 8c 96 9c 93 97 9a 95 8f 91 8d 9c a2 a7 a3 a1 aa ab ad b9 bf ca d6 f2 f9 fc f3 d5 de da d5 d8 d6 cf c9 c4 bc bd b5 af 9c a0 97 95 92 88 7d 7e 82 77 73 71 6e 69 73 66 61 58 4d 48 44 42 33 31 1b 0c 11 0d 09 07 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0a 06 09 0e 1e 1e 22 28 20 2e 38 3b 32 37 31 3c 41 3e 4a 59 5a 5c 74 78 61 5f 60 5f 63 68 68 73 7a 7b 7f 88 89 84 8b 85 8d 83 7c 87 75 87 89 8e 8c 89 94 85 8c 8f 8c 89 8f 94 97 8e a0 9f a5 a1 9d 9b 96 95 8d 91 8b 8f 8b 8d 91 78 89 83 87 87 80 8b 8b 94 9f 9f 9d 9b 99 98 96 95 9e 95 95 99 a4 a2 a9 ac ad a5 a7 9d a0 9f 9f 9f 99 9b 96 85 8a 8e 8b 92 91 98 9b 91 94 91 8c 92 9b 9b 8f 94 89 8a 89 9c 9e a3 9c a7 a7 a6 ad b6 bf c6 da f8 ff f9 fd f1 e9 e9 e7 e3 e9 e9 e4 e5 db d3 c8 c1 ba ad 9c a1 9a 90 8c 84 85 7f 7f 84 89 7f 78 7b 7b 75 5f 52 52 4b 41 41 48 32 29 20 19 08 0c 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 0f 07 0d 13 0a 22 34 2f 28 2b 39 38 3e 45 32 39 39 47 52 5a 52 56 59 5e 5f 69 6a 5f 60 5f 63 6c 75 72 7b 85 8c 92 9d 96 94 91 94 8e 8d 8c 8d 8c 8d 89 94 96 95 9a 94 93 95 92 9e 9d 9f a8 a9 b2 b5 b3 b2 b1 ad ac a4 95 97 9b 97 92 98 8b 8d 8b 83 8e 96 8b 94 9d 9e 9f 9a 9b 99 94 99 9b 91 90 9b 93 9e a2 9c af b5 b8 a9 9e a1 a3 a4 a1 8b 99 98 97 a0 a4 9c ac a3 9d 98 9b 96 96 8f 95 a0 94 9d 94 9c 96 95 91 9b a1 a0 a9 a8 b3 bc bc c2 d2 f3 ff ff fc ff ff ff ff fd ff ff ff ff fe ec dc cd d2 c3 b9 b3 a4 9e 9a 94 8f 90 8a 8b 8a 91 8b 88 81 80 6e 70 60 60 4e 56 44 49 48 45 41 34 22 17 10 0a 06 07 07 01 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0a 17 19 16 22 2e
 31 31 31 32 36 36 39 34 41 47 43 4d 4c 5d 4a 57 5e 5d 5f 5e 64 68 5f 69 74 6e 74 84 85 8f 8d 9e 9f 9e a3 a2 a0 a0 a2 95 9d 97 9a 9e 9d 9e 9e 98 9e 98 a0 94 a6 a0 aa a9 b1 b5 be c8 c4 cb ca be bb ab ab a3 a8 9e 98 92 8e 90 92 92 94 9c 9e a2 a1 ab a4 a5 9e a1 9d a3 a7 a0 9c 96 98 9f 9f a6 ac b0 b1 a5 a3 a6 a7 a6 a1 aa 9f 9d 9a a6 a7 ab b2 b8 b3 b0 a7 a0 a7 a3 a8 a7 a3 a8 aa a5 a1 a9 a5 96 9e 9e ac b0 b9 bc c4 cb ea ff ff ff f9 fe ff ff ff ff ff ff ff ff fa ed e7 e0 db d0 c2 bb ae a9 99 98 9b 99 94 95 92 93 92 86 8a 7f 80 76 6b 5e 60 59 5e 52 56 49 59 4e 47 2d 1d 10 0d 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 10 21 20 28 2b 35 39 3a 36 36 3d 32 43 40 45 4e 50 46 50 52 58 53 60 5f 56 5a 5e 6c 6d 6d 70 76 7f 84 87 8e 91 a2 a5 9f ab a6 ac 9f 9a a3 a5 99 9f a3 a3 a3 a6 a5 a9 af aa a4 a9 a9 a5 a5 bb b5 be cf cb d6 d2 d0 cf be b5 ad aa a0 a3 9d 98 96 92 93 9e 9f a3 af b0 b6 b6 b6 af ae a9 ae b0 ad ad a2 a3 9d 9b a4 ae af a7 ab a5 a4 b0 a1 a8 a4 9f aa ac b9 bd b8 c3 ca c2 bd b5 b6 b8 b1 b6 b1 bb c0 be bf b6 b5 ab a4 a7 ae bc b6 bd c3 cf e2 ff ff ff ff fa f3 fa f3 ff fd ff f3 ff ee f1 e8 e5 ed df d1 c7 ba ae a4 ac 9a 9d 9c 99 a2 a3 9c 99 8f 8d 87 8a 7f 7b 6d 6b 6c 64 61 5b 63 65 63 61 4f 35 1b 16 0d 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0b 10 11 0f 14 2a 31 31 41 3f 44 45 3a 39 33 40 4a 51 50 5c 51 53 55 58 5a 5c 5d 5d 63 60 65 6d 7a 77 7c 7c 82 84 94 91 9b a5 b1 ac b2 ba b0 a2 a0 a7 a7 af ae ae ad aa ae b4 b2 b2 b0 ad b7 b8 b8 b7 be bc ce d3 dc e2 de d7 de c9 be b7 b2 a6 a7 a4 9d 9d 93 a0 a6 b7 b3 c0 c0 c3 bd c0 be bc bd b5 b3 b1 b3 a8 a7 a4 a7 b4 af b5 b1 a4 a3 a1 a0 a9 ac ae af c6 c3 c7 c6 d6 d4 d3 d0 cc b6 c5 c0 c8 d1 c8 d0 d5 cf d0 c3 b9 bd bb b6 b5 be bd c5 c8 e8 ff ff ff ff ff ff f6 f7 ef f8 f4 f3 ed ee e3 e3 e4 f6 ff f6 e1 cc c1 ac a6 a0 a2 9c a1 a2 9e a1 9b 94 a1 9a 9e 94 8e 87 7b 79 7c 6e 6e 6a 6b 79 86 76 75 58 3b 25 1b 12 02 0a 08 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 05 17 19 1e 24 25 35 3d 47 47 47
 46 42 40 4d 52 5b 60 5a 58 58 51 62 62 61 6b 5f 62 62 64 65 70 79 7a 82 85 85 88 8e 9b 96 a4 a9 a3 b0 b1 b9 ae a6 ab a7 b1 ae b1 b6 b4 b1 b9 b9 bc ba be c1 c8 c4 b6 bd c6 c4 c8 d2 dc e1 e4 e4 e4 d8 cc c5 b6 ad ae b0 a7 af ae b5 be c2 d3 cf cf df dd d8 d7 ce d4 c4 cc c9 c0 ba b7 ae b9 ae b0 b6 ba b1 a1 a4 a1 ab b7 b8 b7 c4 cc d7 e1 e2 de dd d7 d7 d8 d1 dc db dc de e6 dd e3 d2 cd d1 c3 c1 c1 c0 ca d0 d0 d4 f1 ff ff ff ff ff ff fe ff f9 ff ff f6 f3 ef e9 ec e1 fa ff f3 f1 e3 cd c6 b9 ac aa ac a7 a2 ab 9c a0 9d 9c a2 aa 9a 99 94 8f 8a 86 74 82 77 79 8c 9a 98 82 6e 52 3c 30 1e 13 0d 05 0f 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 28 27 2c 35 3b 45 4c 62 59 53 5d 61 62 6a 62 63 63 60 5e 62 62 67 68 69 68 6e 73 66 67 68 6f 7f 7e 85 90 94 97 97 95 9e a0 a9 a4 ab a8 a5 a7 a0 a2 ac ae a9 b9 b1 b8 c2 bf c4 c1 c4 c2 c9 c2 c7 cd ca cf d0 d6 e0 dd eb e7 ef ea d4 ce c3 c1 bd c7 c0 c1 c6 cb d4 da df ee f3 ff fe fc f9 f3 fa f4 e3 dc d1 cc c9 c1 c1 b4 bc b0 b6 c5 ba b0 ad ad b9 b8 bf ca d3 d5 df ea f0 f1 f0 ec ed ec e8 ed ed f1 e4 f1 eb e0 e0 d6 d2 c8 cb d0 cc d3 cf d5 e2 f3 ff ff ff ff ff ff fb ff ff ff ff f8 f2 ee e5 ed e6 ec de e0 ed ed ea e2 d0 c7 b5 ae b8 b0 b3 a8 ac b6 b8 aa a3 b0 ab 9d 9d 8e 8b 8d 81 7b 7c 89 9f b0 9f 87 70 56 39 25 16 07 06 06 07 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 09 07 1c 33 3d 43 34 4d 53 64 6e 74 78 75 77 73 74 75 71 63 6b 62 61 6a 6e 70 7b 7f 7f 7f 7e 76 78 73 79 83 8b 92 9f 9b a5 a3 a7 9e a5 a5 a1 a4 a4 aa a0 9f a7 ab b1 b1 b4 bc c1 c1 cd c6 cd cc d7 d1 d9 d7 dd d1 d7 db e3 ec e8 e6 f7 f7 e9 de e4 d7 d4 d9 d3 d6 dc e3 e9 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff fb dc d5 c3 c6 c7 b7 c1 b9 c4 c7 b5 b1 c5 bb cb d0 d5 dd e7 ed f6 ff ff fa ff ff fc fc fb fa f4 f1 f1 ec e9 e7 dc d3 cd c8 ca c5 cb ce d1 d5 e3 fd ff ff ff ff ff ff ff ff fc ff ea ef e9 e8 e8 e7 d5 d6 e0 ec f0 ff ff e9 dd d2 c5 c8 cb c8 c4 c5 c9 c6 b8 b6 b4 b0 b5 a7 a4 96 97 8e 81 85 86 9a b6 bd a7 90 66 51 3c 2a 18 14 0a 10 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0b 05 0d 17 1e 34 4c 4d 57 57 69 65 83 87 7f 83 7d
 6c 72 78 70 6c 64 65 57 64 7a 7a 7f 8d 8a 8e 8e 91 91 86 8b 83 8b a0 a3 9e a0 a6 aa ab a4 aa a1 ad a2 9e a1 a4 a7 ab a1 b4 b1 ac be bb cd ca cf ce d7 d9 db e2 e1 e5 e3 e6 e7 e8 ea ef f8 ef f4 f3 f4 f0 f1 f1 f0 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb d6 ce c6 c9 c1 c2 cd cc be c1 cc cd d0 de e1 ea eb f3 fb ff ff ff ff ff ff ff ff f9 fd f1 f0 e8 db df d8 de cd d3 d4 ca d2 d0 d1 d4 df ed ff ff ff ff fc f9 ff fe f5 f9 f8 f0 ec ea e5 e1 df df e6 ef ff ff f8 ed ef e3 d7 d9 d9 cf dc d3 d6 cd cc cb c7 c0 c0 b8 a8 a2 98 8e 8d 8d 86 8f a4 ca c7 ac 85 64 49 37 20 17 1c 14 12 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 08 1d 21 2e 48 4b 5f 61 6e 6d 75 73 70 68 6f 70 66 6c 68 63 63 61 60 60 65 70 70 78 8b 93 99 9e 99 99 95 9d 97 98 a5 9a a4 ae a5 a9 aa a7 a0 a2 a0 9c a0 9d 9e a1 ac a7 b1 ac a5 b3 b7 bd c6 bf d0 d0 d7 d6 e0 e0 e4 e6 e3 e9 ed e4 ee f2 f2 ff f9 f7 ff f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e3 d4 c9 cf d1 d6 cc cd d3 d3 d9 e3 e3 ea e9 f6 ff ff ff ff ff ff ff ff ff ff ff f6 ee ec e8 da df d5 d8 d2 d7 cf cc d2 cd cc ce d8 e0 f6 ff ff ff ff f8 ff ff fd f6 f1 f0 f3 eb f0 eb ec df d4 e6 fc f3 ed eb f2 ee de d8 d7 db d9 d8 e4 db d6 ce ce ce c8 b8 af 9f a3 99 9b 93 92 8b 94 b4 da cb a2 7f 60 48 38 2a 21 11 0d 10 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0b 1b 27 36 45 50 67 6f 85 8c 8d 88 75 6b 5f 61 6c 66 6b 64 6a 5d 60 6b 6a 6c 6f 8d 85 91 9a 96 96 a4 a4 a0 a8 a4 a6 a8 ab a5 a9 a3 9c a2 a6 a0 9e a5 9a 9d a7 9e a7 9f a1 a5 a9 af b6 bd bc c1 c6 c7 ce db d4 e4 de e6 e9 e2 dd ec ea f5 f4 f1 f9 f4 fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee e2 e5 d8 db d1 e0 db de e0 e4 ed eb ee fb fb ff ff ff ff ff ff ff ff ff fd ff f5 ee e7 e1 db de d4 d3 cf cc cf c2 c8 d2 cb ca c9 d2 e4 ea f7 ff ff ff ff ff ff fb f3 f6 fc f6 f6 ef df dc cd d9 e7 e7 f0 ed f9 f5 dc df d1 dc dd d6 dd de d1 cb d0 c9 c6 be b2 a7 a3 96 8b 95 91 98 9e ac d6 e5 c9 9a 85 5e 4b 3e 2a 24 1a 16 0c 01 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 22 30 32 4c 5a 6a 7e 8c 9d a1 98 92 7d 68 65 69 61 67
 73 6a 6e 73 6c 74 77 76 88 87 8f 96 97 a5 a5 a2 ad a0 a3 b1 af ab ad b1 a6 aa a5 ad a7 9e a1 a0 9e a2 a7 a2 8a 9b a4 a3 b3 b1 b0 be c6 bf cd d2 d7 d7 db dd de e3 ed e9 e8 ea f6 f2 f2 fa f9 fc f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 ef e7 eb ea e3 e2 ef ea f3 ea f3 f6 fe ff ff ff ff ff ff ff ff ff ff ff f1 ea eb f1 e8 db df c9 cd d7 d2 cb c9 d2 ca c3 c6 c1 ca cf e0 ea ef ff ff ff ff ff ff ff fd ff ff fb ea d4 da d3 df e7 fa ff f6 e9 e6 dd d8 d8 d4 dc df e5 db d2 db c7 cb c9 c6 b9 b5 a9 9d 9f 9f a3 9f a4 9e c2 f2 e5 c4 a4 89 67 55 48 31 22 20 1b 0c 08 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 19 27 33 43 53 6a 7d 91 9d 9f a2 95 80 6e 6f 72 75 72 77 78 75 72 79 81 78 7e 88 93 99 97 98 97 9c 99 a2 a7 a3 a6 b3 ad b3 a5 a4 a5 a5 a7 9d 98 a2 9b 93 99 94 94 98 9b a2 a0 9d a8 a9 b3 b7 c2 c7 c6 d1 cd d1 e0 db e5 de df ed ed ec f6 f2 ee f6 f9 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f3 f1 f2 ec ed f2 f0 f3 fc fb f6 ff ff ff ff ff ff ff ff ff ff fd ff f2 fb e6 e7 e4 db d7 d0 d6 d4 d6 d2 c8 c9 c7 c5 c7 c4 c4 c8 d4 d8 e4 ee fc ff ff ff ff ff fd ff fa ec e0 db cd d4 dc e6 fb fd ee e5 d8 d2 ce d0 ce dc e5 de d2 cd d0 c6 da cf ce c1 c3 b7 ab a3 ab a5 a3 aa a3 ab d0 f7 e9 cc af 88 77 59 4b 34 2e 24 12 0c 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 20 28 34 47 5e 79 86 91 96 94 88 82 78 75 75 72 7c 7e 7c 81 7a 76 7c 7f 80 86 8b 8e 90 8f 9b 99 9e 9f a3 a2 a7 aa a6 a5 ac a9 a6 a7 a3 a2 96 98 9b 9a 93 98 95 8d 9d 94 93 a0 a2 ac a3 b6 b5 c1 bf c4 ca d4 d0 df db dc e0 e9 e8 ea eb e5 f2 f2 f4 f6 fb fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f7 f9 f8 fa f2 fb f5 f7 fb ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ef f1 e5 e6 e0 da db d4 d3 cf cd c3 c6 c6 cf c6 c5 bf c3 c0 ca d7 cb d9 e7 f7 ff ff ff ff ff ff f9 e2 e0 df d8 dc ea f7 ff ff ec e2 d8 dd db d9 dd e1 ed dd d1 d2 d1 da e8 e4 e4 d1 c1 c6 b4 bb b8 be ae a6 a1 a3 b2 dc eb ea cb a9 93 6c 59 4d 35 28 1a 18 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 04 07 08 1d 27 32 35 4d 5f 6e 72 7f 7c 7d 75 71 7a 7e 7a 7f 83 89 7e
 81 88 85 84 89 8f 89 90 95 9a 9a a0 a2 a3 a3 9f a2 99 a2 a4 9d a0 9c a1 9e 9d 9d a3 9c 9a 97 93 96 95 8e 91 8b 90 a2 a5 a5 aa ac b8 be c3 cb d2 d7 d1 df d9 da e0 ea e3 e5 ea e6 f0 f0 ec f1 ec f5 f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f0 f0 ea e6 e9 e3 e3 dc d8 d1 d5 cd c9 cc cb c9 c4 c5 c8 c8 c4 d1 cd d0 d3 dd e6 f5 fe ff ff ff ff ff fd fb fc f9 fe ff ff ff f8 f0 ea e0 ec ed f6 eb e7 e3 d8 de e2 f0 f5 f1 f0 d5 d3 cd cd c8 cb c0 b3 b4 a8 ab aa b5 c8 ec eb dd c1 a2 82 60 49 31 1c 0c 08 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 09 0c 0d 14 22 2b 31 41 4c 5d 61 70 6a 6f 72 79 7d 7e 83 85 8c 8d 8f 8d 8e 93 8c 8f 92 91 93 91 93 9c 97 94 9e a0 a2 9a 94 9a 9d 9f a1 9d 9d 9d a8 9c a2 a1 98 96 8f 95 9c 92 93 91 96 9b 9d 9a a4 a1 ab bd bc c8 c1 d1 cf d6 d8 df e6 de e7 e4 e4 e4 e9 e9 e8 ea ee f2 f3 ef f6 f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f6 f5 f5 ee e8 e4 e4 db dc df d1 d5 d3 c7 cc cc bf bd c2 c9 c9 d4 cb cb c4 cc d4 d3 d5 d4 e3 f2 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff fa ee f6 f8 fe f9 ec eb e1 eb f9 ff ff ff f9 eb f2 e7 dc dc d3 cc c2 bf b1 b4 af af b4 cb e6 e8 d7 be 9e 77 60 45 2c 1e 0f 04 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 09 15 23 22 28 36 46 5c 67 61 5a 70 70 72 79 76 85 83 8c 91 89 91 91 9b 90 9a 94 99 91 90 8c 98 96 95 9c 99 9d 9f a1 9d 98 9e 91 97 9c 99 96 96 97 9b 9a 95 9c 91 92 8d 89 8f 94 9d 9b 9d 9d a4 a6 b6 b9 c1 c1 cd c9 cd ce d7 d3 e3 e1 e1 ea ea e9 e3 e1 e0 e0 ec e7 eb f0 f2 f5 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 f2 f1 f0 ed e4 e5 e2 de d4 d1 d4 cf c9 c9 c7 c9 c3 c5 c8 d2 d2 d2 cc cd ce d0 d2 d1 d1 d4 cf e0 e4 e9 f1 f5 f9 f3 e7 ec ec fc ff ff ff ff ff ff ff ff fb fc fb f2 f4 fb ff ff ff ff ff f9 eb e8 dd d9 d3 ce c3 bb af ac b0 ab b2 c2 cc e1 cc c1 99 73 51 34 27 19 13 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 19 20 27 33 31 3e 4c 5d 58 5f 58 5d 68 76 7c 7b 82 80 86 85 8f 91 92
 9c 9f 93 98 9b 9a 90 94 94 9c 99 97 a1 9a a2 99 9d 8f 98 9c 97 95 9a 98 94 94 95 9c 88 8c 8b 8d 8f 93 97 9b 96 93 9b 9d a5 a4 a1 b6 ba bd c9 c5 d3 d6 e0 da d7 e0 e6 e6 e1 e4 e4 dd e4 e2 e8 e2 ed ed ee ef f8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f8 f7 f5 ef e7 e1 e5 e1 df d4 db d8 d1 d1 c8 ce cc c2 c7 c6 d3 d4 d6 d6 d0 d1 d6 dc d1 d5 d3 cf d9 e2 dd e1 d9 e1 db e0 de e5 ef f5 f7 f9 ff f9 f8 ff ff ff ff ff f1 f5 ff ff ff ff ff ff fe f2 ee e8 db df dc c8 be ba a5 a5 a6 a6 a7 b3 bd d1 cb b0 84 61 47 3a 34 16 10 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 21 25 34 39 45 4d 53 56 5a 57 5e 62 67 76 76 7e 81 84 86 8d 93 93 96 97 9f 91 94 96 9b 98 96 93 97 9d 99 9a a1 93 a2 99 8f 96 99 93 a1 9d 9c 90 90 96 93 94 8c 92 90 89 8b 90 95 97 98 a2 a0 a4 a2 ae ba bf bf c3 cc d4 d5 de de e3 e4 e4 de e4 e0 e8 ea e0 de e7 e0 e7 e5 ea f1 ec f5 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fb f3 f5 f1 e8 e9 e7 e0 d7 da d3 d5 cf d2 cb d2 d3 cc cb d2 d7 e0 d4 d8 d5 df d5 d9 cb d1 d7 d7 d7 d7 d8 dc db d5 df e6 df e8 eb e9 ee e7 ee e9 f3 f2 f1 f4 f7 f9 f8 f1 f6 ff f8 fb ff f6 f9 e9 ed f2 e6 e5 d5 ce c6 b2 ad a3 9f a0 9e 9b a6 ae be ae 95 75 58 45 35 2c 1d 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 14 1e 27 3a 4d 5b 5d 57 59 5e 5b 65 6b 72 74 7a 7e 81 84 8f 94 8d 88 96 98 99 95 91 95 9e 91 9b 99 8e 9b 95 94 98 93 92 97 8b 94 8c 92 a0 b2 a2 93 92 8e 91 8c 8c 90 8c 90 92 95 93 96 a3 9c a5 ac a6 ab b4 bd c2 c9 cf d5 da e3 e4 e7 ea e6 e4 e8 df e4 e4 df e3 e4 dc e7 df e2 e5 eb ed f3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f5 ee e9 f2 eb e5 e3 e0 df dc d0 d1 ce cf ca d4 d5 d4 d0 d2 d5 d8 df d7 d9 d5 d8 e1 d4 db d5 da da da e2 db de de e4 e1 e6 de ec e3 ec e5 e2 e7 e6 ea e7 ea ef eb eb ec eb ea eb ed f3 eb eb e1 e1 d7 df d7 d5 c4 c3 b3 a7 9c 9a 9d 98 93 98 90 92 98 8c 7b 6f 52 39 2b 23 17 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 07 06 11 27 26 38 42 49 64 5b 5d 64 5c 70 6b 62 71 7a 82 85 87 8d 8c 8e 92 93 96
 98 96 91 8e a1 94 96 99 92 99 96 98 a9 a2 95 9c 93 91 8e 87 8f 95 9d 9a 9a 8c 86 8d 89 8b 92 94 93 98 96 97 9a 9a 9d 9f a8 ac b4 b9 c0 c0 cb ce c7 d4 de e5 e8 e3 e6 ea e3 e2 e9 de df db d9 e1 e7 db e6 e9 eb ea ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ef ef f0 f0 eb ed ea dc dd e1 dc da df d8 d3 d8 d3 d8 d5 df d6 e1 dc e1 e1 e0 e5 e8 d5 e2 de d9 dc ea e8 e2 e6 eb eb e6 e5 f0 f5 e5 ed eb e9 e7 eb ed e0 e6 e6 e9 e5 e7 ef e5 eb e3 e3 db db d6 d0 cc c7 c5 c1 bd b9 a9 a0 a6 99 9e 9b 99 92 87 8f 89 83 8a 75 58 39 2c 24 18 08 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 0e 16 25 31 35 46 4d 64 5e 66 5e 69 73 6c 73 79 81 82 85 8c 8e 92 8e 95 87 9b 99 94 8e 8d 95 92 97 8d 97 94 96 8e a3 9f 98 99 95 90 91 89 8d 8f 8f 90 99 91 87 92 8d 8a 87 93 94 94 94 9f 9d a3 a0 ab ae ac b2 b5 b9 cb c6 cb d8 d7 e6 e5 e4 ef f1 ec eb e5 e5 e0 dc e1 e1 df dc dc de e5 e7 e7 f0 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f4 f9 f7 f4 ed f2 ee f3 e7 dc e2 e0 df e0 e1 db d8 d8 dd dc d7 e0 e3 e4 e9 ea e1 e0 ec df e2 e7 df e0 e6 e7 ec f0 e2 e8 ed e8 ee e9 f3 ea e8 eb ec e4 e6 ee e7 dc e6 e4 e2 e4 de d6 db df de d6 cc ce c2 be bc b7 ad b0 a6 a0 99 9c 9a a4 94 90 89 79 7e 88 8a 79 60 42 35 25 1c 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 06 0f 12 18 33 4a 4b 56 53 5c 57 56 63 5d 6b 6c 75 84 7d 89 89 8a 90 8d 99 91 90 94 90 8b 91 93 90 8d 96 97 93 8b 95 95 93 95 90 9c 94 8c 85 85 8c 8c 88 8c 91 93 90 81 88 88 87 8f 95 94 98 9a 9b 9a 9b a2 a8 ad b2 be c1 c3 c9 cb d8 e0 ea e5 ea ee f1 ec ec e8 e7 e3 df e7 d3 da d8 e0 da e4 e2 e0 ee f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe ff fa fe f3 f0 f2 f4 f3 ed ec e0 e0 e5 e4 e1 e0 db e4 e1 e4 e0 e3 e5 e6 ed e9 e2 ec ea e2 e2 e4 eb db ea e8 e4 e6 e9 ed ed ec f2 ef f0 f0 eb f5 ea e6 e4 e6 e5 f1 e2 e1 e1 d9 de da d8 d4 d2 cd c3 c4 c2 bd b8 ba a9 a6 a7 a1 9f 97 a0 9d 9c 92 8f 81 7e 7c 7f 92 80 61 4d 39 2f 14 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 03 06 05 03 10 19 2a 55 56 67 61 54 5c 5f 57 5a 62 71 75 74 7a 76 86 87 88 85 7f 92 8e 92 95
 97 90 88 86 8e 8e 92 8e 94 92 8e a1 96 8d 96 98 92 90 8f 8b 8f 8c 85 90 9d 91 92 88 86 89 8d 93 95 98 8f 99 9f a6 aa af b4 b2 bb be cb ca cb cb dd dc e3 eb ee f0 f6 e8 eb e8 e9 e4 e2 dd df dc d9 e6 da e0 de e6 e9 e7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fe f3 fc ff fb f7 f8 fb f1 ee eb e4 eb e6 e4 e4 ea eb e8 f0 e6 ed eb eb e7 f3 e4 f2 e6 eb e3 e8 e9 e2 e8 ea e5 e1 e9 e4 f3 ec ee ee f3 f7 f3 f1 f4 eb eb e4 e4 e8 dc e5 d4 d1 db d6 d7 c8 cf c5 c7 bd b9 b1 b5 ac a3 a6 9d 91 94 9b 92 9b 8f 95 85 88 83 7f 97 9f 83 68 52 3d 2c 18 13 04 00 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 09 1c 25 3a 62 66 66 69 5c 5f 61 61 5f 68 6e 74 7d 7e 7c 84 87 82 8c 8e 8e 8a 8f 7e 85 8a 7e 79 89 81 86 93 95 84 96 96 97 90 94 8e 8f 93 8b 9b 94 90 90 95 90 9a 92 87 8f 8d 90 8d 91 95 9e a1 a5 aa a9 ab bd b7 c2 c3 cc d0 c8 d5 df dd ea ef ed f1 f4 ed f0 e9 e6 e7 e0 df de d9 e2 da e1 db de e2 e7 ea ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff f8 f8 f7 f5 f9 fa f4 f4 f8 eb e7 f0 f3 f6 ee f1 ef f1 f2 ed f1 f1 f2 ed ea ed ed e6 e8 df ea e4 e0 ec e5 eb ed e1 ed e5 eb e9 f4 f5 e9 f0 eb eb e9 e4 ea ed e8 e3 de de d0 d4 d1 d4 d5 c0 c2 bd b3 af a8 a8 a3 a3 a0 a5 90 93 95 8f 8e 9d 8d 8e 78 76 85 94 a5 96 70 58 46 38 2b 1a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 0e 19 31 49 71 76 6d 68 6a 5b 62 60 6c 72 6f 6b 76 80 7d 7f 7e 7f 81 87 82 8d 89 81 82 7c 7d 79 84 82 84 8b 8b 84 86 8e 92 97 95 95 90 9c 94 95 97 94 8d 90 8f 8c 90 94 95 8f 88 93 93 96 9c a0 a1 ab a7 ad b7 bf ce cb d2 d5 d4 da e3 e8 ef eb f0 fa f2 f4 e9 e5 e8 e4 e2 df d6 d9 d3 d4 da dc e1 d5 e8 e8 ec fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 fe f5 ff fe f8 ff f7 f6 fd f6 f4 fb f3 ef f2 f9 f0 f2 fb f3 f6 f3 f7 ec f0 f1 eb e9 e7 ee e2 ef ee e4 ee e6 e1 e6 e6 ea e6 e4 e6 e5 eb ed f0 e7 eb f0 eb e5 e4 e0 e2 de e0 e0 d9 df d6 d3 c9 c9 c2 c4 bb b1 a8 a1 9d a0 99 a0 95 93 8e 90 93 95 8e 8e 8b 86 74 75 89 95 b0 93 7a 55 39 35 25 19 0b 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 10 09 16 2d 42 5e 71 80 73 6b 69 6f 65 67 70 71 76 72 6d 79 78 82 7f 82 80 83 83 81 87 7d
 80 77 7b 80 79 7b 79 81 79 84 87 8d 95 96 9e 96 a4 a0 97 a6 9f 9b a2 96 9a 98 95 8f 95 91 96 9f 98 9b a1 a5 af af b2 ba bf c0 cc cc d1 d2 d8 d8 e7 eb eb f5 ef f2 f7 ee ed f3 ee dd e4 e0 da dd dc de da d9 e0 d5 e7 e9 ed f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f9 fa ff fc fe fc fe fe ff f6 ff fc f4 f6 f4 f9 f8 f0 f2 f3 f0 fe ed e8 eb eb ec ed f2 e8 f0 e4 e6 ea e6 e2 e3 e7 e7 e2 e0 eb e6 e9 ea e6 e4 e6 ee e3 e6 e3 e1 de e1 e0 da d8 d5 c9 cd c8 c4 c2 b6 ad b2 ab a1 9c 9d 94 9a 96 96 94 92 8e 8d 8c 80 7f 7f 7c 7b 81 aa b0 a4 7e 62 4d 39 2e 26 12 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0a 14 1f 2f 44 69 8b 8b 75 73 6b 70 6f 71 6e 7b 77 6f 6f 7d 7c 7d 7a 7a 77 75 76 7e 83 81 79 79 78 82 83 78 7a 83 83 80 7d 85 8d 94 a2 9a a6 a7 ab a9 a7 a3 a6 9f 9e a2 95 97 95 98 9e 9a 9c a0 a4 a9 ac b2 bd c7 ce ca c6 d2 db d8 e7 e0 e2 e9 ee ef f5 f4 f5 f2 f2 eb eb e7 db dc d5 dd e1 e2 df db d9 df e3 e5 ea ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fe ff f6 fc ff fb ff fb fd ff f4 fe fb f6 f6 f5 f6 fa fe f0 f8 ee f2 eb ec eb e9 f0 e9 e0 ee e9 eb e6 df e4 df e1 e4 ea db e4 e7 e0 de e3 e0 e4 dd da d9 db e2 d8 dd d5 d4 d1 cd c7 cb c5 be be bc bb ab af a5 a3 9c 9c 94 94 96 90 8b 93 92 8c 83 84 78 84 7a 84 84 ad c3 9f 88 62 52 4e 39 32 20 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0c 0b 0e 1c 25 39 4d 6f 8d 99 7d 6e 6d 6f 76 71 73 7e 77 7d 7b 73 73 7c 72 79 81 7c 79 75 74 73 84 76 7c 78 82 74 7f 7c 7f 8a 89 8c 90 90 97 a7 a8 ad b0 ad b2 af b1 af b5 ad a0 a5 9d 9b 9f a4 a3 a7 a9 b3 b5 ba c1 be c9 ce db d4 d4 df e0 e1 ed e7 f2 ea f0 f1 f1 ea ef eb ec e4 e5 e3 e2 df df d7 d7 d8 dd dc de e4 e3 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff ff f6 fb ff fb f5 f9 f8 fe fc fc f9 f8 f1 f8 f1 f8 f1 f4 f2 f0 ed ea e6 e0 e1 e1 e2 e5 e4 e3 e7 e1 df e1 d8 df dc dc da db de e2 dd e1 d6 e3 da d8 de dc d4 d3 d2 cf c9 ca ca c9 c6 c1 ba b5 b1 b0 ae a8 a0 a0 96 95 96 8f 92 94 8d 8c 7d 81 83 81 7e 80 74 7d 81 b3 b8 aa 8e 72 64 55 3c 32 20 10 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0f 1a 28 3b 4f 65 7f 95 9f 88 79 76 6f 75 77 73 76 76 76 80 7c 82 81 84 7f 87 7b 72 7d 7b 75
 76 77 79 7a 73 86 77 80 83 87 84 8e 8c 95 9d a3 a6 ab b5 ba c0 c0 b9 b8 b9 b6 ac ae aa 9f 9f aa ab a9 a8 b0 b8 be c2 c7 cd d2 d3 de db e5 e7 de eb e9 f1 ec e9 eb e2 e9 f2 e4 e9 e0 e0 de e4 d7 d7 d5 da de d8 db e3 e2 e3 ea ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe ff fe f9 f7 fe f7 f7 f9 fd f7 fd fc ed f6 f9 f2 f2 f5 f0 f6 ee ee e8 e8 e7 ec e4 e4 dc dd e2 de dc d8 e1 df db df db d5 d6 d5 d8 d9 da d7 d7 d4 d8 d5 d5 d6 db d5 cf ca d2 c3 c7 bb b5 b7 b2 b8 ad ad a7 aa a6 a2 93 94 92 95 98 92 92 8d 8b 8b 86 7f 83 80 80 78 7e 7c 8a ad bc a5 97 77 65 57 45 36 20 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 10 1a 25 2d 42 59 73 8c a7 a5 86 77 7c 75 73 75 77 7e 7d 7e 76 7a 7b 86 86 82 81 7d 7b 7c 80 78 77 74 7f 73 82 7b 80 85 8c 88 8c 8e 97 94 97 aa b0 ba bb c2 c0 c6 c7 ce c0 c0 bd c0 bb ba b1 b7 b5 af bc c3 c7 cd be d3 d8 dc dc e3 e1 e2 da e4 e6 ec ea ee ec e8 ee ee e7 eb eb eb e2 df e7 dc de dd db df dc da e1 e3 e5 e6 ed f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fb ff fb ff fb ff fa fe f9 f7 f9 f5 fa f9 f6 f9 f3 f0 f3 f1 ed f5 e8 ed ea ee e7 e6 e6 e0 d6 df d4 db dd d0 e0 d6 d1 db d7 d4 d3 d8 d3 d8 d9 ce d9 cf cc d2 d2 cf d4 c5 ca c6 cb bc c1 bb be b7 b4 b0 ae a2 9e a2 95 9b 97 99 8e 84 93 8f 91 8a 86 82 7b 78 7e 71 71 80 7f 7b 8d aa bd b0 9a 84 6a 63 4a 35 20 0c 07 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 11 2b 36 42 56 61 7d 95 b3 b4 85 77 77 7b 78 75 75 73 74 7c 77 78 85 80 7f 77 7b 7f 75 76 7f 80 7d 77 7e 84 88 82 8c 88 8d 98 8d 92 9e a3 a9 b2 bc c9 c8 cd c7 ce cd d2 d3 ce cb cd ce c8 c7 c8 cb c3 c1 c9 cd d2 cb ce d2 d8 dd e4 d8 dc e1 e1 e9 e3 e5 ec e7 ee ee ec e5 e5 e9 df e3 e1 dd d6 de da dc d4 de df e5 e3 e3 ec f7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff fa ff fd f5 f8 f5 f6 fa f3 f6 f3 f1 f8 f3 f5 ef ef f8 ef ed ec f0 e5 e4 e3 e4 de df db de df db d8 d0 ce d3 da ca d2 d2 cc cd d2 cf ce d3 cb d1 d0 cd cb ca d2 c9 d0 c5 be bc b5 b4 b7 af b0 ae a3 ab 9e 99 9e 99 97 99 8a 96 95 8c 8d 84 85 81 7d 7d 76 76 64 77 70 72 7b 81 82 94 b6 b3 a5 89 7a 69 55 43 1a 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 20 26 3c 46 5b 76 8f aa bd a7 87 80 76 6f 7b 7d 72 7a 7b 6e 7a 70 7f 7a 76 7c 75 7f 7e 7b 78 80
 7c 7c 81 82 87 8e 8a 91 94 90 9a a0 a3 ad b2 b8 c0 c1 d4 d0 d3 d9 da d7 da df d3 cd d2 d2 c6 c9 cc c5 d0 c9 cc d0 d2 cd d5 d5 da de da d8 db e3 da df e0 e0 ea e7 e4 d8 e4 de e6 de e5 e0 de dd db da d7 d8 cf db e4 e6 e5 ed f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fd fc f9 f6 f2 f7 f4 f9 f2 f5 ef f2 f6 ed ef e6 e9 e9 e9 ef e8 e7 ea e3 dd da e0 d5 dc d4 d7 d4 d3 d6 d5 d4 c7 d4 c7 cd cf c3 cf cb c7 cb c9 c5 cb c8 cb c6 c4 c9 bb bd be bc b4 b5 b5 b1 a9 a5 a3 a0 a0 a2 95 9b 97 90 8c 92 8c 87 81 85 7b 78 79 75 6b 6d 6f 69 67 6b 6d 75 76 76 81 9e b1 a3 8e 78 6f 4b 39 23 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 17 26 33 46 59 65 7f 9e ba b7 9e 80 75 7a 79 76 79 7b 7b 79 7c 7a 7a 7e 73 77 79 7f 7b 7c 78 7f 7c 83 86 82 89 91 8c 92 98 99 9e a5 a5 ae b0 b6 c6 c9 cb da db d9 e1 e4 dc e3 d6 de d2 d9 d6 d1 d4 d9 d0 d3 d5 cb d5 d5 d5 e0 d5 d8 d9 d7 da d1 da de d5 d5 d9 da e5 dd df e3 d8 de e1 de db de d9 dc d1 d9 dc db dc e4 e4 ea f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff f8 f5 fe f5 f3 f9 f7 f5 f2 f5 f0 ea e8 f1 eb e7 e8 eb f0 e4 e1 ed e3 e4 df e0 e4 dd d3 d4 d5 d3 cb ce ce c9 c9 cf ce cc c7 ca c0 c4 cc cc c3 cd c6 c5 c0 c0 c4 bb be bc b7 b0 b4 a6 ad a4 a6 a5 9e a1 94 93 8d 93 90 8f 90 8b 86 83 7e 7e 75 75 70 67 67 6d 6c 6c 67 6c 6f 70 75 7f 8a aa ab 98 80 71 55 37 1a 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 09 28 29 36 57 63 74 90 ab b2 ab 85 71 71 6f 74 72 72 76 74 7c 74 77 7a 72 75 7b 7c 7b 82 78 79 79 7c 87 86 86 89 8d 94 95 92 9a a3 a2 ac b2 bd bc c9 c9 c6 d6 db d6 da de dc e5 e1 d9 db db d7 d9 d5 d3 d9 d2 d5 c7 d1 d7 cc d5 d9 dd db dd dd e4 e1 dc dc de dc db d9 e1 dd dc e3 de df df e0 db df dc e5 e1 d9 e0 e0 ea ea f1 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f7 fa f9 f3 fe f0 f4 f7 f1 f8 f4 fa fb f6 f1 eb ef ef e6 e7 e4 eb e4 e7 e5 dd df db de dc d7 d5 d4 d0 cf cb c9 cd d1 cc c9 cb c9 c9 cd c4 ca c2 c1 c5 c0 be c1 c1 c1 b8 bc c0 ae ac ab ab aa 9f 9d a0 9a 9a 99 93 90 8f 8b 8a 89 85 89 88 77 7c 7b 75 75 74 64 69 70 6f 68 71 6f 6f 6a 69 7d 95 a4 92 89 6b 4c 38 16 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 13 1e 36 43 50 66 83 9f a7 a7 8a 70 6b 65 71 70 78 72 6f 76 79 74 7e 74 73 7b 7b 72 77 79 7b 7c 7b 7d
 8a 81 89 84 84 90 8e 99 a1 a3 ab ae ba b6 bf c7 c5 cc d4 d2 d2 dc dc dd d7 dc df d7 d1 d8 d6 d0 ce d0 d0 cd cd cd d2 cf d7 cc cf d9 d8 df db e1 d9 e0 e0 df e0 dc e0 cc dd df d2 de d6 de e3 de da d5 d9 dc d9 de ea ed f8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb f8 f7 f7 f8 ff ff fc fb ff f8 fd fa f7 fb fc f4 f2 f6 f2 ed ec ec ed e7 e9 e1 df df da cf d1 ca cc cc ca c6 d1 ce ca c6 c8 c5 bf c3 c4 be cc c4 bc c2 bf c1 b9 bd c0 b5 b6 b4 ab ad a4 a5 ab a6 9f 9a 8b 8f 95 8b 93 8c 8b 8d 82 8b 7d 7f 7e 7b 74 64 71 6f 6b 64 70 6d 69 66 67 6b 6e 73 7b 88 a1 9b 7c 64 4e 30 19 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 18 25 3e 4f 5f 7b 94 a6 a6 94 78 6b 6d 65 6e 70 6b 72 6f 70 76 6e 75 73 71 73 7b 73 78 82 76 80 85 81 83 7f 86 88 87 8c 96 9a 9e 9e a9 af af b7 b7 c2 d0 c7 cf cd cf d6 db d5 d7 d4 d3 d7 da d4 ce cb cf d2 c7 cd c7 c6 ca c5 d1 d1 cd de db e2 e4 dc e0 e6 e4 e4 da dd da da d6 d9 db d9 e0 df d1 d6 dc dc d6 dc e3 e4 e9 e9 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 f4 fc f0 f0 eb e7 df e7 e8 dd d5 d1 c6 c6 cb c5 cd c2 bb cd cd c3 d0 c4 c4 be c5 c9 bf c4 bf b9 bd be bb bb bb ab b0 b5 a8 ab ac a0 a5 9b 9d 98 93 95 90 8e 8f 8d 86 8d 87 81 85 77 7b 71 68 76 6b 6c 6c 72 74 69 6e 6b 6a 6f 72 6d 79 7c 94 94 80 68 4d 2d 18 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0a 16 31 40 56 70 81 9e aa a0 7f 73 6d 69 62 6b 6f 6c 6c 70 73 76 7b 79 7a 6d 6f 6c 6f 75 7b 7d 7c 7e 80 89 7e 84 84 88 87 8e 94 9b a0 a3 ad b0 ba bb bb c0 bc c7 c8 c8 ca d0 d0 c8 ce d4 c0 c9 cd be d2 ce c6 c4 cc ca ce d0 cd d7 d5 dd dd db e0 de e6 dc d5 e0 db e2 e4 e1 d8 e1 dc df d9 de dd d9 d8 df df db d7 d5 e1 e7 ed f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fd ff fd fe fe fe e9 f1 de d2 d5 d4 cd d0 c7 ca c7 c5 c4 c6 c6 c4 ce c3 c4 c5 c4 c4 c6 c0 c0 c4 be c1 bc b8 bf b6 bc bc b6 be ad a4 a6 ac 9f a6 9c 9a 94 99 93 97 8d 90 8b 91 84 83 80 6f 72 74 6a 71 77 6f 6e 70 6f 69 6a 6c 6b 71 6d 6c 6a 78 91 93 80 6b 4a 27 14 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 06 0f 16 30 47 59 7b 8b a5 a7 8d 79 72 6c 67 68 64 67 6e 6c 70 76 6f 73 75 78 77 71 6d 73 77 75 73 71 7b 71
 84 80 7a 80 86 86 8f 8e 91 9b 9c 9d a6 ae b2 b5 c1 be bb bd c7 c2 cb c8 d1 ce c1 c5 c1 be be bd b9 b7 bd ce cb cd d2 d0 cf d4 d5 e5 e0 dc e3 df dc df e3 df dc e1 e2 e1 e2 e3 e0 e4 da e1 e0 dd db d8 ea dd e5 df e4 e8 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fc ff fc f8 fa fa f6 f4 ef e8 dd d0 ce d1 c8 c7 c4 c3 bc c0 bf c0 ce c2 c8 be bf c4 c1 c0 c7 be bf bf be c2 bf b9 ba ba b3 b6 ac ab a9 a6 ab 95 9d 99 9e 9a 92 96 90 8a 8e 91 91 89 85 79 7a 73 74 76 77 73 6b 6d 71 6a 71 6c 6a 67 65 64 6d 62 6c 71 87 93 7d 66 40 2c 10 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 05 13 24 41 4e 5f 7d a0 ac a8 88 70 6e 6f 6d 6a 65 6e 6b 6b 65 70 6a 6e 67 6f 70 72 72 70 72 74 72 79 86 81 7f 79 7a 79 83 82 82 86 8e 8f 92 a5 a2 a6 af b5 bd c1 b3 bf b5 bf c7 be c8 c3 b9 bd c1 be bd b9 c1 b9 bf be c9 c6 cf cf d0 d2 db d8 e2 e5 dc de d5 d0 dd da dc e1 ea e4 e4 e4 e3 e2 df e5 e8 e2 d9 e6 e5 db ea e0 ee f3 f1 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc f8 f6 fa ff fb ff ff ff ff ff ff ff ff ff fc fc f7 fc fc f9 fa f1 f0 f1 ea e4 dc e6 d7 d1 c5 c2 be bb c3 c2 be c6 c0 bd bb ba c6 bd ba bb bf bd bb ba c4 bd bd c5 c0 c9 b9 c1 b9 b2 b2 ac ab aa a8 a5 a8 95 9a 97 93 96 91 95 97 92 89 87 88 7e 71 78 72 73 76 76 6a 75 71 78 6d 6e 65 6d 63 6c 6a 68 6f 7b 82 8d 7f 5e 45 2a 10 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 16 2c 40 4e 6d 8a 9f ad 9f 79 75 6f 70 6e 63 63 66 63 6c 71 6d 71 70 6d 6e 78 73 70 71 78 74 6c 7b 7a 75 74 78 7e 7d 7f 7f 85 8b 8a 8c 97 99 9d a2 ab ae b2 ba bc be bd bf c5 bb bf b7 bd be c0 b9 b8 bd b4 be b9 ba c4 bb c2 ca da d5 db e2 e0 de d9 d4 db d2 d0 d8 df e0 e1 e0 e8 e1 e1 e1 e0 e7 e8 e7 eb e9 e7 ed ea ee f6 f7 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 ec ee ef ef fa f5 f1 f4 f6 fb f6 f7 f8 f8 ef f3 f4 ef ee ea ed e7 e6 df d7 d4 d4 db d4 d0 c3 c5 bb bd c1 ba c1 bb bc c4 bc b5 c2 c5 bc b7 c2 be bb b5 b5 b7 bd bf bb bc be be b8 b5 b8 b7 b5 a7 b1 a5 a4 a3 a2 a2 9d a1 95 95 96 95 8d 8c 82 77 7a 7c 76 76 73 80 78 79 76 78 74 71 71 6d 70 6a 67 6d 6b 78 6f 81 8e 7e 66 3b 24 10 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 02 06 05 08 1b 24 44 5f 73 8f a2 ab 8b 73 64 67 6c 6d 63 67 63 64 6b 6c 65 70 6e 64 65 74 6e 70 70 72 75 76 72 7a 79
 80 78 79 7e 7c 7c 79 83 83 8b 90 9e 98 a2 a4 ae b2 b0 ad b8 bc b8 bc c0 bd b0 b9 bf ba b9 bf b1 b7 b3 b3 bd bc b6 ba c8 cc d0 d6 d4 d1 d2 d3 d1 cd cf c9 ce d3 d9 da db dc d8 e0 e6 e5 e7 e6 e6 e5 f1 ed f6 f4 f4 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ef e5 e3 e4 df e7 e7 e9 e7 e3 f0 ec e9 e5 e2 dd e6 e3 e5 df d6 d3 c9 c7 d0 c7 c7 c6 c0 d0 d0 cf bd be c4 b5 bf af b5 b6 b8 b7 be b8 be bf b8 ba b8 be bd b6 bb bd bc bd bb b9 bb b8 b9 b3 ae b2 ac a5 a7 a9 a9 9e a2 a2 9e 9e 94 99 8f 8f 84 85 87 7a 7e 74 79 7d 81 7a 7d 77 75 73 70 71 6e 67 72 6a 6a 6e 6b 6d 6a 8c 8a 77 65 3a 1d 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 15 21 40 61 71 93 aa a0 8b 76 6d 6f 69 67 6a 65 63 66 64 6a 6c 6a 6e 71 6e 71 6d 70 6e 72 82 6f 75 7a 74 79 74 79 7a 7e 7c 85 89 8a 85 91 8e 9d 9a a5 af ae af b2 b5 bb b7 b7 af be bb b0 b7 b2 b3 b0 b9 b9 b2 b4 b6 b6 b1 b4 c5 cd ce d2 d7 ce d1 d2 cd c7 c9 c4 ce ce cd d5 d0 d9 d3 e0 e3 e2 e1 ea e6 f4 f6 f4 f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 e1 dd dc d5 dc e1 da da e0 d5 db df d9 db d7 d3 ca d2 cd c3 c6 bc c6 bb c3 bb bc bd c5 c6 be be c2 bf c0 bb c0 bb b3 bb ba b0 b4 ba c0 be b3 be ae b6 b9 b5 b5 b3 bd b9 bb bb bf bb b0 b3 a8 b1 b1 b2 af b1 aa 9e af 9a a5 99 9e 9c 96 99 89 84 82 83 7f 7e 7a 7e 75 7d 7d 76 73 78 7a 68 67 67 66 67 6d 6a 6a 6c 72 7b 84 7e 5f 37 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 04 06 05 0a 0f 1e 40 61 79 9c a5 95 7a 75 66 6f 6f 6d 68 65 65 67 67 61 65 68 6d 6e 65 6c 6c 6f 6f 6f 7a 72 6f 76 77 77 77 81 81 79 7f 7f 8b 93 88 8b 8f 94 92 a7 ad b5 b0 b2 b6 b7 b0 b5 ba b6 b8 b8 b5 b8 b9 b6 b5 b7 b3 b4 b9 ba b1 ba be c9 ce d4 c5 cf cb cd cb c7 c6 c4 c6 c6 d1 d6 d0 d1 cc d3 d9 dc e1 e2 ea f7 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef e6 d7 db da d9 d2 d4 c8 cc c9 cd d5 cc c8 cd c5 d1 bc bb bb b1 b7 ba c0 bf bd be bd bc bc bc bb c4 be b4 b5 b5 b5 ae ad b5 a7 ac b3 b1 bd af ae b6 b6 b0 b0 b9 b5 b3 b9 b7 b3 ba b9 b7 b8 af b7 b0 ad ae a3 a5 a8 a3 a9 ab 9a a5 95 93 91 93 8e 85 7c 85 82 85 87 7c 80 81 7d 75 77 75 76 6b 6a 6d 64 74 6e 6d 70 6b 82 88 75 5f 31 12 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0d 0f 1c 32 54 77 9a a4 8f 7d 75 72 73 70 69 68 69 6f 68 66 6a 62 64 67 66 70 71 6d 6f 76 72 79 6f 75 73 7c
 78 73 78 7c 7a 84 86 80 89 88 8e 90 99 9a 9e a5 a7 a6 b5 b5 b3 b0 af b0 b8 b7 bc b2 b8 b7 a7 b2 b7 b3 ab b6 ad b0 ad b9 cb c5 cb c5 cc c2 cf cc c9 c7 c9 c2 c7 c6 c8 ce c7 c9 c9 d4 d7 dd e6 e5 f3 f5 f9 ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e6 e3 d6 d7 cd c5 c2 c2 be bb c7 c0 c2 bf cb bf ba be b6 b2 b5 b6 af b6 b9 b8 b7 b5 bd bc ba b4 b9 b7 b8 b1 b5 b3 b2 ad af ad b0 b3 b3 af b1 b7 b0 a7 b1 b0 b5 ba b4 b1 bb ad b8 b2 b9 bf b3 ae aa aa ad a7 a3 a9 a4 a6 a3 a1 9a 96 90 8e 8a 8f 83 88 83 84 82 89 80 7e 82 7a 76 73 6c 6e 6e 6f 70 6a 6f 72 6b 62 6d 74 77 6a 4f 20 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 06 07 1f 33 4f 75 93 a1 8d 78 70 6c 75 73 69 69 69 64 68 69 66 63 6c 67 61 6d 6e 71 70 6e 6d 74 79 6b 75 79 77 74 7c 7b 7b 80 86 7f 85 82 91 93 91 9f a4 a5 a9 ab b1 b5 b3 ad b2 b5 b9 a9 b4 b5 b6 ae af b6 ac ae ab b5 b3 b0 ad b5 b9 b2 bb bd cd ca c9 c0 c9 c2 c1 c0 bb bf c1 c0 bf c2 c6 d2 d0 df e1 e3 e7 f1 ff ff ff ff ff f7 f3 f3 fc fa fe f5 f4 e5 eb ee f6 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ea e6 ea db d6 cb c1 bd bf b6 ba b9 bf bc bf b8 b2 b0 aa b7 b0 b2 b5 b3 b9 bf b0 b6 af ae b1 b4 b8 b3 af ae aa ac b2 ab b0 ab ac a9 b2 b2 aa ae b4 aa aa b1 b1 a9 ab b5 b0 b7 b0 b2 b4 b6 ae b6 b2 aa a7 a6 a3 a5 a1 a0 9a 9c 9a 92 8d 8b 8e 87 8b 8a 82 7b 82 81 7b 7f 76 6b 6f 70 77 6e 60 6b 69 6e 71 65 65 6b 5e 74 79 6a 4f 1d 0f 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0a 0c 19 36 48 6a 88 9f 8d 7a 71 71 69 79 74 70 71 6f 6a 69 6b 6a 69 6e 71 6d 6e 72 79 76 72 73 77 75 80 84 7e 7d 7a 80 85 82 7b 87 85 8b 91 98 96 9d a1 a9 b1 b1 a7 ab af b5 b3 b2 b7 b4 ae b2 af a8 b2 b2 af b0 b2 b5 ad a5 ac b0 bb b6 b7 b3 c6 d3 c4 c3 c4 b9 bc bb b9 b6 b5 c1 b3 ba bb bd c5 d1 d5 dc eb f6 ff ff ff f6 f3 e9 ec e0 e3 dc dc d2 cb c5 bf c3 cb cc dd e5 f6 ff ff ff ff ff ff ff ff ff ff ff ff f0 ea e3 dc d7 cc c0 b8 b4 ad b5 b0 b6 ac ae b6 af a4 ac ac b3 b0 b0 ac ba aa ad b4 b5 b0 a9 b1 a7 a9 ac aa ae a9 ae a4 ab ad a0 a7 a7 a4 ab b0 a9 b4 a4 a5 ad b2 af b0 b5 af b1 b0 b0 b7 af b0 a5 ac a7 ae ad 9f a1 99 9c 97 99 95 95 91 90 77 87 7f 80 85 7f 7d 7d 7a 78 75 6d 6d 71 6a 69 6c 74 71 72 68 64 6b 6c 6b 6e 5d 3c 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0d 18 19 34 4d 6a 88 94 84 7c 6f 77 7a 76 76 77 70 72 6b 71 72 6d 70 69 70 6f 69 77 7c 75 7d 84 7c 7f 7e 83
 83 84 86 84 87 84 84 85 90 92 96 97 9d 9e a3 a7 a7 ae ac b4 b1 b1 b4 ae ad b4 ae ab b0 a9 ab ad b0 b3 ae ae a4 aa ac a4 b3 ad b5 bb bd c5 c0 ae ba ac b6 bc b4 b3 b6 b1 b6 bb b7 bf c3 c4 cd d2 df f6 ff fe f1 e0 d9 d3 d1 d0 d0 c0 bc ac a2 a4 9a a0 a4 a9 b3 c6 d2 e2 ef ff ff ff ff ff ff ff ff ff ff f9 ed e6 e3 d4 cf c0 ad a5 ad a6 ad a7 ab af a6 ad b1 aa b8 af b1 ad ae b2 ae ad a8 b1 a2 aa a5 a7 aa ac a9 ab ac ae a6 9f a6 99 a7 ad ab a4 ac a7 ad a3 b1 a4 aa a7 ad a8 b1 b2 aa b7 b0 ac b1 a8 a2 a6 a0 a0 a0 a4 99 96 94 99 94 93 91 93 8b 8b 80 83 7e 81 80 75 7a 79 78 79 72 6d 71 6a 69 73 6c 6c 6b 74 67 61 64 64 5e 3b 1a 0e 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 05 0a 07 19 2e 46 6d 85 91 85 6d 70 6e 7a 76 79 81 71 70 70 6b 74 6b 68 6f 6c 6c 77 75 78 77 74 80 7b 81 82 84 7e 7c 81 84 87 87 87 87 7f 8b 8c 99 92 9f aa a5 aa ab a7 ae ad ad ae af b2 ab b2 b0 b0 b0 b1 ad b9 a8 a7 a5 a6 a5 a9 ad ab b3 ad b4 bd ca b2 b2 b3 b1 a6 b1 ad b4 a9 b6 b1 af b5 bd b8 cf c7 d2 e7 f6 fd eb d4 c6 c6 c3 bc b5 ad 9c 92 96 87 86 85 86 96 98 9d a2 ab c3 cf e3 f4 ff ff ff ff ff ff ff ff ff eb df dd d4 ce c0 b3 ac a6 9f a4 a4 a1 a8 aa b0 aa ad a9 ab ae ae ae b0 a7 aa ab a8 aa a9 a0 a5 a4 a6 ab 9f a8 a3 aa a8 a0 9b a2 a2 a5 a6 a5 ae a0 a0 9f ab ad a4 a5 a0 a7 ad ad b2 ac aa b0 a0 a1 9a a2 a2 9c a0 97 9d 95 8a 91 88 8a 8e 8c 87 87 82 7e 7e 77 6f 7d 73 78 6e 78 72 75 69 6d 69 6b 77 6c 6e 63 61 64 61 4a 26 24 0e 0c 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 12 17 3b 4e 6f 87 8f 79 72 73 77 77 84 76 79 73 7b 74 79 71 74 72 74 70 6e 72 71 7f 80 7a 85 80 89 85 82 8d 8a 83 89 88 8a 8d 8f 90 99 91 99 9c a0 a8 a5 b1 ae a4 b0 ac a6 ad ac b3 ad a8 b4 b0 b3 ae ae b1 a4 ab aa ad a4 ab aa a7 b2 a5 b2 bc b4 b6 ae a7 b0 ac b0 aa ab a9 ab a9 af b7 ac b3 bb bf c9 e9 f5 e3 d2 c6 b7 b0 b6 a3 94 8a 80 8a 89 84 75 6c 5f 87 8b 8b 93 9d a3 b8 c4 d2 dc f0 ff ff ff ff ff ff ff e5 e2 e0 ce d4 c9 b1 a8 9b 9e a1 a3 a5 9f a7 a2 a7 a4 b2 b3 af b2 aa a2 b4 a6 aa ac aa ae 9f a4 a7 9f a3 a5 aa a9 a5 a8 a2 a2 a2 a4 b0 a9 a4 ab 9d a2 a7 ab a7 aa ab a9 a9 aa ad a6 a4 a0 a5 a5 a1 9e 9e 9f 97 94 96 94 95 91 94 88 87 86 86 87 85 7f 7a 7b 7b 78 77 7d 7c 76 7b 75 71 6d 70 6e 70 6e 69 6d 65 65 66 5c 50 35 21 13 0a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 06 15 13 2c 56 69 81 87 76 79 71 75 77 7a 85 7a 76 7d 80 79 7f 76 76 7b 70 71 74 78 7f 7b 85 88 7f 8a 8e 87
 8f 8f 8e 8b 91 8c 90 92 8f 9f 95 99 a1 aa a7 ad a7 ae a6 ad aa af b1 af b3 aa ac b0 a8 a5 b1 b2 a5 ac a9 a9 ab a9 a3 a8 b0 a1 b0 b7 bc b9 a8 a7 ad af a3 a5 aa a5 a2 a9 a5 a4 af a7 b0 b8 be d5 ea ed db c0 aa 9e 99 90 89 7f 79 73 72 7c 7a 6c 63 48 73 7a 84 80 89 93 9c a6 a8 c0 c9 e0 ff ff ff ff ff ff e7 e5 e3 db cf c0 b0 9f 99 9d 9b 9e 98 a6 a1 ac af af ad b7 ad b6 af ab a9 ab a7 ab a8 a3 a0 9f a7 a1 a0 9e a4 a3 a5 a5 9e a2 a0 a5 a9 9d a5 a6 98 a0 a1 a3 a7 a7 a1 ab aa a7 a9 a7 a8 a5 a0 a0 9b 96 9f 92 91 8f 95 9d 8f 88 89 8a 8b 88 81 83 80 76 75 7e 7a 76 79 76 75 77 74 74 76 75 73 6f 72 6e 6f 64 6b 55 63 52 49 34 27 12 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 0e 09 1b 2c 54 67 85 8e 72 72 6e 71 80 7b 85 80 7e 7d 7b 84 81 7c 7c 76 77 78 72 77 73 7e 83 7e 86 80 8b 85 90 91 97 8e 8c 8f 94 96 9c a0 9a a2 a8 a3 a8 ab a4 ab a8 a8 a2 ac ad b1 ad a9 ac a9 a5 a5 af a9 af a9 a3 ac a7 a7 a8 a5 a5 af ae ba b9 b5 ac ae ac a9 a3 a6 a0 a1 a8 a7 aa 9d ad ac ae b7 b7 cf e6 e1 bf b4 98 81 77 6d 73 6e 6f 75 72 69 66 66 5f 5e 6c 6b 6c 6f 78 84 91 9e 9a a5 b1 c2 ce fb ff ff ff ff e4 e0 dd d9 d1 c9 ad a5 8e 98 9b 9f 9a a1 9e a5 a9 ad a6 aa b4 ac ab af a4 a4 a7 9d a1 a1 9d a3 a8 a1 9e a0 9e 9a a0 a0 a0 9e a1 a1 9b a1 9a 9d a0 9e 96 9f 9b 9f a4 a4 9a 9a 97 a9 9e 9f a2 94 94 93 90 95 95 93 91 92 81 83 85 7f 89 81 7f 89 77 79 7e 75 77 79 76 78 7d 73 84 75 79 74 72 7b 67 6d 70 67 5c 58 61 55 54 41 29 1d 17 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0b 14 21 35 4e 6d 82 8a 7e 6e 71 6f 7e 7d 84 86 84 80 82 7e 84 7f 7e 82 76 7c 7b 80 86 85 8a 8b 87 8c 8e 90 90 8e 91 95 93 9b 99 9a 9a 99 a0 9e a3 a6 a7 a5 a7 a6 b0 b2 a9 aa af a7 b8 ac ad ae ac aa a5 ac a5 a6 ae a5 ac a6 a2 a9 ab af bd c0 bf ae ab aa a8 a1 a6 a6 a5 a3 a4 9c a3 af a8 ad a8 b3 c5 d8 d7 cf b1 98 7f 70 63 61 5e 67 6b 70 6a 65 66 66 60 5b 66 6a 74 70 71 7b 87 8e 8a 98 9b a9 ba d3 fe ff ff ff f3 e5 dc db d3 cb b3 a8 97 92 92 94 a1 a1 a0 a1 a4 ac ab b5 ae ab a1 ab b0 a1 a7 a4 a0 9d 96 9e 97 a3 9d a1 9e 9a 9e a1 a3 93 97 a1 9b 95 9e 98 90 98 a4 97 a3 a5 a0 9d 97 9d a6 99 9b 93 92 94 93 94 94 92 87 8d 90 90 8d 83 8d 7d 86 81 85 7e 7a 7e 7d 84 7d 80 73 75 79 7e 7d 79 75 70 79 72 6c 71 65 6c 64 5f 63 59 58 4b 34 24 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0c 18 27 3e 4b 75 8a 91 80 71 77 72 76 84 83 85 85 88 8b 8d 8d 84 87 83 80 81 82 83 83 89 91 8d 99 8a 90 96
 94 95 97 9a a0 90 a0 99 9f 9f a1 a2 a1 aa 9d a7 a7 aa b4 aa ac b3 b4 a7 ae ad aa aa ab b3 a7 ae a9 a6 a6 ad a7 a9 af ae b3 b4 c1 bd b8 ae ac a9 af a2 aa a7 a5 ad a6 b0 ac aa af b0 a4 af c4 d9 d0 bc a1 7a 69 5a 5a 53 5c 60 60 58 51 51 4b 59 5a 50 56 66 6b 75 7c 7b 80 7d 76 8a 91 8c a7 b7 db ff ff ff f9 e3 e1 e1 d8 ce b9 ad 9d 93 96 98 9d a0 9b 9e ae b1 af b0 ab ad aa ad a9 a8 a7 a3 a6 9b a3 9d 9e 9d a2 9e 9e a0 9e 9d 9b 9a 9a 9f 9f a1 9d a1 98 95 a2 9a a2 9c 94 9a 97 a4 a0 a0 9e 96 96 94 92 8b 91 92 82 97 8a 8b 8b 89 7d 84 81 88 81 81 7d 7e 78 71 75 7c 7a 7b 7a 76 82 75 74 6f 71 71 70 6b 70 6e 6a 61 5d 68 5e 4f 39 27 17 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 13 28 34 50 75 84 8d 7c 6e 6e 73 73 78 7c 7c 78 7d 8a 8d 97 8c 87 81 81 82 81 84 87 82 92 8f 8a 96 90 94 96 99 a0 98 96 9c 99 9d a9 9e a7 a5 a2 a0 9e ac a3 aa a7 a7 a4 ad af a7 ac a6 ad a7 b3 a7 a1 a7 aa a6 a7 a4 aa 9f 9e af b1 b8 c1 bf ba a6 ad ac a4 a4 a5 a9 a0 ad a4 9e a7 a6 a9 a6 b2 b9 c9 ce c3 a7 85 6c 55 4d 4a 52 65 59 4a 41 34 3e 40 3d 44 42 42 52 5f 66 76 7e 81 79 79 75 7b 89 8c a5 c1 e8 ff ff fe ef ed e2 d6 cf be b1 9d 95 8f 94 91 9d 9e a0 aa a4 ae b4 b3 ab a7 aa a6 a4 a6 a4 a3 a0 a2 95 96 a0 a1 9d 94 98 99 90 90 99 92 9b 99 96 90 99 90 93 99 95 97 99 9a 99 9a 95 9f 94 96 96 8e 8b 8d 8f 8d 82 8b 88 8e 8d 7e 87 78 84 84 7e 87 7a 76 7a 78 7c 7a 7a 82 82 7d 78 75 7b 75 72 6f 72 6e 6a 6a 64 67 61 72 69 59 4d 32 28 1c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 06 13 1a 31 46 5b 7c 8a 91 81 74 75 70 74 7c 7a 8a 7f 85 8a 8b 8e 87 91 8c 88 8b 8e 8f 8e 8a 92 92 95 99 99 94 99 9b 9a 97 a3 a0 9a 9d a2 a3 a5 a4 9e a1 a1 a5 a6 a5 a9 aa a7 ac b2 b0 a9 a6 a8 aa a2 a2 a7 af ae a8 a9 aa a7 a9 a6 ba b8 ba b5 ba aa ac ad aa ad a1 a5 ac a8 a5 a0 ac a8 ae af b1 b2 b7 c3 bd a8 89 68 5e 4b 4e 5f 60 59 44 2f 2f 2a 2f 33 39 33 32 36 3c 44 47 61 6b 6e 70 63 66 77 86 86 92 b1 d0 fe ff ff f0 ea e4 d3 d0 be b0 97 9e 93 93 94 95 9c a9 a4 aa a8 ac ac ab aa a7 a7 a2 a8 a5 9d a0 98 93 99 97 98 9e 93 94 9b 94 96 94 98 99 9f 90 92 9a 8e 8c 94 94 9b 97 90 95 8a 96 8f 95 92 8e 92 8b 88 86 88 85 85 82 81 84 84 81 82 81 88 83 82 7a 7a 75 76 76 79 81 79 7f 76 71 7a 79 75 6d 76 69 64 6d 63 6c 68 69 72 75 68 52 43 2d 20 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 1e 22 2b 4a 65 77 98 8f 82 78 77 71 78 7d 7b 81 8b 8c 91 94 92 8b 94 90 8e 85 93 92 92 92 94 99 97 94 9b 9e
 9a a0 9d 9c a4 9d a2 aa a1 aa a8 a3 a5 a9 b0 af ab a4 ad ab ad a6 a6 aa a9 a6 ad a6 9e aa a2 aa a9 a1 a5 a8 a7 ac b0 b6 b8 b6 b5 b8 b5 ae a4 a5 ac ac ab a9 a9 a6 a8 a5 ae ae b0 b5 b2 c1 c1 b6 9c 7b 64 52 52 52 51 4d 46 32 28 2a 24 2e 34 26 27 2f 30 33 3c 39 42 43 59 56 61 6d 7d 87 83 8d a0 c0 f2 ff ff f7 e6 e1 cb c7 b4 b3 99 9d 97 8d 9c 99 a1 a0 ab ab aa b1 aa a3 a7 ab a0 a2 9d 9c 97 9b 9e 97 91 99 97 a1 96 96 91 94 93 93 9b 95 9f 8f 8e 90 88 96 8a 8e 90 94 95 8f 8d 95 8f 93 8d 8f 8a 91 81 89 89 8d 87 8a 81 86 7c 81 85 83 7a 79 83 87 7c 7a 7a 7a 81 7f 7d 7b 83 78 80 71 6e 6f 6f 7a 6c 6b 63 6e 73 71 7a 75 6d 55 51 31 23 19 0b 05 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 1b 26 2d 4e 66 87 9b 97 7f 79 73 74 7a 7b 78 84 89 8c 91 99 97 8b 92 92 92 95 98 99 8c 8a 98 92 99 9e 9c 99 a2 9b a9 9a a3 a1 a9 a5 a0 a4 a0 a4 aa a9 a7 ac a6 a3 b0 ad af a6 ab a4 a9 a9 ad a4 a8 a4 a7 b4 ad ae a1 b1 b3 b1 b2 b6 b6 b8 b1 b6 a9 b1 af b5 b0 ad af b1 a9 a5 ad af ae b1 b1 b5 b6 c2 bb a3 8b 6e 57 4f 47 45 33 34 2b 29 23 23 2c 24 2d 2d 2a 29 2b 2b 2b 34 35 38 41 3b 51 6a 7a 82 8c 8b 9f b7 de ff ff ed f0 dc cb c7 af ab 9f 8d 91 96 9a a2 9d a6 a4 aa b3 ac a9 a4 a1 a8 a0 a5 9c 9d 9c 98 95 98 9a 96 8e 91 97 90 95 95 8f 90 98 8f 8e 8e 91 94 8c 90 94 91 90 92 91 8c 94 8d 89 8f 8d 91 8d 87 87 83 85 7c 81 82 80 87 7d 7f 78 80 76 7b 83 7a 77 7c 7c 7c 7b 7b 7a 80 7a 71 76 76 72 6d 70 70 70 6b 6a 6f 70 72 7a 6e 6a 5d 4b 40 28 1a 0d 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 11 14 21 23 35 4c 69 80 92 9a 7c 77 79 76 7c 83 7b 84 7e 87 8d 8f 93 92 90 8f 90 8f 96 94 95 9a 8e 99 9b 9d 9e 9f 9c 9f a1 9e a5 ae a9 ac a8 aa a7 a5 aa a9 aa a9 a3 ad a5 b0 a1 ad af ad b4 ad a1 a5 a4 a9 a3 a0 ac af a7 a8 a9 af b6 af b9 b9 b4 ac b1 ae ae b0 b6 b1 ad a5 a9 ac ac af b0 ae b3 b6 b8 b6 bd 9f 71 5a 50 49 3b 30 25 29 27 27 24 25 24 21 1d 28 25 28 2b 28 2f 2e 2d 30 35 3e 47 50 60 70 84 95 a3 ca ff ff ff ef ec e4 cc bb a7 9e 94 90 8d 94 95 9a a6 ac 9a a7 ab a8 aa a1 a3 9b a1 95 97 9b 9a 98 94 97 9a 96 96 94 93 99 92 90 90 93 97 94 94 90 8c 88 87 90 8b 8c 8c 86 8d 93 8c 8e 8c 8b 86 86 81 89 7f 81 8a 86 7d 78 78 83 82 87 7d 7a 78 7e 7d 7c 7b 72 7e 7f 7c 78 7c 78 75 77 71 75 68 70 71 6c 6d 69 74 6d 74 67 79 75 66 61 45 3d 28 1f 15 0f 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0e 1a 26 30 46 5c 6e 80 9e 97 85 82 75 83 78 81 82 84 8d 8f 91 90 94 9a 95 97 8e 90 8e 96 9a 9e 9f a3 a2 a1 9e 9f
 a9 a5 a1 aa 9d a5 af a8 a9 a6 a7 ac a8 a9 a7 ac b0 aa ac ab aa aa b6 ad ae a5 a3 a5 ae a5 a5 a9 b1 ae b3 ba ba ae b2 ad bb b0 b2 ad ad b1 ad af b8 ab b1 ae b4 a6 b2 b7 ab ad b2 b7 be c4 ae 8d 5b 4b 3b 2a 2c 23 25 23 1d 20 1e 19 1c 1e 20 24 18 15 21 22 26 2d 26 34 36 35 39 3c 48 5f 7b a8 cb f1 ff ff fc e9 dd d6 c5 bb a4 9b 92 97 95 96 9c 91 9b a2 af a3 ae a7 aa a5 9c a2 a3 9e 99 a4 96 9b 9e 97 94 91 95 8d 92 8b 90 8a 92 90 92 90 8e 91 94 94 91 88 8a 85 8e 8d 82 90 89 8a 7e 85 89 88 85 83 7d 85 82 7a 7c 80 82 85 7a 7e 80 7d 89 7b 82 7d 79 82 81 7b 80 79 77 7a 7e 79 7a 6c 6b 70 75 6b 6a 6c 71 6a 70 6e 76 7b 6e 68 59 44 39 29 1b 10 06 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 06 0b 0a 24 21 38 4a 57 73 8f a1 97 8b 7c 76 7f 83 7c 83 89 7f 8c 90 96 95 98 94 9b 98 9e 93 9b 96 91 9b a0 9f a1 9e a4 a9 a9 a9 a7 a3 a6 a4 ac a6 ab af a8 a5 af a8 ae b3 ae b1 a7 ac a8 b0 a5 b0 aa a5 ac a2 a8 ad b2 b1 b3 b1 ae b3 aa b4 b7 b8 b4 af af b3 b0 af b1 b3 ac ad ad ae b2 b0 b4 b1 b5 be c3 b9 b9 a5 84 51 3b 29 1c 27 1f 2a 1e 1b 19 17 10 15 1a 15 14 17 1b 1c 22 20 1f 25 2c 34 2c 3a 35 42 51 75 98 b3 ed ff ff df dc c8 c6 b6 b8 a0 99 93 93 90 8f 98 9f a1 aa a7 a9 aa a8 a7 9c 9d 9e 97 98 8c 9f 94 99 97 8f 98 99 95 95 8c 93 8f 8f 89 8b 8e 8f 90 8a 8e 8d 8b 89 8b 84 7e 82 84 8d 7d 82 7e 81 7d 7d 81 7c 7a 7c 7c 7d 7f 7f 79 7c 7b 74 7e 7a 81 75 75 82 73 7a 80 7c 78 76 76 75 6d 6e 6f 6e 71 69 70 65 68 71 74 6c 6d 67 7b 70 6f 67 56 48 33 2b 15 13 07 0e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 11 13 19 23 3b 44 5b 80 91 a6 99 7e 80 7d 80 85 83 8c 7f 89 90 8f 94 93 96 94 91 90 94 93 9a 97 9d a1 a2 9b a4 a4 a7 aa a1 a9 a4 a3 a1 9a ae ae a9 a0 a9 a7 a6 ab a9 b0 ac ad af a9 af af b4 b2 b3 a4 ae ab ae b5 b3 ae b1 ae b8 b2 b3 ad b2 b7 ab b4 b3 ae b5 b2 b6 ad ae ac b3 b4 b1 ae bc b8 bd bb c7 c5 c2 ae 75 49 2b 14 21 13 1b 1d 22 0f 16 0c 12 0c 14 15 14 11 15 0e 14 1a 14 1d 26 25 2f 32 30 35 48 5d 7a a3 df ff f6 d6 c8 bb bf b2 aa 97 95 8f 95 8c 90 93 a4 a1 a7 a3 a6 aa a9 a7 9d 9d 9e 9f 9b 97 98 92 90 95 90 92 8b 8d 8c 8e 8d 85 91 90 89 8b 7e 8c 85 89 84 8b 8c 8a 81 7a 8a 84 82 7b 80 82 7f 81 74 81 7f 78 7a 78 7a 76 78 78 74 74 7f 7c 77 7e 7b 82 7b 7f 7b 81 75 7c 72 76 71 6b 6f 67 65 68 65 6b 71 71 73 70 6a 64 6f 76 76 70 63 5b 4e 47 38 23 19 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 0d 1e 24 2e 3c 47 60 7b 90 b1 a0 86 7f 72 7f 80 8f 8f 8a 8d 8a 85 8e 8d 91 95 8f 9b 94 95 94 9d 97 9a a1 9d a3 9d a5
 a3 a0 a0 a7 a5 a4 ac a7 a4 ab aa aa aa a7 a8 ae a6 9f a6 af a8 af b5 a3 b1 ab af ab b0 a7 ac b3 b1 b0 b2 ac af b3 b3 b9 b5 b0 b5 b6 b1 c0 b2 b5 b8 ad b0 b5 ac b3 b1 b6 b5 c3 c7 c5 c3 bf a2 6a 2f 22 1f 14 1a 1e 16 14 1a 10 12 0d 0b 12 0f 0a 0e 15 0d 10 15 1c 1c 1f 1c 1c 2b 3a 35 44 52 69 93 cd f0 e0 bd b0 b0 af b2 a5 96 98 98 94 95 95 97 9f 9f a8 9f a2 a2 a6 a1 a0 a5 94 9b 9b 95 9a 91 90 86 8b 91 94 91 8c 89 89 90 8b 88 8b 8c 8e 94 80 8b 8e 85 8a 85 89 85 83 86 84 7b 80 7c 7d 80 79 7e 73 71 75 7f 7f 77 77 71 7b 79 78 7a 7a 7e 79 79 84 79 77 76 71 78 71 6d 66 6a 60 73 6a 6e 6c 70 6c 70 7a 76 64 64 67 73 79 71 6f 66 53 49 36 36 20 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 10 08 19 2e 27 3e 54 68 80 96 a5 a2 87 7f 7a 76 7e 84 85 84 87 8d 87 93 86 86 92 8e 8b 91 92 94 a0 9e 9f a1 9f 9b 9e a9 a6 aa a6 a1 a7 a8 a9 9d b4 a9 9e a5 ac a6 aa af a2 a7 a9 ad ab ab ae ac b0 a7 a4 aa ac ad ae ae af b0 a8 b5 b5 b6 b2 b0 b8 c0 b5 ba ba b6 ae b4 b5 ad b1 ad b3 b7 b2 bc c0 bd c6 c6 c7 c1 a1 65 36 22 11 18 0f 0e 15 14 0b 10 0b 0e 05 10 06 10 0d 09 0d 0d 0e 0c 0b 0c 15 1a 22 2e 3a 3a 4a 61 89 be d6 d3 ad a8 a0 9f a0 99 95 9a 8e 96 95 9d 9b a2 9e 99 9d 9f 99 a2 9c a1 9c a0 94 90 99 94 95 92 8e 8f 8f 87 89 80 86 81 81 89 85 8d 8b 83 88 82 8b 84 78 7a 88 87 84 7f 77 80 80 70 76 7f 7b 7a 74 75 72 75 75 79 7a 6f 78 77 75 79 7e 7a 7a 7b 7e 7b 7a 7e 7c 6d 6e 74 69 72 70 65 71 71 69 6b 64 75 73 7a 70 65 66 6a 76 77 6b 6d 62 57 49 41 2e 23 1b 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 1c 22 29 3c 44 57 6f 81 97 a1 9e 84 82 74 7d 7f 78 88 8b 88 8d 82 92 88 89 87 8f 91 8f 93 95 90 97 9a 9d 9a 9b 9e 9a a2 a2 99 a5 a8 a1 9f 9f a3 a5 a0 a4 a4 a5 a6 a3 a3 af a5 ab aa aa b1 ab ae a6 a7 a8 a7 a8 ad aa b0 ae b1 b9 ac b6 b8 b5 b8 b7 b0 b9 b6 b8 b4 b7 b7 b5 b1 b6 ac b0 ba c0 d0 c7 ca c5 c5 bf 9c 51 2f 22 10 0e 0f 15 14 0a 05 00 08 05 03 00 06 05 06 02 06 0a 0d 0b 0f 0f 12 1f 16 2e 2d 37 41 4e 80 b3 d6 be 9f 9d 95 9f a1 9e 95 94 91 97 98 95 96 a0 9b a3 9e 9c a5 9e 95 9c 9f 9b 94 98 95 94 92 94 91 92 8e 8e 89 86 8b 83 82 88 85 80 81 82 8d 7c 85 84 7d 7c 81 80 7e 7f 76 77 78 73 7a 7b 6c 6b 71 76 73 70 75 6f 6e 72 71 70 6b 73 76 74 7a 6b 77 7d 78 70 6d 68 74 64 6f 74 69 68 67 6b 62 6d 6a 6b 7c 70 68 5b 59 6c 72 82 70 6f 63 5a 5b 41 33 25 15 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 15 11 1d 29 35 4b 5e 74 8e a8 a8 9a 7b 82 7a 85 7b 81 87 7f 88 87 89 8a 8b 8a 8a 8c 86 8b 96 8d 94 9b 99 96 a0 96 a2 9d
 9f a1 9c 9f a6 aa a1 a9 a3 9d a7 a5 a5 a4 a4 a5 a0 a6 ac a0 aa af ad a8 a6 a9 a7 ab af b0 ae ad ae b8 b6 b6 b3 b6 b4 b5 b7 bb b5 b9 be b5 ac b7 ba b3 b5 b9 b0 b9 be be c5 be cd c9 c5 ba 98 53 37 1f 0f 20 0e 0a 12 07 05 06 09 09 03 05 06 05 04 00 06 06 0d 0b 0b 08 13 1f 1a 20 1f 3e 47 46 6e a2 d6 b7 94 95 8b 96 9b 9f 9b 95 96 9c 9b 9c 97 9c 91 9b 94 a0 9c 9f 9e 9a 98 9d 94 95 8f 93 93 94 92 8e 8f 89 90 88 8c 84 81 84 84 82 85 83 89 7e 7b 89 86 7e 7a 7b 7e 76 84 7f 70 72 73 7d 6f 74 72 6b 6e 75 75 6e 71 76 77 72 71 6e 75 7b 72 7f 73 7b 74 69 6e 64 72 6f 72 68 69 69 70 65 6d 6d 78 79 72 72 66 57 5b 62 70 7f 77 71 6c 5a 4b 46 36 25 16 19 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 06 0a 0c 11 1c 33 41 4e 5d 77 89 a0 b4 98 85 7b 72 7d 83 81 86 7b 81 8d 85 8b 88 84 8a 86 88 8f 88 8a 9a 8f 9a 97 92 96 9d 9d 9a a1 9c a1 a4 9b 9d a1 aa a4 a3 a6 a3 9d a2 a5 9f a9 a5 ae a5 a5 a9 a5 aa a1 ae a9 a4 b0 ad b0 b7 b2 b6 bd b7 bf ba bc be b6 b1 bb b1 bb b8 b4 b1 ad b2 bd b6 bc c5 c3 c3 cb cb c8 c3 bb 95 5e 35 1a 0e 10 05 03 0a 10 0a 01 07 05 03 03 06 06 03 00 06 0a 03 06 06 0a 12 18 1c 14 22 29 42 47 64 a6 be a7 93 93 9c 9b 9f a0 9b 97 96 9c 94 96 97 9f 96 9d 98 9c a4 9c 9c 99 98 a1 90 99 97 93 8b 94 8d 85 90 88 8d 87 83 85 85 86 8a 84 86 7e 85 7e 81 81 7a 7a 7f 81 78 79 7a 77 75 74 76 74 6d 6c 72 74 70 6b 66 70 6d 74 71 73 6f 7d 6f 7a 75 70 76 72 6f 68 68 66 6c 6e 64 6b 6b 67 71 63 68 6c 72 7b 76 69 63 5f 5a 5f 6d 7c 7d 77 66 68 5f 50 3e 33 1f 19 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 0f 19 2d 33 3e 51 64 7e 96 a4 a5 97 7b 79 79 72 88 83 7e 84 83 8c 8e 8e 8e 87 8d 88 85 86 8e 99 89 95 95 95 8c 91 a1 9d 9b a0 a2 9a 9d 9e 9f 97 a4 a0 9b 9d 9e a2 a2 9e a3 9f a6 a5 a5 a9 9d a6 a9 ac a9 aa a4 a0 ac af b8 b6 b3 bf b7 b3 be b9 b7 b8 b1 b0 ba aa b5 bb b8 b8 b8 ba b9 be bf c4 c3 ca cd c9 c6 bb 9c 5a 2f 18 08 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 06 0a 0f 10 19 22 3a 44 5b 94 ad a0 93 90 8c 97 9e 9f 9e 99 92 8f 93 99 98 94 99 99 90 98 94 96 98 93 97 94 94 96 90 94 89 8d 87 86 83 8c 80 84 84 81 7c 79 7b 79 7b 83 77 7d 7d 83 77 7b 82 73 73 75 6e 74 6e 6f 71 70 6c 6c 71 65 65 6d 6a 70 76 6e 72 75 71 78 6f 74 71 76 6c 6c 63 64 67 66 6a 70 6d 65 67 6c 6b 70 71 74 74 77 6a 65 62 5b 55 5d 75 78 77 76 69 61 54 55 41 33 23 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 10 15 22 31 40 55 67 83 9c a3 a7 90 6f 70 71 79 81 7e 85 88 89 8b 88 8d 8e 8b 8d 85 84 88 8a 8f 89 8e 88 98 96 96 a4 93
 97 9a 99 92 a3 95 9f 9e a0 aa 96 9c a8 a2 a2 9a 9d a3 a1 a4 a2 9c a4 9d a6 a5 aa b4 ab b2 b1 ae ba b7 bb be bb bb bb b3 c1 b9 b9 b8 ba b3 b1 b0 b5 bc b7 bb bd b7 bb c7 cc c9 d6 c7 c0 b6 a2 71 38 16 06 05 0a 04 0f 07 08 00 06 05 03 05 06 05 03 00 06 06 03 00 06 05 11 0e 08 1b 14 22 3d 50 66 8f a1 94 95 90 8e 92 a2 9a 9a 97 94 96 9d 8b 97 97 9a 91 96 8f 94 9a 97 9f 96 96 9b 8a 8b 91 90 84 8c 89 85 83 82 84 89 84 83 7d 83 7e 76 7f 79 7b 82 7f 7c 75 78 7f 77 6f 71 6f 6e 6e 74 65 75 6b 66 67 62 68 69 71 70 70 6d 6c 6b 6b 74 6c 70 6a 6a 74 68 69 67 5e 6c 66 6e 6b 6e 73 6f 73 6f 6f 78 6f 66 5e 5b 57 56 5a 6d 7b 75 72 72 62 5f 59 4a 33 21 20 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 13 16 28 34 47 56 6f 7f 98 a4 a6 8d 7b 76 74 6f 7b 7a 89 8d 87 8e 8d 8c 91 87 81 89 8c 86 90 90 96 8e 8e 95 91 90 98 96 99 9e 99 99 96 9d 95 97 9f 9c 9f 9d 9e 9f 9f 9c a2 a3 a7 9e 9f 9f 99 a5 a3 a3 ac ab b0 ae b2 b5 b9 ba be c0 b9 bb bc bb bc b0 bc ba b0 b4 b5 b2 b9 a9 bd b8 ca c4 c4 c6 ce cb cc c5 c0 bc ad 84 36 1c 07 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 0a 0d 0b 0c 15 16 30 48 61 91 99 94 99 90 95 98 96 9f 9d 94 8d 94 95 8d 90 96 89 9a 8e 91 96 91 9a 9c 92 98 90 98 8f 8f 8c 8a 8f 8b 86 88 85 86 7f 7f 83 7d 85 7e 79 7e 81 79 7c 80 70 6d 7b 74 71 73 6d 6d 71 6e 6c 76 71 6c 6d 68 6b 64 6d 6f 6b 72 6f 67 73 7b 6b 72 68 6e 5f 65 61 69 6b 66 66 6a 78 74 6d 6e 6f 6b 72 6f 70 5f 5e 5d 55 54 57 68 6a 7f 7d 76 71 65 60 52 51 3d 2b 22 10 06 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 13 22 29 37 52 54 69 79 92 a5 9f 84 7c 73 72 78 7b 7a 7d 8c 85 80 8e 8b 89 91 8a 87 88 89 87 89 8b 8c 91 95 95 8a 91 97 95 91 94 99 93 99 93 9b 96 99 9c 9c 99 9d a0 9b a1 9b 97 9e 9c a3 9e 98 a1 a0 a4 a7 a8 b2 b7 ba ba b4 b9 b9 bd b6 b3 b4 bb ab b4 b4 aa b3 af b5 ba b4 b3 bd bd c0 c6 c6 ca c8 cd c3 bb b1 a5 7f 2e 11 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 0a 0d 06 14 16 2a 50 72 8b 93 94 96 8b 98 8c 9b 90 8b 8a 84 90 8e 8e 91 90 91 87 8e 8c 8e 98 90 8d 8e 8b 91 90 8e 91 88 83 86 85 81 7e 83 83 7d 75 80 80 7b 7d 80 75 7e 77 71 7d 74 78 78 75 71 6d 6e 70 66 76 69 69 6d 65 6b 64 5e 68 65 70 6a 6e 70 74 70 73 6a 65 66 64 66 61 62 66 62 60 63 67 6d 73 6b 70 6b 69 64 6a 69 5d 57 58 55 52 50 5f 66 7b 79 70 76 6a 61 5c 54 44 2b 1d 15 07 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0d 16 26 3a 4e 54 66 7f 9a a0 ad 8d 79 76 6c 72 80 78 7e 80 83 82 8c 88 98 90 87 89 89 8e 87 8d 87 8a 86 8d 8b 97 96 8e
 92 97 97 94 9c 8f 97 90 94 9d 92 95 9c 96 94 9c 9b 98 a2 9a a7 a0 9d 9c a3 a6 a5 b0 aa b6 bc bf bb b8 ba be bb b5 b4 b9 b7 b6 b2 b2 b1 aa a9 aa b1 ba b5 b5 b7 c3 bc c4 c3 c4 ce c1 b4 b7 9f 77 29 0f 06 05 0e 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 0d 0d 0f 10 18 2f 55 7c 98 98 93 91 92 8f 94 8d 87 85 8e 87 96 8c 8b 8c 88 8b 91 8a 83 8d 87 91 94 90 94 92 8b 88 8c 8f 83 8b 88 7e 84 85 78 81 7f 82 75 7b 74 77 75 7a 75 7a 7b 76 70 71 71 6d 6e 66 72 71 70 68 70 69 6f 68 62 61 67 66 63 69 6d 6e 70 68 70 67 65 65 63 60 65 62 62 63 68 6d 67 75 72 70 6c 68 63 68 60 61 58 56 5a 55 55 54 58 69 7a 7a 78 6e 6f 5f 58 4e 3d 2e 21 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 13 1e 2e 45 47 5f 6a 84 9b aa a3 8c 71 70 6d 71 7b 76 7c 83 88 80 85 8d 8d 8a 85 89 83 87 96 8a 87 93 90 95 91 95 96 97 91 91 95 8f 96 94 8f 93 91 94 98 93 98 93 97 98 a0 99 98 9b 94 a0 9e 9f a3 a5 a7 af b0 aa b1 b8 b5 af b9 ba b6 b0 b5 b2 b8 bf b8 b6 ae b0 a4 a9 b0 af b8 b5 b8 be bc c3 cc bd c5 bd b8 af a0 84 3e 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 10 0d 18 0e 0c 26 4a 7a 99 93 9a 91 8f 89 88 92 8f 89 83 86 8c 89 84 8b 91 92 91 8c 86 8c 92 8c 8f 89 8b 8e 8f 96 86 88 89 85 89 79 83 7f 81 82 7b 81 7c 77 79 79 7d 7a 76 79 7c 74 76 75 77 6a 6a 77 6b 6e 66 6b 66 6d 6f 67 68 69 69 71 6a 67 6f 74 6c 69 6a 63 64 67 61 62 64 65 67 68 6b 72 70 75 79 6e 68 66 62 63 62 60 5e 51 55 55 4d 4f 52 60 71 7e 78 69 6d 63 51 4d 41 31 28 15 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 0f 21 29 41 53 60 76 83 9c a9 9f 92 74 77 70 77 7a 77 7b 80 7e 7f 89 87 8a 8c 89 82 84 85 89 8f 8c 8f 90 92 8a 90 93 8f 8a 99 8d 88 92 96 8b 92 96 98 8b 8d 92 94 92 94 9a 90 90 9b 9b 9b 9b a3 a3 a1 a5 ac ae b2 b5 af b3 b9 b4 b9 b3 ae ac b2 b0 af ab aa aa a0 aa a5 b0 ab a9 a0 b0 b9 b1 b9 c0 b6 ba b6 a6 ab a6 8f 31 08 06 05 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 08 0c 0a 0e 0c 12 18 4e 83 94 96 9a 8c 87 8a 8c 88 8a 87 8c 8a 8f 8a 88 8b 8b 88 87 88 8e 8e 8d 95 91 89 8a 86 8b 8b 88 8b 8a 83 81 86 81 81 7e 79 81 77 7b 7a 74 7c 76 74 6b 70 7b 73 75 75 64 66 69 6b 70 5f 65 65 67 5e 70 60 66 60 61 6e 6a 69 6b 70 6b 64 64 58 64 5e 66 61 63 66 66 6e 6e 6f 6c 71 72 67 63 5d 62 62 60 5c 5e 4e 4e 51 4e 51 4f 63 71 78 75 6e 74 65 61 51 43 33 29 16 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0a 1d 23 2f 44 45 5f 73 8b 98 a7 a9 91 7b 72 70 75 75 74 74 71 7b 86 8b 87 8a 85 85 84 8c 89 8c 8c 8b 8c 90 8e 8e 8d 86 91
 8c 89 8f 8b 88 8d 8a 8e 90 8f 8e 89 91 92 93 98 97 8b 91 9e 94 9f 9d 94 a7 9b a9 a3 ad ae ad af b6 b1 b2 b2 a7 a8 b2 a6 a5 b0 aa af a2 a6 a0 97 a7 a3 a8 ae b3 b4 b5 b1 ae b0 b0 ad ae a2 a2 89 40 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 07 06 07 05 10 1e 4b 81 87 92 89 89 88 87 84 8d 87 7e 83 86 8e 80 80 81 82 8d 89 8d 83 8f 91 8b 82 8b 94 89 8d 7d 8c 83 86 83 7f 89 78 7b 7b 7d 80 7b 80 78 79 71 7c 73 73 76 73 71 67 6c 6c 6b 71 63 6d 67 6c 66 6e 68 60 68 65 63 66 6c 69 70 69 62 67 5c 66 63 63 63 61 66 5f 6e 5e 66 72 6a 63 6f 63 55 60 67 58 5e 5d 5a 57 4f 5a 55 4c 4a 4f 58 70 79 79 70 6b 67 62 55 4a 3a 2e 16 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1e 1f 3a 48 52 5a 6e 8a 95 aa a1 90 7c 6e 76 71 6f 71 75 78 72 7b 86 84 87 89 86 86 84 89 8b 89 89 89 8e 8a 86 8e 8e 8a 8b 8c 8c 87 90 91 95 8b 8f 8e 8f 8f 8f 91 87 8c 92 9d 99 99 94 97 97 a4 9f a4 aa a5 a6 af ac b1 ac b0 b4 b2 af af ab a7 a8 a4 ab a5 a5 a4 99 9c a3 9b 9f a4 a9 af a7 ab ae af ac a9 a5 9d 98 88 41 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 0a 0c 08 07 18 44 78 87 8d 89 8b 8c 7e 7f 84 84 82 81 81 8c 85 86 87 83 84 8c 81 89 88 89 8c 85 87 87 86 86 85 8f 87 82 85 7e 82 82 83 79 79 7a 74 79 77 7b 76 7b 79 73 76 70 6c 70 71 65 6e 63 72 66 65 6b 66 66 62 66 6b 6a 6a 65 70 6e 6f 70 68 66 57 64 62 62 5b 61 5f 64 62 64 68 6c 6a 69 63 65 62 64 6a 5f 61 58 5e 55 54 50 46 4c 53 4f 5f 72 72 79 70 70 68 5d 55 4a 41 36 17 09 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0f 1b 24 32 44 51 66 74 87 8f a9 a6 9b 76 73 6f 73 76 74 72 70 72 75 80 84 88 85 86 88 89 82 87 84 87 8f 88 8b 8b 83 86 84 84 83 89 86 84 8e 85 89 91 94 8d 8a 8b 8c 91 8d 92 8f 92 93 90 96 9a a3 9a 94 a0 9f a2 9e a7 ac b0 af a6 ae aa b3 9c aa a5 a0 9f 9f 9c 9e 9c 9e a0 9c a1 99 9d 9f a0 a3 a2 a0 a6 a0 9e a2 96 82 48 12 06 05 03 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 06 09 09 07 15 4b 70 8a 8e 81 75 79 85 81 81 7c 7f 80 7d 80 80 82 83 85 88 85 86 80 84 88 88 85 87 8c 89 89 80 8c 7f 8a 87 78 84 7c 80 80 7e 78 75 7c 75 75 76 6a 77 71 77 6e 6f 6e 6b 6a 70 67 66 5e 61 68 67 67 62 66 68 63 62 64 69 6d 65 5f 61 5f 61 5a 66 5f 61 60 64 6e 65 6c 6f 66 63 62 62 5e 62 5e 60 5a 59 57 56 58 57 52 4f 4f 4e 4d 5a 63 75 76 74 6c 63 5f 5a 4b 41 2f 19 08 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 0a 18 25 35 42 4b 66 6e 86 98 a0 ac 94 80 7b 65 69 6d 6d 6b 75 76 75 6f 7d 7d 7b 90 82 85 7d 82 84 87 8b 85 88 8d 84 81 84
 7f 8c 87 87 7d 86 85 83 8a 85 86 8c 8c 80 90 90 8a 91 92 9a 92 96 9a 97 99 a2 97 96 a1 a1 a1 a4 a7 a2 ad ab a4 aa a6 a0 a2 9e a0 a1 94 9c 97 9c 93 8f 99 9c 92 9b 9e 95 9c 9f a2 a1 97 9b 8f 84 51 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 09 05 1f 4b 74 82 89 8b 7b 7d 81 7f 85 81 82 80 84 75 7c 81 80 89 86 84 86 8e 85 88 83 8a 7f 8a 7e 8b 82 85 7c 86 88 80 89 81 7d 82 71 7a 7d 76 7a 6d 77 75 72 72 78 6f 6d 6a 6b 6d 69 6a 60 66 61 66 66 6f 62 5b 60 65 65 6b 62 61 64 60 62 5d 5a 5e 5f 5c 65 6b 62 65 63 66 67 64 5d 65 5a 57 5d 5d 58 5c 57 58 4c 56 4a 54 4c 48 4b 49 4f 62 6f 7b 6f 74 69 60 59 4c 43 35 1b 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0b 0f 1b 23 37 4d 54 69 71 86 9a aa a3 97 83 6f 6c 70 6e 6a 74 69 76 6f 6d 70 76 83 87 84 88 84 79 88 81 7c 88 84 82 82 85 8b 80 8b 84 82 86 87 8b 88 83 83 85 85 86 90 88 8d 86 8d 90 8f 92 8e 94 91 9b 9b 94 a1 9d 9c a0 a5 a4 ad a1 a3 9e a4 a2 a7 a8 9f a0 a3 8f 93 92 87 94 94 96 8f 92 8d 91 95 9c 92 9c 90 9d 90 93 84 55 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 0a 05 13 4a 71 7a 85 7d 7c 7b 75 80 7f 80 7e 7f 80 81 80 78 7f 7e 83 86 7e 80 7c 82 85 84 83 8e 80 8e 86 84 89 84 84 82 7a 80 7c 7c 72 76 7c 74 72 79 6c 79 7d 70 72 72 6d 6f 70 65 66 6d 66 68 6b 67 62 62 63 6a 65 6b 5f 62 62 67 68 61 65 5e 5a 5e 61 61 62 6e 64 74 69 66 6a 5f 63 60 58 62 5e 62 5c 61 5f 56 55 51 52 4f 4b 4d 49 4a 51 67 6e 74 7e 6d 67 62 5e 47 3a 38 1c 12 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 26 2b 3e 4f 52 67 71 8a 9c a4 a6 a4 8a 79 74 6f 70 78 77 6a 6e 6f 6a 78 7a 7b 80 7f 85 85 80 84 86 7b 7d 7f 88 83 87 81 81 82 85 89 81 80 84 8a 87 8a 82 81 89 85 89 89 87 8e 8c 8b 8d 8d 97 8a 96 95 93 9a 9a 92 9f a2 a0 a4 a8 a4 9d a2 a3 a1 9e 96 9c 9d a0 96 92 93 8c 8b 8d 98 93 96 95 98 92 8c 9a 8c 8b 92 96 89 5b 14 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 09 03 11 10 40 74 79 82 7d 77 7a 7d 7e 7b 83 7b 7e 79 7d 82 7e 7f 79 82 7e 86 87 88 87 7d 82 82 83 86 7d 80 83 84 85 82 79 7e 78 76 76 83 78 7c 75 74 6f 71 67 74 6e 6a 77 61 6e 6a 65 6a 67 65 64 61 5e 65 65 65 67 6d 64 61 64 69 63 5e 5f 61 58 57 62 5d 5c 62 70 6e 68 65 66 66 57 60 5e 5a 5f 59 5d 59 5b 5f 54 56 51 46 52 4c 56 47 48 49 63 6d 76 7b 75 6a 60 59 4c 3b 30 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 14 15 22 3a 4a 4d 5f 75 88 90 9a a6 95 7f 7a 6b 68 63 70 6f 68 72 6b 6e 71 6f 78 74 7b 81 7b 85 81 85 86 7f 80 86 81 84 81
 87 80 7f 7f 7f 81 84 85 7f 86 7e 8a 84 7f 82 88 83 83 89 89 8b 89 90 94 9b 94 8c 94 97 99 98 9d 9e 98 93 a6 a3 9e 9b 9c a7 8e a2 94 8c 91 89 92 89 85 8c 8a 85 8f 89 88 92 89 8d 8c 88 8a 7f 7f 5c 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 07 0c 37 6d 75 80 7e 78 78 76 79 7a 76 75 75 75 7f 7c 80 7d 7f 7e 7d 7a 85 80 84 84 86 7c 84 85 84 78 79 81 80 7e 7b 7b 80 83 7c 75 70 75 74 6c 73 6d 72 6c 66 6a 6c 66 67 6c 68 62 65 67 62 5c 63 64 60 66 5f 61 69 59 5a 60 61 64 5b 52 5b 54 5d 58 62 62 6f 6a 74 5b 64 5e 5b 5d 60 59 5f 57 5a 5b 5b 54 4e 55 58 47 4a 47 4d 48 4a 48 5a 6f 79 75 73 6b 61 59 4f 3f 35 14 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 14 18 29 39 49 55 6b 71 84 95 9f 9a 99 7e 79 68 6c 64 68 70 70 66 6d 6f 72 74 6f 6d 70 7a 7c 84 8a 84 82 80 84 81 85 85 85 7f 85 76 83 87 7b 88 84 86 80 7e 85 81 80 8a 86 7b 86 85 84 85 85 87 8d 8d 90 96 92 94 91 8d 95 9a 9e a3 a2 9e 9c 9a 95 9d 9c 95 93 8e 96 95 8f 8c 8c 83 92 8f 81 89 8b 83 85 86 87 7d 87 85 84 58 16 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 01 0f 35 62 74 79 7f 75 75 7b 78 7f 7b 7c 79 7d 7e 7c 73 70 78 78 80 80 7a 7c 7e 7d 7a 78 7e 81 83 7f 83 77 7f 77 82 7b 77 74 7a 79 72 71 66 6c 75 6d 6b 70 6b 6e 6e 61 63 63 67 69 64 5c 64 63 62 63 65 62 5f 62 62 69 5f 68 5f 5f 5d 60 64 5c 57 62 64 64 65 73 69 60 62 5e 5e 60 59 5c 5d 52 55 58 52 51 4f 56 50 54 52 4f 46 49 45 50 5b 65 6f 71 6f 6f 5f 54 4c 3e 35 1e 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 15 11 24 3a 45 52 65 6d 83 8b 9c a0 91 7e 71 68 64 69 60 68 67 65 6c 6a 6c 6f 6e 70 72 6f 7f 82 88 90 8d 85 84 85 7f 82 7f 85 82 85 7c 79 81 81 7c 7a 82 7d 7f 84 89 81 7f 84 85 85 86 87 87 8c 89 89 8d 8d 8b 88 8d 98 95 9d 97 9d 9a 9c 9a 9e 9d 9d 96 95 92 8e 8f 89 86 8c 87 89 84 83 89 89 89 83 83 84 82 7d 89 83 78 57 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 09 05 03 09 06 30 60 7b 78 82 77 72 7d 75 77 81 74 77 73 74 76 7e 78 7c 78 7e 74 74 7f 7e 75 7e 7b 80 7b 7d 7e 7e 75 7c 75 7d 7f 78 71 76 7a 74 74 6e 69 66 6d 69 6d 69 6a 63 6f 68 63 66 63 60 62 5b 62 64 63 62 60 5f 61 61 5e 66 66 56 56 5c 5c 67 5b 60 5b 62 62 6e 6c 73 6e 5f 5d 54 58 59 56 60 59 5c 5b 57 5b 4d 51 54 51 4d 4a 4c 47 3f 46 52 64 6c 71 6e 67 59 59 4d 43 36 1e 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 14 29 3e 45 58 62 7a 7a 91 9c 95 81 6a 67 68 67 6c 65 6e 63 6a 60 6a 65 68 72 6b 70 6f 74 83 87 87 8c 93 95 8e 8a 8e 84
 82 7f 7e 7a 7f 78 7e 82 80 80 7e 7d 7a 81 7f 84 89 84 7e 88 81 85 89 89 92 8b 8a 84 88 8e 8f 8d 94 91 90 98 99 9e 8d 96 96 90 8f 90 8a 8d 83 88 8c 87 85 86 7d 88 82 84 7d 7a 85 83 87 7d 80 7b 57 1b 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0c 1e 5d 71 79 79 6d 75 76 7c 77 75 7b 7a 77 79 7b 75 78 78 7b 79 7c 71 76 76 7d 81 80 80 84 76 7b 7f 73 80 78 7e 78 76 77 7a 73 70 71 71 65 67 64 65 69 63 6a 64 66 63 66 65 61 61 5a 5f 64 5f 59 63 62 5f 6a 61 5e 5e 59 55 5b 5c 54 58 57 58 55 64 6a 62 64 67 66 62 66 53 55 55 5e 4e 60 60 56 58 52 50 55 4e 4a 45 4b 4b 47 42 39 4c 56 6c 6e 6d 6a 5d 5c 47 40 37 20 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 11 1c 27 39 44 54 65 75 87 90 94 93 7b 6c 63 62 64 64 6e 64 68 68 6d 74 67 6d 6d 69 70 6b 6e 81 80 86 8b 8e 95 95 93 89 8c 8d 87 89 83 87 80 82 8b 7e 84 80 83 87 87 79 84 88 81 8d 87 80 84 86 87 90 94 86 94 8c 8d 93 96 98 9f 9a 9a 90 93 92 90 92 90 8f 90 87 87 88 8b 8d 86 85 88 83 84 80 77 82 7e 76 83 7e 7c 7c 75 5a 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 01 07 1e 5c 6e 7c 77 73 76 74 72 78 72 74 73 6f 7b 79 75 78 7d 79 80 72 79 7d 75 7f 71 78 77 79 7d 79 7d 77 75 74 75 71 71 6a 6c 69 69 75 72 6e 70 69 70 68 6a 6e 60 60 60 5d 5a 63 5e 61 60 63 60 5e 5d 62 5e 65 59 56 59 5a 55 5f 59 58 5b 54 5d 64 6b 71 67 66 6c 6b 5f 64 5a 5c 5e 5b 54 56 54 59 61 54 56 56 58 4c 50 4a 46 47 42 41 48 4d 66 6e 69 6f 6e 5f 54 45 36 21 17 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 09 1c 23 3e 49 5b 69 6d 7d 93 90 87 74 65 64 64 67 6e 6c 6b 63 72 63 6f 5f 64 6d 70 64 67 6d 6a 79 81 86 8c 8b 8d 8f 8b 8f 89 8d 89 83 87 80 85 7e 8b 84 7b 84 84 86 80 8a 87 8b 85 8e 89 8e 8a 89 83 89 8f 91 93 8d 92 98 93 93 9a 96 9b 9d 93 94 9b 8e 94 8e 8c 89 8d 8f 85 87 7e 83 88 8a 85 83 88 87 8f 84 7e 85 7a 76 5f 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 56 75 7e 7c 76 6a 75 76 73 79 6f 7a 6f 79 7a 79 70 78 79 72 72 72 7a 79 70 78 7a 7b 74 7e 76 78 74 75 73 78 6e 6f 77 6e 6c 6e 6b 63 6b 69 68 69 6a 66 62 6e 69 5f 63 64 5d 60 69 58 5f 63 62 66 63 63 5c 55 52 58 5c 56 57 5a 57 52 59 60 6a 65 62 6c 6a 74 67 6a 61 5f 5d 5c 59 59 56 5b 5c 5e 59 56 4d 55 58 50 50 47 4c 3e 4a 43 51 59 65 6c 63 65 56 50 46 35 27 11 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 10 19 2d 33 51 54 5e 77 82 90 94 8c 6e 5c 5d 5e 61 66 62 6e 60 5b 61 61 67 69 5b 67 64 63 63 67 72 77 7a 84 93 85 87 8a 8f
 88 8f 85 85 88 8c 85 8b 89 89 7e 8b 85 7c 8b 8a 88 8b 8a 8d 8e 84 8f 8b 91 85 8a 8a 89 90 98 94 96 93 94 9b 93 96 94 93 9c 8a 8d 8e 93 90 8d 90 8f 85 88 85 89 8c 8a 84 8a 7b 84 82 7a 81 80 76 5a 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 17 4d 72 74 78 6c 76 6e 70 72 6e 75 73 69 70 73 70 78 77 6a 76 77 70 72 6c 77 76 75 7b 7b 71 73 74 6a 76 6e 74 70 6b 6f 71 6b 70 65 65 64 67 60 65 5d 67 66 60 60 5f 66 69 60 62 5d 5f 51 5d 5a 58 59 54 55 63 52 53 5e 50 59 58 5a 5d 66 62 6e 63 62 6b 65 62 61 5a 59 58 5f 5a 60 55 5b 5c 5a 5f 59 4d 5a 51 56 4e 4a 44 43 3f 42 3f 43 51 5e 65 70 5d 66 4d 40 37 20 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 12 16 2a 38 44 5c 5f 74 84 8f 8d 80 68 62 52 5e 5c 60 5c 62 65 66 66 63 6a 6d 68 60 64 71 67 66 70 6a 76 7a 85 8a 8b 92 90 90 88 87 89 7f 86 81 84 8a 87 85 88 87 8c 7d 89 8c 83 8d 8b 8a 93 89 93 90 96 90 94 8e 93 95 94 91 96 93 99 92 90 96 97 92 97 9b 91 8c 8d 89 8f 92 8b 8e 8f 8f 8a 89 87 8d 90 8d 88 80 84 7a 7f 63 2a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 17 48 6a 76 7a 76 6f 77 71 76 70 6b 78 6e 78 77 71 78 73 76 76 6e 72 75 73 77 72 6e 74 6e 77 6b 73 76 77 6c 78 69 6e 6a 65 5f 6b 64 67 67 68 65 68 67 5d 62 5c 57 57 5e 5c 62 61 5e 5a 5d 5e 59 5d 56 50 58 54 53 57 57 56 5f 5f 5f 5b 66 5b 59 65 5e 64 69 60 69 5e 55 55 58 5f 5c 5a 53 59 65 62 62 50 53 57 50 4e 4d 48 3f 3b 37 3b 4b 4c 5c 6a 63 65 5a 50 3f 32 24 14 07 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0d 1a 26 3a 4c 5c 63 76 84 88 98 82 67 5c 5a 54 5e 5b 61 5c 64 67 68 68 67 67 71 6f 62 68 5d 63 6a 6c 70 76 7e 78 80 83 8b 8d 94 91 88 88 85 8d 8b 86 91 8c 8a 87 8a 85 83 86 8f 8b 94 8c 91 98 94 9f 8f 94 94 9d 94 98 98 92 9c 90 9d 99 97 90 98 91 9a 91 97 97 8f 95 98 8d 9a 99 8f 8f 91 91 93 8d 8e 94 91 89 8c 87 83 6c 2f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 4a 71 83 89 85 81 70 79 7f 75 70 76 71 78 7e 81 73 7a 7d 7b 75 78 80 77 78 7f 77 74 7a 75 71 75 72 6a 7a 75 6c 6e 70 6e 64 69 68 64 63 62 60 65 64 66 64 69 61 5c 69 5f 63 60 5b 56 50 58 58 58 5b 54 52 58 51 55 5b 5d 63 66 68 67 6a 68 70 73 69 6d 65 77 6b 5f 5f 5f 52 61 64 5f 64 5d 6b 67 5e 5c 53 55 52 4b 53 48 46 4c 3e 40 46 4e 57 6b 66 61 53 48 42 30 22 13 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 17 23 3e 46 54 6c 76 7b 87 87 80 64 56 5a 4f 52 5b 58 51 60 5f 68 69 6e 72 70 6b 69 62 60 62 5f 61 65 6d 78 6d 6f 72 7f
 8c 8f 88 85 8c 83 89 8a 86 87 7e 8a 8b 85 86 88 7f 8e 86 92 89 91 91 91 93 8c 94 9a 8f 90 94 97 8f 90 89 87 93 93 85 94 8d 94 93 90 94 93 90 84 98 90 94 9b 93 92 93 96 94 92 84 84 85 87 85 86 79 30 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 04 06 12 3c 78 8b 8a 7f 89 78 84 79 87 80 7b 7d 82 7d 76 80 79 7c 7e 78 73 78 6c 78 7b 7b 7c 78 71 6f 77 6b 74 71 72 70 6b 68 67 66 5e 66 63 6b 67 61 60 64 5c 65 61 5c 5c 61 5e 5b 59 55 53 54 4e 57 54 56 51 54 58 55 50 4f 5d 6b 69 6b 63 65 60 67 72 71 77 7f 78 63 5a 5f 4d 56 5b 63 61 66 64 6d 6d 6b 59 57 50 50 4c 4a 47 46 3e 44 39 3e 47 48 67 63 64 5b 4a 40 34 1c 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0a 21 34 45 56 60 71 7e 8d 8b 79 67 52 5a 55 55 55 4d 5a 54 5a 61 62 6f 72 71 6f 76 63 63 64 61 5b 67 61 6a 6d 71 7c 76 75 81 79 84 86 86 86 88 8b 8b 84 81 83 82 88 89 8a 86 8c 8d 8d 85 8d 8b 92 8c 92 91 92 8f 8d 89 8d 8f 8b 96 90 8a 88 90 8d 91 8e 81 89 8b 87 93 8e 88 8a 94 91 92 8b 90 8b 93 91 89 87 8a 8d 81 72 37 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 3e 79 97 9a 91 84 88 80 89 86 7b 7d 79 77 7e 83 7e 7b 7c 7d 83 7b 7d 7e 7c 7c 80 7b 7e 74 75 72 6a 6a 77 6b 69 6b 69 6a 64 63 6d 65 62 60 65 62 60 5d 66 5a 59 5a 61 5b 5c 55 57 5a 57 5a 56 54 51 50 57 4f 52 5a 66 60 69 6c 70 64 63 69 68 6c 79 7e 80 79 62 5e 54 53 5b 50 5a 5a 67 6e 6f 6b 5d 5d 50 4d 45 4b 4b 4d 47 40 43 3a 36 44 52 59 60 62 55 4f 40 36 1d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1e 37 4d 5c 68 78 7d 88 8a 71 64 53 57 4e 5a 52 5b 4d 55 52 54 5f 5d 62 6b 6a 65 62 64 66 66 6f 69 66 6a 63 6e 77 6d 74 7b 7d 7b 79 79 7a 82 7c 89 81 84 8d 84 8b 83 85 8b 91 8e 8b 8c 88 8f 8b 8b 93 8d 92 90 81 8a 8b 84 87 8a 83 86 89 86 87 7d 7f 7f 85 7c 83 85 87 89 88 80 89 8f 91 84 8e 8f 88 8c 89 8b 85 83 69 3b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 08 2a 79 90 97 95 8c 8d 8d 8d 83 84 7b 76 80 82 84 85 8a 7c 7c 82 87 85 84 89 85 7e 81 74 73 6d 75 71 6f 66 6d 69 64 6f 61 62 62 61 5c 5f 63 63 59 5e 5b 61 5a 5a 60 59 64 5f 5f 58 55 4e 54 56 58 5e 53 52 52 54 5d 6d 73 79 7e 76 76 67 6a 6d 70 7c 85 7b 71 5b 59 50 59 55 5d 5b 5f 6a 6a 76 6c 60 50 5a 56 43 4e 4d 48 4f 41 3e 3d 3d 47 52 59 68 5e 57 4f 3c 31 20 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 22 2f 45 54 62 79 7e 88 89 76 5f 56 57 4d 57 52 58 56 4b 4e 58 53 5f 5f 65 68 66 67 69 6b 68 69 5f 62 63 63 69 68 6e
 6a 72 70 6f 77 77 7a 7b 84 77 7f 7b 85 88 7f 7f 8b 83 83 80 87 87 82 89 8b 84 7f 7d 87 80 7d 84 85 84 7b 7f 6f 7c 7e 79 81 72 79 79 7f 72 73 78 7c 7e 78 82 7a 7b 80 75 82 7f 78 76 76 86 7c 77 6d 43 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 6e 8c 92 94 8c 89 8c 84 89 85 82 77 86 89 78 8b 82 8b 84 83 84 7e 84 7f 78 7a 6f 6e 6b 6c 6e 64 69 66 6e 69 68 63 5c 60 62 60 62 60 5f 5f 5e 5f 5f 59 59 56 54 5b 5e 56 5a 52 52 57 53 57 54 55 51 53 5f 5b 66 70 7a 70 73 6f 65 61 63 69 65 6b 72 67 61 55 58 52 53 55 57 59 62 67 75 6c 66 58 55 55 52 46 49 52 4b 46 41 44 35 39 46 44 59 65 5e 59 48 39 2d 16 0c 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 16 29 46 4e 5e 6f 7d 7f 88 72 64 4d 4d 54 57 55 5f 56 51 56 55 58 55 56 5f 61 68 67 72 6b 63 68 5f 65 69 69 6e 6c 5d 64 6a 67 61 6a 6b 6d 69 6f 74 7a 71 77 77 73 7e 7b 7b 79 79 7d 79 85 74 7e 79 7a 77 79 76 75 7e 79 75 7a 6e 77 75 76 6e 76 6c 73 71 67 69 6c 73 6f 71 68 63 6c 68 70 6f 6e 71 6b 6d 63 71 71 70 63 35 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 2a 66 83 89 8e 7a 7f 83 84 7f 7f 7c 7b 86 7e 82 7c 85 7d 81 80 85 85 7f 84 86 7c 7b 71 74 6a 6a 64 60 67 64 5d 64 67 68 62 61 5f 5c 56 62 58 64 5a 57 5d 5e 57 53 59 5a 52 4c 4c 4d 54 56 52 56 52 57 53 5b 5b 63 5e 5f 66 65 62 65 5e 63 67 6a 6b 60 60 57 5a 59 5a 54 56 5b 5d 68 6f 67 69 58 50 4b 4e 4f 50 4a 51 40 40 3e 3f 43 3e 48 41 54 63 5b 5b 40 33 27 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 2a 3b 53 5a 66 7e 88 88 75 63 5b 4e 49 50 55 55 52 50 4c 51 57 55 56 5e 5c 61 5f 5f 6f 6c 69 69 63 63 69 6b 66 65 6a 68 66 66 66 6b 65 70 68 6d 6a 6e 73 72 6d 6d 77 70 77 71 70 77 71 78 72 70 71 66 65 73 69 6f 6e 64 64 70 6c 6e 70 61 69 6f 6f 6e 68 6e 61 67 67 60 68 70 63 64 6c 63 66 5f 6a 67 5f 62 5e 5b 53 3a 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 23 51 77 7c 7e 70 6f 74 7a 74 7c 7b 7c 7a 7b 81 77 84 80 80 81 7b 81 83 7e 7e 71 6a 73 6a 66 6c 62 64 60 6e 5d 6c 6a 64 67 62 60 60 56 5c 5b 61 59 5e 5b 55 53 5b 5c 56 50 54 52 58 58 55 53 53 56 55 57 5d 55 60 5a 5b 5c 62 5e 63 63 5f 61 5c 65 5f 54 5f 56 57 56 55 5c 57 61 69 60 6c 57 5a 55 4f 52 4f 41 4c 4f 4b 45 42 3f 37 3d 49 4d 4f 63 63 57 49 38 1e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 08 21 33 47 61 6c 70 7b 86 7a 6d 59 50 56 4e 56 5f 51 53 57 51 51 55 5a 58 57 52 60 60 6b 74 72 6c 70 6a 67 64 65 66
 65 68 68 64 64 64 67 67 61 65 65 6d 6f 6b 68 61 70 68 64 6c 66 68 62 66 66 67 63 6c 62 63 63 63 67 62 5e 63 63 5f 5f 60 6b 61 66 6e 69 5c 66 65 63 65 64 6a 5f 65 6d 64 5c 64 64 65 5f 61 5b 5a 52 42 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 19 50 6b 71 6d 70 73 6c 6e 6f 6e 6a 66 6c 72 75 75 77 72 75 76 73 7e 79 79 78 75 73 6d 69 6a 6a 5a 61 6d 60 64 5f 5c 66 59 5c 62 59 64 65 63 62 62 5e 60 5f 57 4e 5e 58 51 55 4e 5a 58 58 50 5f 5d 59 62 5b 58 55 50 51 57 5f 5c 64 63 69 62 63 62 60 5b 55 62 54 4f 51 59 5f 60 64 5b 5d 58 55 5a 57 4f 51 4b 52 46 42 49 44 48 42 41 3d 42 4c 60 59 57 3d 24 19 08 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0d 14 2a 39 52 67 72 81 8e 80 67 52 52 49 51 4d 54 4a 57 4e 56 5d 58 55 56 52 4e 57 56 66 69 69 5f 61 6b 6c 66 65 6e 66 67 61 5c 61 64 5d 5b 60 61 64 5a 67 61 6f 64 60 5f 6a 5e 64 62 61 67 67 65 5a 64 57 5d 5f 5e 59 5d 5d 61 61 62 64 5b 63 60 65 62 5d 63 66 5e 5b 64 66 5a 61 64 68 64 5c 5c 5c 61 58 5e 58 56 50 30 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 3f 61 66 68 6a 61 68 61 6f 5f 5f 62 66 6e 6c 6d 6d 69 6b 73 69 74 72 67 72 70 6b 6b 66 65 67 68 5f 63 5d 60 5e 64 64 61 62 63 56 5b 5e 5b 5d 58 5c 58 57 5b 5a 54 56 50 4f 54 55 59 52 53 5d 5d 60 5e 56 56 55 4f 54 58 5f 5b 5f 62 66 64 61 56 5d 5d 5b 58 50 4b 51 59 54 5a 5d 55 5b 59 4f 4e 4f 46 4f 41 46 47 47 4b 41 49 3a 37 3c 43 53 5c 55 3e 34 23 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 10 1f 3c 55 64 67 89 8b 85 6e 55 4d 4c 54 51 4f 52 51 52 4f 53 53 50 52 55 56 50 53 58 60 65 64 6d 70 61 6b 67 69 73 67 64 63 62 66 65 60 67 67 5e 66 56 6a 63 5e 63 5d 5a 64 5b 56 64 5a 5d 5d 63 5e 5b 5e 5a 5b 59 5b 5e 5b 56 56 5b 62 64 61 5d 5e 5d 5f 62 56 60 58 5e 5e 5f 58 5b 56 53 5f 60 58 59 5f 5c 53 4c 3a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 35 60 64 5f 6a 69 66 6a 63 68 63 60 67 62 64 6b 67 67 65 6b 65 6a 63 6d 64 61 66 6a 63 64 64 61 68 63 68 6a 5f 61 5b 5c 59 56 56 5f 5c 5b 5f 62 5f 63 56 5f 62 5a 54 52 50 4d 5a 59 52 62 60 5e 58 5a 5e 54 55 58 5b 60 63 70 64 62 63 5c 57 5b 6d 59 5a 55 5d 57 54 5d 5d 62 58 53 50 54 4c 5a 4b 44 51 49 4d 4e 4e 4d 47 43 47 3b 40 49 48 50 4d 3a 2f 1c 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 08 1e 39 4a 61 6d 7b 8e 85 77 59 53 4b 4d 55 54 53 51 46 4e 50 61 50 5b 58 55 51 4e 5b 58 59 5d 63 64 68 64 5e 6a
 6c 5f 64 60 63 65 5a 5d 66 61 67 69 60 5e 61 59 5d 5e 58 64 5c 59 61 51 5e 59 55 5a 54 5f 62 5d 5e 5a 60 5d 59 5e 5a 5e 5c 59 57 5b 5c 54 5e 5b 5c 5d 5c 58 5c 5f 55 5b 55 60 5e 5f 53 5c 55 50 53 41 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 34 58 59 6a 63 64 63 61 6e 5c 62 51 59 5f 5d 5e 60 65 64 60 63 63 5f 61 64 67 5f 62 60 62 66 61 5e 58 5b 60 5e 63 5f 59 5d 64 5f 61 56 5b 58 5f 58 5b 59 4f 5c 53 5c 50 53 59 55 62 5b 64 66 60 5d 5a 5c 61 64 66 65 69 6f 66 6a 64 62 56 58 63 65 68 63 5b 5e 55 59 59 58 5d 63 56 51 55 51 4e 4b 41 51 4c 4d 43 4c 4a 44 41 41 3e 3e 3f 44 4b 3d 33 22 14 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 10 17 25 3f 56 6b 79 83 82 73 5a 50 51 4f 52 56 56 55 54 4f 50 4f 4a 56 51 4f 4f 4a 49 59 4d 51 56 56 5a 5c 63 64 62 67 64 61 5a 5e 5c 62 5d 5f 57 66 62 5b 5b 5f 58 5f 58 5e 53 58 5e 64 5f 5c 5c 56 51 4d 5a 57 57 5d 54 52 59 52 4f 54 55 54 56 57 53 5f 60 59 59 55 58 5a 58 54 59 53 54 57 5a 5f 57 5c 51 53 4c 3f 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 2e 61 66 63 6a 60 5c 5f 5d 62 64 60 5c 66 59 62 61 5f 5c 59 5f 5a 5a 63 5d 60 5b 59 61 5c 62 61 5a 58 62 56 61 5c 56 5e 5a 5d 5b 57 5c 5c 5b 59 4f 4e 5c 51 52 4d 56 53 4f 60 61 5a 65 60 5f 5d 5c 5a 5a 64 69 6e 69 69 5f 5d 66 5e 62 60 5e 5e 62 5e 67 5d 5f 60 5e 67 62 64 64 57 59 57 4b 4a 47 4b 53 4d 45 42 4a 46 46 3f 40 44 3e 3a 37 3d 2f 22 18 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 05 0b 1a 20 3c 4b 5c 7e 80 81 75 5b 51 51 55 55 50 48 50 4e 4e 52 4f 52 4e 5a 4e 52 55 52 4d 4c 58 56 56 5d 50 5e 5f 61 5f 62 5f 5d 5f 5c 5d 63 5f 66 5c 5c 5e 64 5c 57 5e 5e 5f 5b 5d 5e 5b 5a 55 57 52 59 57 5c 5b 5c 5d 51 54 51 56 5a 56 5d 50 56 53 51 58 5a 59 52 54 57 58 4f 5f 55 50 5a 52 55 50 5c 52 59 51 46 3a 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 2e 5a 63 66 58 66 5f 61 5b 5d 60 54 61 63 60 55 58 5c 60 5d 5c 5e 54 5c 61 5b 5c 52 62 5d 5c 5d 5d 56 5c 5d 5e 5b 55 59 5c 62 5f 4d 62 5d 58 5a 54 4d 5e 53 50 54 54 4d 51 5f 5c 5e 64 5d 60 60 5d 59 59 62 60 65 64 60 65 5f 57 68 6b 63 62 63 6d 6d 66 62 5d 5d 61 6a 5f 68 56 5c 54 59 50 4f 4c 52 51 4b 43 49 48 49 46 40 42 32 41 40 3a 3d 21 1d 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 13 14 22 3f 60 6d 8c 85 72 63 57 4e 49 52 4f 51 4e 4a 4e 4a 46 59 54 55 52 47 4a 51 4e 59 52 56 55 4d 58 5a 5c
 5e 5a 58 5c 61 5b 57 5e 5d 5f 57 56 5d 60 5c 68 5e 5d 57 5d 5f 5a 55 56 5c 5a 51 54 56 5a 5a 53 56 54 4e 5d 4d 59 4d 55 56 54 55 54 54 55 57 54 5d 59 56 54 57 54 4c 4f 54 4f 59 59 47 56 51 4f 54 42 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 29 56 58 5c 63 5f 61 5e 64 60 63 57 5e 5e 5d 5f 5f 59 61 65 5b 5d 5d 5b 5d 57 5a 5c 63 51 67 54 61 5a 61 5c 5f 5f 60 5c 52 5a 5e 58 58 56 54 55 56 51 53 54 54 5d 50 5a 59 57 65 62 65 56 57 64 57 58 52 5f 61 60 5a 62 5e 67 64 61 69 69 5c 68 70 61 69 65 5c 63 59 66 67 6a 5e 5e 59 5e 5b 51 4f 55 48 4a 4c 49 4d 48 48 45 42 41 3f 3b 33 34 23 11 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 19 1f 32 50 6b 7d 7c 70 5e 52 4a 4b 52 4e 4a 46 4f 52 4c 44 47 4f 52 52 4e 4d 51 55 4e 50 55 47 4c 4b 4a 53 51 59 52 54 4e 4c 4c 56 5a 4b 57 4f 4d 5b 52 57 58 51 5a 55 49 5a 54 54 4b 50 54 4e 4c 4c 51 4c 57 54 56 57 4f 58 54 4e 57 51 52 5a 5c 55 56 55 58 51 5d 52 50 54 57 53 55 4f 52 4e 54 4d 53 54 51 3a 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 23 4f 5a 61 5a 59 5e 60 5b 5f 65 59 60 5f 62 5a 62 63 66 5e 5c 5e 5a 5f 62 60 65 56 5f 58 60 5f 5c 5b 56 58 58 5b 59 50 5a 54 54 5a 56 54 56 61 52 55 57 4f 53 53 4f 4f 55 64 69 62 5f 59 55 59 56 52 58 55 5a 5a 58 5e 5d 65 62 5f 66 6d 6f 6e 62 6c 64 58 62 63 60 6a 65 68 61 60 62 62 54 62 53 54 52 4a 4e 44 4c 47 46 53 3d 46 38 31 34 2e 1e 19 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 0a 09 1b 2f 48 65 74 86 75 5c 4e 4e 4b 52 53 4b 4d 47 51 4b 47 4a 57 4f 51 51 50 55 50 4d 4e 51 50 4c 4f 4e 53 4c 54 50 46 4a 4d 54 4d 46 51 40 4a 4d 4c 58 53 52 50 51 4a 44 4a 4f 4b 48 4c 4c 4d 47 4a 50 56 5b 58 53 52 51 50 5a 54 51 54 53 55 56 55 49 56 58 4b 55 54 53 4b 4c 4e 53 54 54 56 51 59 47 4f 42 41 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 23 49 59 53 60 5d 5a 5e 5c 5d 56 58 63 65 5d 5a 56 63 61 5c 63 59 5d 5c 61 64 62 5e 5c 5c 69 58 5d 56 5f 58 57 55 64 5c 59 5f 4e 58 58 58 5d 5b 59 54 58 59 54 58 5a 53 5c 59 62 60 61 5e 57 57 51 56 5a 52 56 54 54 5d 53 60 57 65 6a 7c 74 74 72 75 65 6d 6a 64 64 5b 64 5b 61 64 64 67 61 60 57 5e 52 4b 44 45 47 51 4c 4d 45 3d 40 33 3a 20 16 16 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 01 11 08 0a 17 23 33 56 70 85 72 62 54 4b 4c 51 4f 44 4c 53 4e 4b 51 4a 47 4e 4e 50 4c 53 4b 4e 51 4f 4b 50 4d 51 4f
 52 4a 4c 47 51 49 41 4d 45 4a 4f 4c 49 50 4a 42 4f 4c 4c 4b 4e 49 4d 41 4d 4c 52 45 46 4c 45 52 4a 4d 4d 50 4d 57 56 50 51 4e 52 53 54 53 55 53 52 52 55 4c 57 4c 51 52 4e 51 53 4c 48 4f 50 4d 42 3f 15 06 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 1c 4e 5c 52 60 58 50 5e 68 59 57 5a 5e 5c 56 5d 5d 64 65 65 65 67 67 69 64 61 66 62 5f 60 61 61 61 5e 57 5f 5e 5a 5e 5e 53 52 5b 58 5b 5a 54 57 56 56 58 5d 60 63 5b 58 5d 61 61 60 63 56 57 60 5f 5a 4c 4c 51 52 53 57 56 60 64 6f 85 79 7a 7b 81 7d 7c 69 70 66 5c 67 5a 62 5a 67 5f 66 62 5f 5f 5a 5a 4f 48 47 4c 4f 46 47 3f 3d 38 34 34 20 14 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0b 0b 16 1d 2b 47 62 7c 74 58 5c 4f 46 50 4e 4b 49 47 51 47 48 4b 52 4e 4c 4a 4b 52 4f 4b 4e 4a 4d 44 47 45 52 49 49 4b 45 48 4b 44 50 48 4b 4e 4b 47 3c 4e 46 46 45 45 4c 4b 41 47 46 44 4a 42 44 3d 48 54 4e 4f 4d 43 45 5a 54 58 51 54 59 5b 57 50 4a 50 50 54 52 4e 53 4f 49 50 50 4c 4c 4e 45 48 4a 4c 4c 49 34 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1c 47 54 56 5d 56 5b 59 5f 59 59 58 5e 5f 56 61 5a 5c 67 62 65 69 63 61 6d 67 66 57 6b 58 63 59 5c 59 56 51 5a 5e 56 59 5a 58 56 50 5e 52 54 64 57 57 62 5c 5f 5e 61 63 56 5c 55 5b 5f 5f 57 55 5a 55 53 4a 4b 4b 52 54 5c 61 68 76 72 84 81 84 8c 87 80 7d 76 76 68 61 61 61 65 65 64 6a 5b 59 5d 58 58 4d 47 45 41 49 4e 4c 45 46 39 3d 25 1f 0c 10 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 07 0f 10 1b 2c 4f 64 76 5f 50 55 42 4f 4b 4c 46 47 4b 46 4e 52 43 4b 49 49 50 47 4d 4b 46 4c 4e 49 4e 4f 50 49 4f 49 41 49 41 43 48 43 4e 44 45 49 43 49 48 48 4e 4b 49 3d 4b 3f 42 4a 46 44 44 3f 4a 44 4b 49 3e 4e 4c 4a 4a 54 4d 4d 50 51 50 57 45 4b 4a 4c 47 4a 4b 47 49 47 51 4a 41 4a 49 47 4c 43 46 45 3b 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 17 4b 53 55 59 4f 51 57 59 51 54 5c 5e 59 5a 54 62 5a 61 5f 64 66 65 6b 6e 71 67 64 62 5d 5d 5c 5a 55 59 51 5f 56 58 57 53 55 57 5a 52 57 61 62 62 5a 5d 5b 61 5e 55 63 52 5c 60 53 5a 54 58 52 52 4d 4a 4b 50 49 4c 51 5c 61 71 75 7b 83 8a 90 90 90 90 7e 7f 71 6d 6a 63 69 64 67 63 61 59 5d 56 54 4f 4d 4e 47 43 48 45 41 3e 37 38 2a 21 1c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 06 10 09 11 16 1a 2e 44 5e 6f 62 55 51 4c 4d 46 4b 4b 48 4c 52 4d 43 4c 4c 45 4b 4f 4f 55 4b 4e 4f 50 45 4b 4a 4a
 45 4b 4a 50 4d 4b 47 47 48 47 45 47 4a 43 42 46 4d 4f 46 4b 44 46 4f 42 50 45 49 46 3e 44 44 4c 4b 41 45 49 47 4e 49 4d 56 53 50 57 51 48 46 4a 4d 49 4d 47 48 46 53 4a 49 48 4e 4a 48 46 45 3d 4b 44 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 12 43 4e 59 55 57 53 57 50 56 57 5a 5b 5a 4e 5f 58 65 65 60 69 6d 68 71 75 6c 72 67 5f 62 5c 5b 58 59 59 54 54 55 56 56 5b 5b 5e 5a 52 63 5a 61 65 61 60 5f 65 62 65 5c 5f 5b 52 57 5b 50 59 50 4e 50 4e 50 4b 4c 53 52 57 5e 6b 78 89 85 96 99 93 9d 94 8a 8b 84 80 74 6b 72 6d 68 6f 5e 5f 60 56 56 50 47 4c 4d 4c 54 42 45 45 36 36 27 20 0f 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0d 0f 09 15 1a 2e 3d 58 60 5a 56 52 4c 4d 4c 47 44 44 4f 48 41 47 46 4b 4d 4a 47 47 4a 49 4e 4b 51 48 4e 4b 4a 4a 4c 3f 4a 46 49 42 45 44 40 3e 3f 40 4b 43 49 45 43 46 45 46 45 47 45 46 47 50 47 3c 39 45 47 3f 44 47 44 46 45 4e 49 52 53 51 54 4c 4f 4f 4a 4c 45 45 46 46 4c 47 48 44 4c 4c 47 41 4e 45 47 44 41 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 3c 55 57 54 53 49 55 50 57 5e 57 5d 5e 5c 5d 5b 59 5b 5e 6b 61 64 71 73 72 6a 62 67 5b 5f 5b 53 55 52 50 55 55 4f 53 54 55 5b 5b 5e 56 58 5f 5d 5a 5d 60 5e 61 62 57 5e 4e 52 50 57 4e 59 4a 4f 4e 49 49 4b 50 53 53 54 5c 6a 76 81 90 9c 9c a0 a1 a1 92 87 81 78 7b 72 6d 6c 67 63 64 5a 5a 54 51 49 4c 50 4b 45 4c 50 48 37 36 28 26 1f 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 05 03 0f 0c 15 22 2b 52 5b 5c 51 49 4b 4f 4e 49 4d 43 45 50 43 42 4c 48 49 44 47 41 41 4f 4e 44 53 49 4b 48 4c 4b 46 3f 44 47 47 39 46 3f 55 3e 3f 48 50 42 43 3e 44 40 47 49 3f 44 42 47 48 4e 35 43 41 47 49 3d 3d 3e 4e 40 41 43 48 52 4e 4b 52 50 53 46 4e 4f 44 45 4a 3d 4a 43 47 4b 47 47 48 47 41 49 47 46 44 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 39 52 4a 56 50 51 4f 52 55 54 48 5c 54 51 59 5d 59 5d 54 5c 63 64 69 67 6f 71 69 5b 54 5b 52 59 5d 58 5a 56 5a 52 5f 50 56 5d 57 59 55 55 54 56 5d 5e 4e 50 56 4f 59 4c 5a 55 53 56 57 54 4a 46 42 49 45 4b 4e 4a 51 53 5a 65 66 70 82 8b a0 a4 a1 a1 89 85 7b 76 75 6a 6f 70 63 69 5b 5b 59 54 4b 4f 55 4d 4f 49 4b 41 3c 31 2c 2c 1e 10 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 10 12 12 12 1b 25 35 3e 54 55 58 4d 4f 4e 4d 4d 49 45 50 50 49 44 4b 44 4c 4c 47 4c 4a 49 4a 4a 50 41 41 41 4c
 47 4c 49 48 47 48 44 50 44 41 4b 48 3f 43 45 4a 45 49 3f 50 46 4e 44 3d 47 45 42 48 44 44 48 49 47 43 3a 42 39 43 49 44 47 42 4b 4d 47 4f 4b 4d 4a 4a 4c 50 44 50 47 44 45 3f 4b 45 48 40 49 45 48 42 2e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 38 4c 52 54 4d 4f 59 5f 4d 4f 4e 58 58 51 55 56 57 5e 58 5b 5c 62 65 61 5e 6a 63 66 57 5b 57 55 55 5b 57 55 56 54 53 54 53 55 52 51 52 58 51 52 58 5a 53 56 5a 52 53 49 57 51 4a 4c 4b 52 53 4e 50 4c 49 4b 4e 4a 4b 58 5a 62 62 6c 78 87 8d 98 9a 95 8c 82 73 72 71 64 61 66 62 64 56 57 59 4f 4d 51 54 4a 4d 4f 46 45 41 2f 2c 28 18 13 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 09 0b 09 13 15 15 23 2f 32 50 56 51 47 4c 56 4f 49 4a 47 46 45 4d 4e 45 4d 4d 43 45 41 4b 49 50 46 48 45 44 4a 45 47 4f 49 46 46 3e 3f 4d 43 49 43 48 43 44 49 42 4a 44 40 43 41 49 47 45 48 40 3f 49 48 46 49 43 48 46 43 46 46 3a 3f 42 4a 46 47 4b 3f 49 45 45 4f 49 4a 4b 3c 49 4a 4b 3a 44 4a 44 48 44 45 4a 41 48 2c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 30 4f 50 51 51 4a 52 4d 4a 51 4f 58 54 4f 4f 5a 50 5b 59 5d 5b 5d 66 60 60 66 65 5e 55 5a 58 5d 5a 56 54 56 57 51 50 52 55 56 53 50 4f 50 51 52 51 54 50 4f 5a 56 56 52 56 4d 4c 4f 4c 4b 53 4a 4a 47 4b 4d 45 4f 53 50 55 54 61 64 70 77 7f 91 90 94 80 77 77 72 64 67 64 65 55 63 65 5b 58 54 50 4b 46 4c 55 53 4b 45 3d 33 27 1e 1c 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0f 10 12 25 29 3b 46 50 53 4b 52 4a 44 4a 46 45 4c 42 49 3b 3e 47 42 52 4a 48 42 43 41 42 48 40 45 41 49 3e 4e 41 4a 40 3c 40 42 40 41 47 40 42 40 38 4b 42 45 48 49 3f 45 42 45 45 44 3b 4b 3d 3f 41 44 3f 3f 49 44 4a 3a 3e 44 41 42 3d 3b 3c 40 44 42 4c 43 49 44 41 49 41 42 43 43 4a 48 44 41 46 4c 49 45 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 27 4c 54 56 53 48 4a 53 43 58 47 50 4e 4c 52 50 54 58 59 52 59 54 57 5a 56 65 5f 5d 5a 55 5d 52 57 56 55 56 56 4f 51 4f 51 5c 54 50 56 5a 4a 4f 55 56 52 52 56 50 51 50 59 50 4a 4b 48 4e 49 4b 52 4e 48 4a 58 4d 53 54 55 56 50 5b 61 65 71 72 73 85 76 78 7b 70 69 60 5b 61 5a 5f 5e 54 61 48 4a 50 4c 4e 4f 49 4b 44 3d 34 25 21 11 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 12 12 13 20 31 37 47 4e 54 48 4d 4f 44 4c 46 44 4d 45 4f 3d 47 45 44 4c 4b 42 40 4e 44 3f 44 40 50 48 4f
 3d 44 44 46 4a 48 3d 46 4b 44 4b 44 43 46 49 45 46 40 40 45 47 45 41 4c 4b 44 44 41 45 46 47 3c 44 45 3e 45 3a 3e 42 44 45 3b 3c 37 3f 3d 3c 41 49 47 47 45 41 4d 4b 43 44 4b 46 44 44 4f 51 4d 3f 3d 2c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 27 4e 4d 57 4a 51 52 53 4c 4b 4b 52 55 54 52 52 5b 56 5b 56 52 5e 53 56 58 5a 57 5a 58 5e 55 56 53 52 5c 59 52 58 54 4f 54 58 52 4a 52 54 5d 58 55 53 52 52 5b 5f 55 52 49 4f 4e 4b 48 4e 4b 48 4e 44 45 4f 51 47 4c 57 4a 58 5a 60 5b 61 64 6d 6a 78 76 75 7a 6e 6b 63 5e 5c 54 54 5e 58 5c 54 53 50 46 47 4f 4e 45 4b 3a 2c 23 13 0e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 02 0f 1e 1f 22 27 45 4c 54 53 48 4c 48 47 48 47 45 39 3e 45 49 45 46 3c 45 42 49 40 4f 45 4a 4a 4a 49 3f 47 49 42 45 4a 44 3e 45 41 3f 40 46 45 3d 43 46 44 41 4c 3e 3f 45 48 46 46 44 44 43 41 3f 46 44 4b 44 3d 3b 3f 41 48 42 42 3c 41 40 3d 3e 3d 3e 44 3b 42 4a 42 42 44 44 42 45 47 4f 44 47 46 3f 43 35 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 1b 43 49 56 50 47 49 4f 4b 4c 4f 50 59 4b 50 52 4c 5e 57 51 50 59 56 56 55 55 59 59 52 55 55 5a 55 54 5e 5e 5a 60 56 59 55 5c 53 55 4d 58 57 4f 51 56 52 4a 50 52 4d 4c 58 55 51 4a 4a 4d 45 46 50 48 40 42 50 4e 51 4a 52 58 4a 58 54 56 5a 63 65 6f 66 6f 64 64 6e 59 54 51 52 55 52 53 59 4f 51 4d 4c 4c 4a 47 4d 36 3a 23 21 15 0a 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 0a 0e 10 16 1e 20 32 3f 3f 4c 4d 4f 48 42 44 4a 4a 41 4b 47 49 3f 4c 48 40 42 49 4c 43 43 4b 4e 42 44 42 3d 44 42 44 45 40 42 4b 40 4a 46 43 42 44 45 40 46 47 46 44 43 39 4a 4a 45 4f 4c 40 40 44 45 47 4d 4a 38 3f 43 43 37 3d 3d 39 40 41 3e 3f 3d 32 40 42 3e 3e 3f 42 41 3f 46 3b 44 3b 41 40 40 3b 3c 36 38 2a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 18 45 4c 4f 55 4c 52 4e 4c 44 4d 4f 4e 51 51 4f 58 4c 56 57 53 50 53 50 54 4f 59 52 57 5e 5b 60 5a 62 61 53 63 5c 51 53 53 51 4c 52 51 51 51 50 50 4f 50 53 50 45 52 52 51 47 4e 54 45 54 50 4e 4b 53 4d 4a 4e 48 50 4d 50 52 4b 53 55 55 52 53 56 59 64 5f 67 61 60 5c 56 57 51 4f 54 54 5c 54 4c 50 4f 49 43 45 3e 3a 2d 21 10 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 09 13 12 12 1f 2b 35 43 55 4d 4d 4e 41 41 46 42 48 45 46 4a 42 41 39 41 41 41 49 4b 45 48 49 4e 43 4b 4b
 40 48 4d 3a 44 3f 45 47 46 3e 49 48 4a 44 3f 43 41 43 44 45 3d 42 47 40 46 42 42 42 44 41 4f 37 22 2f 49 47 3f 3a 36 3c 3e 41 3e 38 35 36 36 3b 43 3c 42 3c 36 38 3d 3b 45 3c 3a 3b 40 44 35 35 3d 33 2a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 24 49 4a 53 4e 4c 54 4d 52 52 4f 4c 55 4d 4e 51 4d 54 4c 53 58 54 47 57 5b 50 51 59 59 5b 54 5b 63 5b 5a 5a 52 50 55 4d 57 4e 4a 45 48 53 57 4c 49 55 4b 4d 51 4e 4f 50 4f 4c 4a 49 4a 53 47 4b 4d 4e 51 4a 4c 4a 47 49 56 50 53 51 54 5a 50 49 56 54 57 5a 5c 5b 5f 5a 5a 59 56 51 57 57 55 4e 4e 4a 49 50 44 41 3e 2f 2e 15 0d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 10 0f 13 1b 1a 25 3b 40 4f 53 4e 4d 4c 43 48 40 41 47 45 45 49 40 45 43 47 46 45 48 47 42 44 48 44 48 43 42 44 44 46 44 46 44 47 44 46 4b 43 4d 45 3b 43 45 3b 45 41 46 48 43 3c 4a 40 40 4a 3f 47 42 40 45 47 4a 3f 3a 3e 3f 3d 43 3a 39 3e 38 38 3a 34 34 36 34 3e 43 41 3f 46 3c 40 3f 3e 33 3b 39 3b 36 34 2d 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 3c 44 4d 4f 4d 4f 54 4e 51 4b 53 55 44 52 4f 4c 53 4f 58 55 4c 50 4c 4d 49 4e 56 60 59 5b 5d 5a 52 50 55 5a 52 47 4f 51 4f 4d 4e 55 57 51 50 50 46 42 51 51 4b 46 4b 42 54 45 45 4e 56 44 4e 4e 4d 52 4b 51 4e 46 4e 49 58 49 51 42 52 4c 52 5a 55 54 56 5c 53 5a 5c 5e 54 4d 59 50 4f 54 53 55 49 4b 49 3b 44 3d 31 2d 1c 10 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 02 0b 0e 16 20 22 2f 3a 4f 53 4f 54 4f 44 48 46 3a 42 43 46 44 48 45 44 3e 46 41 45 39 46 45 42 49 41 44 43 3e 42 3f 43 4c 40 44 46 40 3e 3c 46 4d 3e 3f 45 43 41 3e 43 47 40 45 48 4a 41 48 43 3d 4d 45 40 3a 3d 43 34 3b 3e 35 41 3f 3d 3f 35 3d 37 3b 3f 39 37 37 3d 3c 37 40 35 37 38 35 39 3e 2e 3a 37 31 2d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 3c 45 53 55 47 57 4f 55 5f 51 56 4f 52 4c 52 4f 57 4d 54 4e 4f 4f 52 55 52 52 5d 4e 5b 58 54 52 50 44 4c 49 4e 4f 4d 54 47 4c 47 49 46 50 53 46 4b 3e 4b 4e 4c 49 49 49 4b 45 46 48 4d 43 4a 44 4c 46 50 44 50 43 4e 4f 48 4b 4e 4b 4d 4b 50 53 54 4d 50 52 54 59 55 5b 57 4b 54 4b 52 52 4a 48 50 41 40 3d 3a 37 20 1e 10 0f 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 1b 2e 1e 29 33 4d 4e 53 51 49 4b 44 40 3d 44 3e 46 3f 44 3b 38 44 45 4b 44 48 45 41 43 3b 4a 47
 3f 44 4e 3f 48 40 44 41 40 45 41 42 3b 48 46 47 3d 3f 41 49 3a 3e 39 3e 44 4c 3f 3b 44 3c 41 44 44 3c 3e 44 3c 39 37 3b 36 3d 45 42 3a 38 31 37 3b 3e 3c 3f 38 3f 35 3c 3e 36 3a 40 3b 38 3b 33 33 2e 1d 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 10 3f 43 4b 4c 4f 55 5e 5a 5a 52 5a 59 59 53 56 52 54 5a 59 56 52 57 59 58 53 54 53 4f 52 53 50 49 4f 4d 51 4e 4c 52 58 55 4b 43 45 48 47 41 4d 4e 4b 45 4b 45 44 4a 50 45 48 51 4e 52 47 4b 4e 4c 4c 45 43 4f 50 4c 4c 4f 4e 42 50 4b 4b 4d 54 54 57 55 4d 51 4f 5d 5c 5d 56 52 51 4c 51 4d 4f 4e 47 47 4a 38 36 2d 29 1f 16 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 14 0d 13 21 27 2e 3b 49 4d 4c 51 4a 4c 43 44 48 3e 3c 44 3f 3f 3f 3c 46 42 49 3c 47 42 43 48 40 48 48 46 40 4a 42 43 40 45 4b 45 42 43 47 43 43 41 45 41 48 3f 43 43 41 42 45 44 38 42 46 42 43 44 42 44 41 4c 43 3b 44 3e 45 4a 3a 41 3d 3a 37 43 35 30 30 3d 3f 42 41 40 3c 3c 37 3a 3d 2f 33 3a 36 34 36 24 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 3c 4d 51 4c 56 5d 5d 54 5b 57 5e 51 61 55 59 59 6c 5b 56 59 5a 52 55 55 57 5b 5f 5b 5c 4e 51 54 4c 4e 4a 47 48 50 56 51 4a 48 3e 49 44 44 4f 46 44 46 4b 40 49 4e 48 55 49 46 4d 4a 4c 41 4a 4a 4a 48 4c 52 4b 52 50 54 51 48 51 47 52 4b 52 4d 4e 51 55 55 5a 5f 5d 57 53 51 52 4f 4f 4f 46 49 49 4a 47 3c 33 3b 2f 1a 14 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0e 1c 18 25 39 40 49 4c 4d 46 3b 45 39 42 49 41 47 41 47 3e 44 3d 43 40 45 41 46 48 44 46 40 4b 49 3e 3f 44 42 45 46 47 3c 46 48 42 42 44 3e 3f 45 3d 4b 45 41 45 44 41 41 47 49 50 3d 36 3e 3e 45 43 40 41 3a 3c 3d 3d 49 39 33 39 39 41 3d 3f 37 3c 3e 37 34 34 35 32 35 38 3e 44 3b 3c 2f 39 34 31 1e 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3b 47 46 55 54 5a 58 51 55 57 5f 55 52 52 4f 52 57 57 55 4e 5a 4d 50 54 59 58 5d 57 52 47 4f 41 4c 51 4a 4e 4b 42 50 49 42 48 46 4b 4a 4b 49 43 4b 4b 47 50 4a 42 46 49 4f 41 44 41 4b 46 47 48 45 46 4e 4a 4c 49 4a 49 55 4b 4e 51 49 54 50 4c 55 4b 52 50 5a 60 5e 54 5b 52 4f 4a 44 4c 4e 45 3f 38 44 3f 39 33 21 1b 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 11 11 17 28 30 3c 44 4a 48 44 4b 50 42 48 3d 40 40 3f 40 43 42 39 44 3f 4d 3e 40 44 43 41 3f 3e
 3e 42 47 39 45 41 40 41 45 3f 42 44 3b 40 3f 42 50 43 3d 47 43 43 4a 42 4f 3e 3d 42 3f 3d 3e 3c 48 3b 3e 43 44 38 3e 44 40 36 42 35 33 3b 32 3e 38 34 3a 40 42 39 3a 3a 3f 35 34 39 38 39 30 38 34 38 25 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 37 48 4e 52 4f 4f 54 51 5a 4c 5d 5b 54 49 4d 50 50 58 4f 50 4b 49 55 49 4f 4f 50 51 52 4f 4e 4d 44 4c 45 3c 42 43 4a 4d 49 3b 43 51 43 47 47 3b 4b 46 3f 4d 42 4c 4a 4a 4c 41 4d 48 4a 49 49 50 49 47 4b 47 48 4c 51 43 4b 49 4b 4c 49 48 4c 5a 54 51 4b 56 54 59 5b 59 51 4d 4e 4d 53 4a 3f 49 45 3f 3e 3d 2e 2e 1a 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 08 0a 10 1f 22 1f 2a 42 39 42 48 4c 41 45 48 4e 3e 44 3f 4b 3a 3b 43 3a 43 44 4a 48 48 46 42 44 43 3e 45 48 41 47 44 43 42 43 3c 3f 43 3e 3f 46 40 43 40 3d 44 48 41 4d 4e 46 45 42 43 41 46 3c 3f 3c 41 3c 3c 3f 3e 3c 3d 41 3e 37 3c 41 3b 39 39 44 3a 40 38 3e 37 46 3a 38 34 3b 3a 3a 3c 3b 36 39 30 2a 21 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 33 4b 51 5d 53 5b 57 4d 50 49 4a 4b 49 4d 4d 4d 45 47 4f 47 4b 43 52 4d 59 45 45 52 50 4b 52 4d 50 4a 41 48 45 45 4a 43 4e 41 4d 41 49 4d 47 49 45 4f 48 44 48 4e 47 4e 45 45 4d 3e 4d 49 44 56 4b 3f 47 48 57 54 53 4c 49 43 4f 4a 4b 52 4b 4f 54 4e 4f 5a 58 54 52 53 56 54 4f 50 50 53 42 4a 44 3e 3c 39 32 2c 1f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 16 12 1f 26 2b 3d 40 41 49 42 41 4b 4b 49 43 3c 48 46 41 43 3b 46 43 46 48 41 4a 44 43 42 4b 3d 3d 4e 44 46 46 45 41 43 48 43 42 47 48 46 40 48 40 3b 3e 3e 3a 44 43 49 44 42 49 44 3f 41 3b 40 46 43 46 45 49 3c 38 3b 39 36 44 37 3c 35 38 3a 37 3c 3d 3d 38 3d 34 3c 38 35 37 39 38 34 37 39 35 30 2a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 26 4a 56 57 52 4c 4b 4a 51 4a 4b 4b 47 4d 42 47 47 43 4b 47 4c 42 4d 4a 4e 49 41 4d 4a 49 46 48 4e 40 4e 44 4d 45 4a 49 46 48 46 3b 44 46 48 48 47 41 3d 4e 49 4b 50 4b 44 49 48 49 46 48 41 3f 4b 48 56 45 4d 4b 4c 47 51 47 42 44 4a 59 4d 52 59 50 4a 51 4c 4e 4a 4a 4f 50 50 54 5b 4c 47 4b 40 3c 3d 35 33 23 1a 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 09 13 16 1e 26 36 47 40 45 48 3e 47 47 4b 48 46 3b 49 3c 41 3e 47 45 41 48 42 48 46 46 44 3e 45
 4c 47 40 44 40 47 43 44 3e 3c 44 49 3b 3c 43 4b 3f 44 43 47 3c 47 44 44 45 3f 41 45 44 3f 3e 41 3d 42 3d 43 3c 3a 3e 3e 3a 39 3e 39 37 35 37 3c 3b 33 3b 3b 37 3a 43 38 37 36 3b 3e 38 3e 2c 35 2e 32 31 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 18 42 44 50 50 44 4a 47 48 48 44 45 45 42 4b 3f 4f 3a 45 47 45 47 43 45 43 41 4c 44 43 46 48 44 42 3d 3f 4a 42 42 42 44 3f 48 3d 41 47 41 41 42 42 47 42 48 49 48 43 41 41 3f 4b 47 49 51 4b 4e 4e 43 44 3f 47 49 4f 4b 4b 4c 4b 46 53 52 4c 51 49 4d 53 51 51 52 54 54 4f 51 53 52 46 4b 46 49 47 40 37 30 27 27 14 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 0e 1d 19 2a 39 43 44 48 46 43 44 4d 4b 4a 48 44 45 3e 40 45 46 44 45 40 3e 46 46 42 44 46 4e 42 40 41 3f 3d 44 42 42 43 47 45 3d 39 45 48 46 47 3d 42 4d 42 3c 49 41 41 46 44 47 43 42 3f 49 43 44 3c 38 3e 3d 3c 40 3f 36 3d 39 37 3f 2e 3d 3b 35 35 3d 3d 3e 3f 36 30 39 32 3d 37 39 38 35 35 37 2c 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 40 3f 4b 44 41 45 49 4f 43 42 43 40 42 45 41 43 3f 46 3f 44 45 46 4b 3e 42 48 47 4b 44 54 3d 44 42 46 4a 48 43 41 44 3c 3f 44 48 49 48 4c 3d 49 45 49 4f 4a 49 4d 4c 51 47 46 47 4f 50 43 47 49 44 4d 45 4c 4f 50 4a 54 4b 4a 50 47 43 52 4e 55 4c 56 5d 56 57 58 49 56 4c 57 4e 4f 50 44 41 3c 35 3e 32 28 26 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 11 24 29 3a 3e 3c 4a 42 3f 47 3d 4b 44 49 41 3e 46 45 3e 3e 44 46 3d 45 43 42 43 3e 40 4a 4b 4f 3d 41 45 45 40 41 41 48 3e 47 47 45 48 45 48 45 43 48 3e 47 48 41 44 43 41 49 44 4b 4a 45 42 42 42 3b 3c 3a 3c 40 3e 36 3b 40 3b 41 32 3c 3b 36 36 3c 2e 40 36 3e 34 3a 3a 3a 3f 36 30 2a 30 2d 2c 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 35 42 42 40 45 44 44 46 43 42 47 45 3d 3e 39 44 3e 44 48 43 42 41 45 4b 40 43 49 44 41 4a 44 44 3f 48 40 4a 3b 46 45 3d 41 41 40 46 44 49 4c 45 48 46 4c 4a 41 47 4a 48 49 49 47 45 4e 4a 4a 47 41 52 4d 47 4f 4d 44 4e 4b 4f 4c 54 4d 4c 52 52 4a 55 53 56 5d 52 55 4e 4b 4d 4c 48 49 48 47 40 40 3b 2d 2e 19 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 18 1b 20 2a 3f 4d 42 40 46 48 46 46 4b 46 45 45 40 44 36 3a 3b 44 3e 3d 41 45 46 44 43 40
 3a 45 3b 3f 3c 3f 40 43 44 4c 44 44 44 45 43 41 3f 3e 4b 4a 42 44 46 40 3d 40 39 41 3d 44 3e 42 40 3b 3c 3f 3a 42 3d 43 3b 37 39 3c 35 39 38 39 39 31 39 35 39 38 33 35 37 38 3e 35 39 3b 3a 2f 33 29 35 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 2f 3c 45 44 49 3e 38 46 3a 42 3f 45 41 3c 42 42 48 46 41 47 48 44 41 41 3d 41 41 3e 44 44 37 47 41 3f 3d 44 41 41 42 43 3d 3e 48 40 45 45 4a 4a 47 45 3e 55 46 41 48 4b 43 47 48 4d 50 4c 46 40 45 41 4d 4a 49 4b 47 49 42 4a 4c 4c 4b 47 49 54 4e 52 52 52 4f 52 43 4f 51 49 52 49 49 41 40 40 31 37 31 17 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 10 13 1f 2d 38 43 47 44 44 3d 45 42 4b 40 42 46 45 41 48 3c 3e 44 42 40 48 48 3d 3e 3f 38 41 43 3a 3d 3c 3e 43 3d 46 3d 42 3f 3e 43 43 40 41 40 49 45 48 42 42 40 41 3f 47 43 40 43 47 3d 43 44 42 44 36 3d 40 40 3f 3c 42 3d 33 38 42 3a 44 35 3c 3c 3b 36 34 2e 34 41 3e 3c 3e 36 33 35 2d 27 31 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 33 38 42 44 45 46 47 44 3d 3e 4d 43 44 45 47 44 46 40 41 49 41 40 41 40 3e 41 37 3f 3b 3b 44 37 42 3c 47 46 38 3e 3d 47 3a 3a 45 42 46 42 4c 4d 50 4d 47 46 46 46 45 46 45 53 4c 4e 47 41 4b 44 43 4b 47 45 50 51 4b 4d 44 48 4f 4c 4a 50 4a 56 4d 4e 4e 53 4c 57 46 59 4f 48 47 45 50 44 49 46 34 2d 2c 16 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 11 13 18 2f 37 3d 47 45 41 3c 44 45 46 55 49 4b 48 3e 3b 40 3e 48 3e 3e 4a 42 47 48 3f 42 3e 45 3b 46 3f 3f 41 43 44 4d 3b 43 40 43 48 4a 46 44 45 3f 3e 49 40 40 44 42 49 41 40 39 3e 4a 3e 42 4b 3c 42 3d 3b 3a 3c 45 3b 43 37 37 3e 38 3c 41 39 3a 3a 41 3a 39 36 2f 3c 34 34 38 32 38 32 31 2d 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 2d 3b 40 44 46 4b 47 3f 3e 44 3d 44 44 46 42 3d 36 46 3c 44 42 47 46 45 3e 43 3b 41 3b 44 3e 3f 43 3e 41 3d 43 46 3d 43 43 44 4e 43 40 4a 46 46 45 43 48 49 47 45 43 49 40 48 4c 47 46 41 48 45 48 50 4a 46 48 58 4f 4e 49 4a 46 48 49 4a 45 4a 51 4f 4c 4f 52 52 4c 4f 45 52 4d 4b 46 45 3c 41 31 2b 1f 0e 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 12 12 24 29 37 49 4a 46 4a 4a 52 4b 43 42 40 47 3b 41 39 3d 44 3d 42 3a 41 3b 3a 3e 41
 48 3e 47 3f 45 44 3e 41 3d 39 45 48 40 3f 3e 41 50 3e 4b 44 45 3c 3f 46 42 46 45 3f 3c 3e 3c 3e 42 39 3e 3f 3a 3b 3b 3b 3c 44 46 3e 3a 34 36 38 35 33 39 37 37 40 34 34 31 32 2d 3f 38 33 2c 30 32 32 2d 1e 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 2f 38 41 41 42 45 45 47 46 47 40 46 44 41 39 44 44 38 41 3f 44 44 39 3d 37 42 43 3e 43 43 3d 3a 3c 41 3e 45 38 35 41 42 42 3d 49 48 4b 3e 4a 47 42 47 49 44 46 4f 41 45 47 46 3d 4d 42 4d 4a 45 4d 4d 45 48 3d 47 4b 46 45 4c 4f 4f 4b 4d 3e 50 4e 42 51 4f 4e 4b 51 4e 4c 4b 46 49 4a 49 3f 37 2d 27 14 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0f 13 0e 1b 29 2c 43 41 43 44 45 47 4b 44 4a 50 47 44 3b 42 43 44 3c 40 48 41 49 45 3e 3d 42 3d 45 43 3c 40 42 3e 3b 47 41 3d 44 47 43 44 45 45 4a 42 3c 49 46 46 47 3f 46 49 3b 40 48 3f 44 3f 41 41 41 3b 49 45 39 3a 40 3a 3f 3e 39 41 39 3d 3e 36 3b 40 35 39 3a 39 36 3c 37 36 38 30 34 30 2b 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 32 33 39 41 3e 44 3e 3b 37 46 40 3e 41 3e 40 43 45 49 3b 44 43 3d 3f 3e 3e 46 3e 43 41 45 3f 40 3f 47 44 3e 37 42 3e 3b 45 43 50 4c 4b 50 42 46 4a 43 48 4d 48 48 49 43 48 4f 48 50 45 40 51 4f 4d 46 42 46 56 4a 45 44 49 4c 4c 4e 49 4e 4d 4d 47 44 48 52 4c 49 4e 46 4c 4b 47 4b 48 3e 37 3f 28 22 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 09 0f 0e 24 22 30 42 3e 3f 48 48 49 4a 44 46 49 3d 3d 3b 3f 3e 3e 44 45 3e 41 3f 41 41 40 43 44 3e 45 3d 45 3c 42 3b 45 46 40 44 47 3f 4d 40 3e 42 4f 3b 3b 4d 44 47 50 3d 4a 44 40 3b 41 49 3d 4a 44 3b 3c 3b 40 42 3f 40 3d 37 3a 37 43 39 3c 3e 32 3a 3e 36 33 38 36 38 41 33 41 38 31 2f 2d 2a 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 2c 3e 3a 49 3e 46 3c 3d 3c 3f 46 41 41 3d 3f 3f 3d 41 42 46 40 3c 3b 40 39 45 3e 43 41 42 43 3f 49 49 44 47 3e 3f 47 44 3f 3b 45 45 45 49 47 42 4f 4b 4a 4a 45 41 4a 4a 3a 50 48 49 4e 44 47 4c 46 46 49 4a 4c 48 4b 46 4b 46 49 47 47 4b 50 4c 4b 4c 50 45 4d 49 47 47 48 46 47 45 42 41 41 36 28 18 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0b 0f 12 1f 2b 32 39 41 46 3d 45 45 4f 52 40 4b 42 46 3e 3a 43 3d 40 3b 3a 3a 41 43 40
 48 3d 3e 3d 46 45 40 3b 41 41 42 43 41 46 4a 46 45 44 42 44 39 4d 43 44 40 45 47 43 41 3e 49 42 39 41 3e 3f 48 3d 3b 41 3e 41 3e 43 3c 37 3d 3f 3c 34 39 3c 34 36 37 38 37 31 35 37 34 39 32 2f 2e 2a 29 21 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 33 42 42 40 3f 3b 3f 3b 3c 4a 3b 3d 45 39 3f 44 3e 47 41 3e 41 41 40 33 3b 42 48 39 46 40 3d 41 3d 3e 42 3c 3c 3f 42 46 42 47 4d 47 51 4a 48 44 4c 50 4b 4e 44 46 4b 45 46 4e 4c 4d 45 4d 43 41 4b 48 45 47 46 4f 46 45 48 49 43 4b 4d 48 54 4b 41 44 4a 40 48 53 4e 3e 4a 47 47 44 33 38 34 23 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 00 0a 06 0f 13 1b 2a 33 42 47 44 45 44 4a 4e 4c 50 46 45 3b 3f 3e 42 43 46 46 48 45 40 3b 43 49 4b 47 3a 3c 3f 40 42 40 40 44 3c 45 41 46 48 43 44 3b 4a 3f 4e 40 3e 3d 3e 3a 41 3d 42 39 41 41 3b 42 3e 42 43 40 42 40 34 46 37 40 43 40 3d 3d 3a 34 39 39 2f 36 33 3b 39 37 35 32 30 33 2c 2c 29 36 2b 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 24 3d 3e 43 42 46 3b 40 32 39 3b 3f 41 3e 3d 47 40 3e 38 3e 3f 41 37 40 40 45 3c 44 3e 41 3f 44 42 44 41 47 3e 3c 4a 46 48 43 4c 47 45 46 45 49 44 42 48 48 4e 46 47 4b 47 43 46 49 49 45 4b 44 44 49 46 44 52 4e 48 48 4b 4a 4c 42 45 4a 45 4e 48 4f 48 54 4a 49 45 46 47 44 45 43 44 3a 38 2a 19 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0a 06 11 14 1a 24 32 34 33 36 41 46 4f 50 4a 46 48 45 40 41 43 43 44 48 4f 46 43 44 4a 48 4a 4a 52 4a 41 3e 41 42 43 43 42 44 4a 3e 41 47 4b 40 44 42 45 40 44 41 3e 46 3b 45 3e 3e 41 42 46 3d 3e 44 43 3a 3e 40 43 44 3f 3d 45 39 34 3e 3d 40 36 3a 39 36 2f 32 3b 35 36 38 30 35 30 2b 2e 30 2a 22 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 3b 3b 44 3e 43 35 41 35 39 36 39 3f 44 3c 42 3b 37 42 43 4b 3c 47 46 3c 3d 3b 48 47 47 44 40 40 41 44 46 41 3e 4b 47 40 49 44 4a 4c 49 4d 46 42 4d 44 52 4b 4b 43 47 44 49 4d 4e 50 51 44 48 45 4b 4a 4d 42 4b 46 48 49 50 47 4d 4a 4b 46 4b 4c 4c 4b 49 4c 4b 4c 4a 4b 4a 46 43 3e 3e 32 2a 1a 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 15 18 25 33 39 35 3d 47 4b 4c 4e 3f 43 48 3e 41 3e 40 45 51 4d 44 4b 41 41 4d
 58 51 53 4f 41 43 48 44 49 49 49 45 46 41 40 47 4b 46 41 47 44 47 3a 3a 4b 41 42 3f 39 42 3e 3e 41 43 3a 3e 3a 40 3b 40 45 35 35 37 35 37 36 3e 33 3e 3a 34 40 30 38 41 37 39 32 34 3a 36 30 2f 2e 33 2e 26 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 31 45 35 37 36 37 3a 3f 3d 44 41 38 44 3d 44 39 3c 3e 41 44 3f 47 3f 41 46 3e 43 41 49 46 40 46 3e 42 41 3c 3b 3c 41 49 4e 44 49 45 44 46 45 4b 4a 49 4e 46 4e 47 44 44 4c 41 4b 45 41 47 41 44 42 48 44 44 44 41 40 41 3e 4d 43 46 4b 49 49 49 40 50 49 41 46 49 4a 45 44 45 46 40 38 33 24 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0e 0d 25 29 30 31 37 41 3c 45 4a 42 46 48 43 3f 3c 3d 44 4b 49 41 4d 3a 39 48 40 52 53 4e 49 4a 3d 47 46 40 47 43 4b 3d 4b 48 49 41 46 4a 41 43 42 47 42 45 40 36 3f 3b 3f 40 41 3f 3b 3e 3f 3d 3b 3b 3d 3e 35 42 3d 3b 43 37 3c 34 34 31 35 38 39 36 34 39 31 38 38 2f 2f 33 2b 34 27 2c 1d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 33 3c 39 38 38 32 34 36 3a 40 40 3a 3c 42 3b 41 41 49 40 3c 3d 3a 41 46 49 3e 3f 40 43 3f 3d 40 47 40 3b 41 3c 4a 45 46 3f 47 4a 47 47 50 4b 49 41 47 43 42 4e 4c 4b 4a 49 45 50 44 46 41 41 42 47 42 43 45 49 41 45 3a 49 3c 40 3c 4e 4c 4a 47 4f 41 49 50 4a 48 41 4b 49 49 43 3d 39 28 1d 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 07 10 14 19 22 31 34 3c 3b 41 43 44 4a 44 49 44 42 3e 45 42 41 4a 48 4a 47 44 3f 46 4b 56 56 50 49 46 44 43 42 46 4a 4c 40 4f 45 4c 47 40 4c 47 3c 46 42 41 49 3d 40 49 35 40 41 3f 43 43 3f 39 3a 34 41 3e 3c 3c 3c 38 31 41 3e 38 3e 3b 35 3d 2d 37 39 2f 32 39 3d 33 32 3a 35 31 32 33 31 29 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 17 34 44 3a 3e 41 3d 3c 31 3b 3e 39 40 3a 4b 47 44 3e 36 37 43 3a 43 44 3c 3d 36 3c 41 45 48 3f 3f 3f 40 41 41 3d 40 40 44 45 4e 4a 4d 46 43 46 47 48 4c 46 46 4b 4d 42 4a 45 45 47 43 42 44 47 42 4a 45 42 42 4b 47 46 3f 46 44 41 47 43 44 46 47 4a 49 51 4b 45 4e 46 44 43 4d 3b 3f 2e 1c 12 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 14 1e 24 36 36 35 40 3a 3d 48 49 48 43 3f 3d 3e 3c 4d 41 41 45 3e 36 3b 4a
 4a 57 4b 4d 46 47 38 43 43 3e 45 45 48 4b 4b 42 43 47 3e 41 46 44 47 41 40 3d 3b 41 40 41 43 43 37 41 3f 40 36 3b 3e 39 3b 33 3f 35 38 3c 37 38 3a 35 35 38 35 37 37 32 38 2f 37 2f 2c 34 32 32 33 2c 26 28 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 32 36 44 37 36 35 41 3a 3e 3b 3e 45 3f 42 37 41 3c 39 3f 3e 44 39 39 3a 40 3d 43 4a 37 41 3e 48 40 3d 44 37 43 43 3c 41 4b 42 4c 45 44 45 4e 46 44 47 4b 48 4a 42 49 44 3d 44 44 4a 44 47 3c 42 49 43 3d 47 3c 40 3e 48 42 3d 4d 3f 46 43 4b 4c 4b 46 40 48 46 4e 43 43 45 3f 39 3c 33 1b 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0a 18 16 22 32 2f 31 3e 40 46 42 49 45 44 40 43 39 3e 47 42 40 43 3d 45 3f 3a 4a 4f 54 51 47 4a 3b 3e 41 40 3e 40 44 48 40 3d 3d 3c 3c 47 45 43 46 36 40 41 41 3f 3e 3c 3d 43 40 3d 42 3f 38 3b 41 3a 3c 41 44 3c 39 38 3c 3a 32 36 35 3a 39 3b 3a 31 37 30 35 36 38 2c 30 30 30 2e 2a 1c 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1e 30 38 39 3b 40 37 3a 3a 42 42 3f 36 3f 47 3e 42 3b 36 40 37 45 39 40 3b 3b 43 42 40 44 35 3d 3e 39 34 42 43 41 3f 40 46 44 44 40 44 46 42 49 45 43 45 44 49 45 49 4c 41 41 3d 46 46 49 47 44 3e 3a 47 3f 3f 49 3d 41 3f 43 4d 40 48 4b 44 4b 44 43 48 42 4a 50 3d 44 48 3a 41 39 3c 18 17 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0a 09 1c 20 27 35 35 3a 3d 43 40 4b 48 43 38 3f 42 3a 3e 48 42 49 3e 3d 44 3f 4d 4d 4b 47 41 47 44 42 3c 3f 3d 41 3f 49 42 3e 45 3c 46 44 3f 43 42 40 44 4c 39 43 44 3a 41 3f 3b 38 39 41 38 38 3a 3d 3d 3a 34 34 44 38 3c 3f 40 36 38 36 39 3a 39 32 35 2f 40 39 39 2f 2d 2f 29 2e 2a 24 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 3b 41 33 3c 36 36 39 36 3b 3b 34 39 3e 3b 41 3d 3e 47 3b 3d 3e 36 40 3d 3a 45 3d 45 41 3b 3f 46 42 4a 48 45 3d 47 49 43 3d 40 41 46 47 41 47 48 44 4f 44 46 45 4b 45 47 3d 41 45 48 3f 45 42 44 47 42 43 48 47 48 3b 3e 42 39 41 41 3e 4a 45 4a 43 45 40 40 3f 45 46 42 48 49 3a 30 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 09 0c 13 1c 1e 29 2b 2f 3e 3d 48 48 44 3e 47 40 43 44 44 44 43 47 42 46 46 3b 4a
 44 4d 3e 3f 3b 49 3e 45 3f 44 35 3e 38 42 45 3b 42 43 3e 4d 46 3d 41 42 43 3c 41 42 3a 43 3e 48 49 3d 43 40 38 47 3f 3f 41 3b 35 40 42 3c 30 33 3a 36 39 38 35 35 35 29 3b 2c 31 34 34 39 34 2e 24 2c 2c 27 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 33 36 3f 3e 34 38 3e 34 3f 3d 42 41 39 3f 42 3b 3b 38 3b 3f 42 3d 48 39 44 3a 3a 35 43 35 35 3d 3c 40 3b 41 41 4a 46 42 41 40 46 3b 3f 48 2f 4f 49 3f 4a 3f 41 41 49 43 45 43 45 3f 42 47 43 3a 3f 3d 3f 46 46 3a 41 45 41 44 40 41 49 49 47 4a 45 45 43 46 4d 4b 44 40 43 3e 3e 28 17 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0a 17 11 1e 25 2c 36 42 35 3f 47 41 44 41 3f 3d 3e 37 43 48 4b 44 3e 3c 3d 44 3d 39 41 3b 41 3c 39 3f 3e 3e 45 3d 3a 42 3e 47 45 40 44 48 41 42 36 3f 3e 44 44 3c 3d 41 3c 3f 3b 3d 44 3f 39 35 3b 3d 3e 38 38 3c 36 34 3e 3d 3a 2f 3a 32 34 32 2b 31 39 37 3a 32 2b 2e 2d 2d 26 2a 27 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 28 34 3c 37 35 3a 32 30 38 3b 32 38 38 3e 40 3a 3b 3c 40 40 3c 3d 34 36 3b 3b 38 3b 3c 3c 40 32 3e 3c 44 3a 3e 45 3b 3f 49 3f 40 46 40 47 4b 3b 3f 42 41 38 42 3b 44 47 42 3f 48 45 42 47 4b 3f 40 3e 3c 3b 42 37 46 3d 3d 42 40 45 45 47 46 44 44 47 4a 4c 42 40 3f 45 49 42 2c 1d 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 0c 1f 20 1f 30 39 42 40 39 43 40 3d 43 39 43 3e 48 48 45 48 4a 3f 43 40 3a 3f 42 3c 3b 47 3e 43 3c 42 41 40 38 3f 3b 41 46 48 40 3f 42 47 45 41 3d 3f 41 3a 40 43 47 3d 3e 3e 3e 44 3e 3d 42 3b 39 3c 31 43 3e 36 33 35 3c 35 37 39 3a 38 34 39 30 34 32 31 2b 33 30 30 2a 25 25 2c 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 29 38 39 37 38 39 38 35 30 3d 34 42 38 31 3f 3a 3e 40 3b 3d 36 3e 3c 39 41 36 41 37 3d 32 38 38 3f 3b 43 47 44 45 41 3b 41 44 3d 41 39 42 40 3c 45 41 49 47 3e 48 43 42 4c 42 44 41 3b 3c 3f 40 39 37 3b 46 3f 3f 40 40 3b 45 44 40 44 41 4b 45 47 51 41 47 48 44 40 46 42 37 31 1b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0c 10 17 1e 21 2b 2c 36 39 41 3b 45 44 42 44 45 4b 45 47 47 51 50 46 47 3c
 3d 41 40 3c 3b 41 3a 3e 3b 41 3d 44 44 3c 3b 3e 42 3e 3d 44 3b 42 45 40 47 3b 3e 3e 40 45 4a 46 3f 42 3f 48 3b 3a 36 40 3b 35 39 40 40 42 33 3a 39 39 32 3d 3d 34 3a 3c 34 30 3e 30 35 34 34 2b 2b 2e 22 24 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 28 35 35 31 32 32 41 38 34 3a 34 38 3b 36 3a 3c 3e 36 3a 37 37 3a 3e 39 3c 36 3c 38 39 3e 2e 3c 44 41 42 3e 40 42 3c 47 43 3e 3d 39 41 3e 48 43 45 44 3c 44 46 41 40 42 45 41 40 49 3a 3b 3b 38 41 41 41 3b 3c 3d 3e 3b 42 41 40 42 4a 46 40 45 4f 4d 46 51 44 40 45 3b 41 34 22 10 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 0d 0f 13 18 2b 30 32 31 40 3d 3c 42 44 3d 34 3f 44 3c 49 43 44 43 3d 3a 40 3b 43 38 3f 3b 36 42 44 41 39 44 37 37 3d 3f 3a 3c 3e 4b 39 3f 43 35 3e 3a 3d 38 3d 37 3a 43 48 3b 38 42 39 36 3d 3a 3c 33 3f 37 38 3d 32 3d 39 3b 2e 33 37 39 37 36 3b 34 34 35 34 32 31 3b 2d 2e 22 27 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 21 25 31 41 36 36 37 32 38 3a 38 2f 39 35 37 38 38 36 32 3c 36 34 3b 3d 3a 39 3a 39 37 31 39 33 36 3c 35 41 3e 3b 3e 37 39 3f 42 41 3c 3d 40 41 3b 3f 3c 46 41 42 3b 3f 3d 36 3c 3f 40 47 43 3b 40 36 3e 44 42 36 3e 3d 3a 37 4b 45 43 42 42 49 46 41 44 41 42 49 42 3c 34 27 1b 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 13 1a 1c 23 26 25 33 2e 41 3f 42 45 42 45 41 4b 44 48 4f 3d 4a 43 46 42 44 41 3e 47 3a 3e 34 35 4d 43 44 3f 3c 40 3f 3e 3d 44 41 44 33 3d 3d 41 3a 47 48 46 39 3e 3d 3e 3b 3f 44 32 3a 36 33 34 3b 39 3f 34 3c 35 3e 33 34 3f 37 36 3d 3c 38 35 31 39 37 39 33 2e 32 2a 28 2c 2b 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 25 36 37 3c 32 32 39 33 3d 37 3f 34 39 3d 41 35 3e 31 38 3e 35 3c 34 39 32 31 3f 3c 43 33 3c 3e 33 3c 41 3b 42 35 43 3b 3b 42 42 44 31 3f 3b 3f 41 47 41 3f 4a 42 48 42 3d 3b 43 3e 3d 3b 41 39 36 35 40 38 41 42 3f 41 3b 3e 39 42 3f 45 40 3a 41 4a 49 4c 46 43 43 2f 30 1e 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 0d 1c 20 27 2c 25 2e 25 43 40 3a 3c 3e 42 43 47 45 3f 44 44 3b 3f 45
 47 43 47 3e 3d 3f 3a 42 38 36 3d 3f 38 44 42 41 3f 40 45 46 3d 43 42 44 3a 45 3d 3f 3b 35 41 3e 41 40 42 41 3d 3e 3b 3f 44 41 41 39 3c 42 30 3a 3b 3a 35 3e 38 3a 3d 38 3a 36 2d 36 33 32 36 39 35 2b 2e 20 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 28 3d 39 36 37 36 3b 35 41 32 3e 3b 38 3a 3b 35 3b 40 3b 42 35 3a 3f 36 3d 3a 37 3b 3c 30 3c 3e 35 3e 3a 3a 3b 3e 43 3f 3d 3b 38 3a 37 3d 3d 3f 47 3b 3d 46 3b 42 4a 44 39 47 42 3f 38 3d 40 36 3b 3e 3c 3d 3f 39 3b 3d 3b 4d 40 41 49 3a 49 41 4a 43 46 4c 49 3d 45 39 23 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 13 10 19 1b 21 27 2b 2f 32 35 37 46 3a 43 45 3e 49 42 40 3c 3e 42 40 43 48 3e 42 40 37 36 35 3c 36 38 35 39 43 41 39 40 41 3e 3f 41 33 42 45 49 47 44 47 3e 41 40 3e 3e 47 43 3c 39 3c 3b 3f 41 37 37 38 3c 3b 3c 39 35 35 34 3c 3c 39 3c 37 30 3c 2a 38 30 31 31 31 32 2d 30 27 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 37 38 3b 33 37 32 27 3e 39 34 32 37 3a 3d 31 2f 30 39 3c 39 35 3c 3c 3c 3a 41 34 33 36 34 36 2f 3b 44 38 3a 3a 3f 3b 3c 35 3d 41 42 40 3c 3d 3c 45 40 3d 3f 43 45 3c 3c 40 45 3e 49 39 40 3c 3e 3f 3b 3b 3e 33 34 38 3f 36 35 3b 44 48 43 3f 42 42 3f 42 38 41 37 26 20 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 09 0f 1c 26 25 28 33 36 38 39 35 43 3a 3e 3f 42 42 46 3c 39 41 3d 44 49 40 42 3b 3e 34 41 38 3f 3e 44 3b 3b 3e 3d 3d 3f 49 38 3d 3d 32 42 3f 3f 3f 3f 40 44 43 47 3f 45 3e 40 3f 45 3b 3f 41 37 3c 43 36 3b 3e 37 3a 30 31 38 35 39 35 37 39 39 3c 3f 2c 38 2d 33 35 2a 27 2a 21 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 24 3e 37 33 36 37 33 3d 3a 38 31 2e 30 3e 38 37 33 3a 32 34 37 35 35 34 3d 39 41 3c 34 38 2d 34 38 3f 3b 3a 3e 3a 39 39 3d 44 43 48 39 38 41 35 38 3b 47 39 3a 47 42 41 41 3a 3b 3e 35 3a 3a 3c 3b 3a 37 3a 40 39 2e 38 40 3c 3d 3e 42 39 42 48 40 4a 45 47 3e 3d 39 22 10 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 09 0d 23 1b 1f 24 29 2c 34 33 3e 3d 39 4d 4c 3d 44 48 40 3b 43 44
 43 47 42 3f 3b 37 3e 3f 3b 3f 36 3c 39 43 40 3f 45 42 3e 41 47 3a 3c 42 3d 40 49 44 41 44 3e 3b 41 40 42 45 3f 40 3c 3a 43 3e 3c 3e 33 40 32 38 44 38 38 40 40 38 32 3b 31 39 33 30 2f 30 36 34 3e 32 34 28 1c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 31 37 38 3f 35 3d 3f 3d 38 34 3c 3c 3f 38 36 39 38 3a 35 40 33 3a 34 30 2b 33 38 32 38 35 35 43 39 38 44 35 3f 3d 37 41 38 3a 41 40 3c 45 3d 3f 3c 42 3f 44 47 3b 3e 37 3d 44 3f 3d 3f 42 3a 3e 3a 3c 3a 37 36 43 40 41 44 3c 3f 40 45 40 40 40 49 46 42 42 36 2d 1e 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0d 14 1f 22 22 2a 35 34 35 35 37 44 41 46 47 40 44 3d 42 42 45 3b 45 47 3e 44 3e 38 3a 3c 39 39 39 35 43 3e 38 41 3d 43 42 38 3f 3c 40 3c 45 3b 42 45 4b 45 3e 3e 44 40 3a 3c 3b 3f 3e 44 3a 3d 39 37 3f 32 37 3b 37 35 3f 2f 36 40 33 36 37 35 38 2c 36 35 30 34 2f 29 2f 1f 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 17 34 2e 3d 32 31 39 36 35 3e 3e 3c 39 37 26 35 33 35 3b 32 39 33 32 3c 3e 35 44 36 38 34 36 3e 3d 3e 3c 3c 39 30 37 3c 41 42 35 38 38 41 40 3c 3b 43 3a 40 3e 41 3d 3c 41 3a 3e 3e 39 2f 41 33 43 42 3c 3e 34 3b 3d 41 48 3f 40 3f 3c 3e 42 40 4a 4e 4b 45 33 31 1d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0e 1f 21 2b 24 30 35 34 34 39 3e 38 3c 3b 3f 44 40 3e 40 3e 41 4d 49 40 40 3b 38 37 41 34 39 43 3c 3a 38 3b 40 3b 41 44 3e 39 43 44 40 36 3b 42 40 42 41 3c 3e 3b 3b 45 3d 3d 39 3a 3e 39 3a 3a 3a 3d 31 39 33 31 33 30 34 34 36 35 39 2f 36 3b 30 33 37 2e 2c 2a 30 2b 1e 0c 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 31 35 3a 3b 35 3c 39 3d 36 3c 2e 30 2d 37 32 31 38 35 39 34 30 38 3c 35 37 36 2f 34 38 33 34 3d 3b 31 37 38 3d 35 3a 3d 32 3d 40 3d 3a 38 3c 3f 3e 3e 3d 3a 3b 36 3a 39 39 41 3f 3e 42 3c 39 3b 36 3a 41 38 40 39 2d 39 40 3a 39 43 40 48 44 3d 40 41 36 3c 2b 11 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 0b 17 23 20 20 27 2f 32 32 34 3f 41 3f 40 3a 43 40 3c 3d 45
 3e 4a 4d 44 3c 3d 3c 36 3b 3d 42 44 39 41 3a 38 46 3e 44 44 3d 42 3c 39 46 44 47 43 41 3d 41 49 49 46 4a 41 45 3e 3b 43 38 39 3f 37 3e 37 33 39 3e 3d 3c 3b 35 32 2e 36 2c 36 37 37 2f 36 37 35 2e 2f 36 29 21 07 06 05 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 35 39 3d 35 2e 37 2e 34 3e 36 37 38 3e 3b 33 35 34 39 33 38 39 37 34 34 30 3e 34 30 2e 2e 3b 30 35 37 3b 37 34 33 41 36 3d 3d 36 30 3b 3f 3b 40 38 38 42 3b 36 39 38 35 43 38 36 3b 3e 3b 3c 3a 3b 3e 46 37 38 3c 35 39 39 40 39 42 44 42 3f 3b 42 44 45 2a 1f 14 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 18 1a 23 29 27 35 34 36 33 36 3e 3f 3c 43 45 3b 4a 3e 40 40 44 46 4a 3f 43 40 40 3c 3e 3a 40 3d 3f 3d 41 37 38 3b 43 3b 3a 49 3c 45 40 40 3e 3c 49 44 45 49 3e 3e 45 3a 3f 41 3e 3d 38 41 3c 3b 39 3d 42 3c 42 3f 35 3b 39 3b 30 34 34 34 3b 34 3a 32 32 32 31 32 29 28 05 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 37 35 3b 31 35 39 2e 32 32 32 39 3a 32 37 38 31 34 3a 26 30 35 35 38 2c 35 39 37 37 39 31 3c 34 38 3a 36 36 35 40 38 2b 40 39 42 38 33 3c 40 32 43 36 3f 41 37 3e 3b 3d 37 3e 46 36 3f 40 32 35 38 34 3b 3b 46 3b 39 3c 36 3d 45 43 44 45 3e 4f 3f 41 38 23 1f 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 10 1b 29 20 24 2c 33 2f 38 3e 36 38 3a 3a 43 40 42 41 42 45 44 3f 45 3d 36 32 3e 38 43 3d 3b 3a 3d 44 3e 3b 37 3f 42 44 42 3c 3c 39 38 43 44 40 44 43 46 44 45 43 3e 3d 42 40 3b 3e 3f 3d 43 3b 39 39 41 3a 36 32 2d 30 35 36 38 2f 32 31 32 39 32 3b 34 2f 2b 2e 25 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 33 34 33 33 33 38 32 3c 31 2e 37 35 2b 39 34 39 35 38 35 32 35 34 2d 2f 32 38 3b 38 2d 3a 2d 37 33 31 3d 32 39 30 36 36 37 36 38 3d 41 3e 31 39 39 32 3a 36 3c 3b 36 41 3e 42 3f 3e 36 36 33 3b 43 44 3c 38 2b 44 34 34 44 34 46 41 48 49 45 4b 3f 3f 35 24 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 10 1c 1a 2d 27 27 2f 2c 35 3c 3a 43 44 3f 38 3f 39 39
 3f 45 41 40 39 41 39 3f 37 3b 3e 3d 3b 3b 36 40 3d 3e 3f 3e 40 42 39 41 3d 3b 42 41 3c 42 41 47 48 43 4a 4d 43 46 46 3d 47 36 44 42 3a 3c 38 40 47 42 3f 37 35 35 34 3a 34 2f 35 35 31 3d 32 34 2e 29 33 30 28 11 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 2b 2e 3b 32 32 3e 2e 30 38 39 35 33 36 34 39 31 2d 35 32 3b 34 35 33 30 39 34 37 3a 32 37 37 3a 37 3b 3d 3b 37 35 39 37 39 35 40 3c 40 3d 3e 3e 3a 40 36 35 3d 3d 35 3b 3f 3c 3c 3d 35 3a 37 34 36 39 40 3b 35 35 33 3b 3b 3f 46 3f 42 3a 22 35 3c 3f 2e 19 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 12 17 28 20 25 2e 2d 2e 34 36 3d 3f 2f 40 3c 35 44 3d 3f 40 48 3d 36 3e 3f 3d 3a 44 3a 39 3b 34 43 3b 37 3f 36 3c 39 44 41 3d 38 40 42 44 3c 42 3f 41 4c 4b 44 4d 4f 4b 47 46 41 3e 42 36 3d 44 42 41 41 41 41 3d 32 36 30 2f 37 3a 2e 2f 34 36 2b 2f 34 33 2d 27 29 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 26 30 37 36 39 38 2c 2c 38 33 35 3b 33 37 2a 30 31 35 36 36 35 29 2e 30 32 34 2f 38 36 34 35 2e 36 33 3b 33 37 3b 3f 41 3f 35 3c 39 37 3c 36 33 3d 3c 35 39 38 36 35 43 35 47 38 40 35 3c 36 3e 3f 3f 49 37 33 3f 3a 3c 3e 40 3a 45 40 45 3f 3c 2e 33 1f 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 18 20 21 1f 25 2f 31 30 37 39 3f 46 40 3d 42 41 42 3f 41 3c 40 3f 3f 39 3f 38 37 3d 37 40 43 35 3b 34 42 3f 3f 39 2e 3e 3f 46 3d 37 41 3c 41 43 46 4a 4c 4b 54 4b 43 45 43 46 44 49 48 3e 44 44 4c 42 3c 36 31 30 35 2f 25 2c 33 35 2b 35 39 2d 30 30 2e 2e 25 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 2e 36 36 2f 32 33 30 3a 35 34 27 31 35 31 32 2f 32 2e 2a 32 30 32 30 30 34 38 33 36 34 35 2f 37 36 38 39 36 3e 3c 3e 34 30 36 3a 3a 3f 41 3c 40 34 3a 44 3c 39 32 32 39 39 3d 39 3b 45 3e 3a 3f 40 46 44 47 41 42 3e 3e 43 42 49 3a 43 3e 39 3d 29 1f 10 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 13 1f 25 2a 2c 23 27 36 30 3f 3d 3b 3d 3c 43 41
 42 43 35 3b 3e 41 38 37 3f 44 41 3e 3f 41 3b 3b 37 3a 41 3b 3a 3b 3c 41 47 3d 3f 3b 33 3f 3f 46 4c 45 4e 54 54 4c 4b 54 3e 44 46 46 43 42 44 46 51 4b 4b 3a 3b 36 31 38 2f 2c 34 30 32 36 31 34 2f 31 2d 26 29 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 23 2e 34 32 28 3c 34 38 36 36 35 30 3a 31 35 30 30 35 35 36 32 2c 33 31 2b 39 37 36 32 35 34 38 37 3b 3d 35 38 31 32 38 37 3b 3c 38 3e 35 3c 33 36 39 42 3d 3d 46 3a 48 3c 3f 3c 3b 3e 43 44 45 47 44 48 51 53 49 45 4b 43 47 49 3c 44 3f 39 33 22 15 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1a 1c 1b 20 2b 29 33 33 35 37 43 3e 42 41 38 39 35 35 3d 42 3b 3d 40 34 3d 3b 3b 39 3a 38 39 32 3e 35 3b 36 3b 3e 41 40 3a 43 3c 42 41 43 47 46 47 4f 56 47 50 50 4b 45 4e 4d 4e 49 56 49 52 4e 49 4c 42 35 3b 2f 34 34 2f 32 32 33 2b 2a 38 28 31 2e 31 25 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 22 36 36 30 2e 33 32 31 37 2f 33 37 31 35 31 35 35 36 35 35 32 37 36 2f 2e 2f 32 3b 36 34 32 33 35 41 37 34 33 36 3c 3a 3b 38 35 3c 37 38 38 39 3c 3e 3a 3e 39 37 31 3e 40 49 44 41 4b 49 4d 59 58 5d 5e 5e 55 5a 4f 54 45 48 40 44 47 39 33 2f 15 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 14 20 21 22 24 2a 2a 2a 2f 34 3e 3d 45 47 3b 43 3d 3a 39 3d 39 38 39 3a 3e 32 3a 3a 39 42 35 31 39 39 3e 39 43 41 3b 46 43 45 3f 3f 40 3a 48 44 50 47 4d 54 4a 4b 53 4a 4d 51 4f 52 53 52 58 56 4d 48 3e 3c 31 35 31 30 2b 36 32 2e 32 2c 2c 2e 2a 30 29 29 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 1d 34 32 2f 32 37 32 37 32 34 39 38 32 32 30 32 31 30 35 2f 2f 33 2f 36 2f 33 35 31 34 2c 32 34 2d 3b 35 31 30 31 35 33 33 39 3b 37 38 38 32 31 3b 3b 3e 2c 38 38 3d 3b 40 3f 48 4a 57 5c 60 60 70 6d 6b 6d 63 6a 5e 5b 5c 45 45 3d 3c 39 2f 1b 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 14 16 25 25 2c 28 2c 31 34 3b 49 48 41 3e
 44 3a 40 44 31 42 3c 41 3e 46 3a 3d 3c 3d 39 3f 38 36 39 40 37 3d 38 3f 42 47 41 3d 3c 44 41 49 41 45 4d 57 4c 52 57 54 59 50 54 52 4e 59 56 5c 60 4f 4f 43 36 35 36 39 32 2b 35 36 3c 2e 2e 2c 2c 30 2a 2a 22 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 39 3a 32 30 36 2a 33 39 36 2f 34 2e 32 2f 36 36 3c 30 37 2f 2e 37 39 2a 33 2a 36 30 32 33 2f 33 39 36 36 36 33 35 3b 34 33 3b 39 36 35 35 3a 39 34 3b 38 3b 3e 40 45 46 59 62 63 6b 66 6e 79 7c 72 7d 7a 73 78 68 5f 57 49 40 3e 3c 33 1c 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 19 22 25 2a 27 2f 2d 32 3e 3b 42 3a 3f 39 43 41 3d 3e 3e 3d 3f 40 41 3e 3b 40 40 38 44 3b 39 3c 3a 37 3b 40 3f 49 41 43 3c 40 45 44 4b 51 52 53 4f 57 57 57 4f 52 50 55 59 5b 5b 58 5a 5e 56 46 43 42 34 39 32 39 32 32 38 36 39 30 2d 30 2e 27 2a 2a 21 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1c 37 36 36 28 37 2e 2d 2e 32 33 2b 3b 35 28 2f 38 30 34 35 33 39 39 30 32 35 33 2f 34 2b 32 3a 2d 32 31 38 2c 37 38 37 3d 43 3c 37 2e 38 37 37 3a 39 41 40 3e 46 4d 4f 5a 66 71 74 7c 77 7e 7f 79 7b 7d 80 81 73 63 6c 59 43 43 3c 35 28 0f 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 10 20 28 26 29 2a 30 32 38 39 36 3a 3f 4b 39 42 39 44 41 39 3e 41 3b 3d 38 42 36 37 30 3b 35 3b 3a 38 3e 3f 3f 45 38 3e 3f 3c 42 4b 4b 4e 4f 54 5c 59 54 5a 52 4b 4c 59 56 5b 64 66 5d 50 43 3d 3b 41 33 30 3b 2f 2c 29 33 32 31 2e 2c 27 27 29 26 16 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 16 26 33 3a 31 37 2c 30 2d 2d 30 33 36 34 2e 2a 31 34 33 32 2b 33 30 31 2e 31 33 35 2c 2b 2c 36 34 36 33 37 2e 3c 33 30 36 36 37 32 37 3b 3b 39 3c 3c 3f 41 47 57 5e 62 6b 6f 74 71 7a 81 78 79 7f 75 7e 8a 7d 76 6b 64 5b 48 3c 33 27 18 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 13 1d 20 27 2a 33 32 35 3a 36 44 3d
 3c 42 41 45 3f 41 3a 40 3d 40 3b 36 3a 3e 3e 3e 37 38 43 37 3f 3e 37 3b 41 3b 36 36 36 42 4b 4a 4c 4d 52 59 63 64 57 51 53 52 57 60 5b 5e 54 63 62 58 52 49 37 3c 32 35 37 35 2b 2a 2f 30 32 31 2e 2c 28 33 20 1d 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 29 30 35 2f 3a 34 31 35 33 33 2b 31 28 33 34 31 2e 35 2c 25 29 36 36 2d 2e 2a 35 32 2d 31 38 37 39 39 39 3f 3c 31 31 39 3c 33 31 44 35 31 3b 42 46 48 50 60 6a 6d 74 78 76 7d 79 80 73 7a 78 6e 73 72 78 7c 73 64 60 53 48 3b 28 1d 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0c 13 25 18 2b 25 27 38 36 39 42 3d 44 4d 4b 45 43 42 38 44 3f 46 40 36 3c 3e 34 35 3d 34 34 3d 36 3c 36 3f 3c 35 38 39 42 45 46 45 49 58 58 61 5d 64 60 59 5f 57 5e 59 5a 66 69 64 66 54 48 42 39 36 37 34 32 36 35 37 33 35 32 25 30 2a 2a 2a 28 1f 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 2c 36 39 30 36 31 2e 35 36 2a 3a 2d 33 31 2d 2f 33 2d 2f 31 2c 2c 2d 34 36 2c 29 2e 36 33 35 39 35 2d 31 30 2a 3d 38 36 3a 37 35 42 39 3d 46 48 51 58 69 6e 73 79 75 7e 76 81 7d 7d 5c 75 74 75 77 7d 71 75 72 65 57 4a 41 32 20 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 14 15 20 21 29 2b 2a 32 2f 36 35 4a 4a 49 50 4a 48 43 39 3b 40 3a 44 3d 3f 38 42 34 42 37 36 32 34 37 34 38 43 3a 40 39 3d 41 4a 48 52 59 58 4e 63 59 5c 55 54 5c 60 61 5f 68 60 5c 51 47 45 38 39 3a 2d 33 2d 29 30 31 2d 20 25 2d 2c 34 29 2b 1d 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 2c 30 31 29 36 24 3e 36 2a 2f 2d 2f 37 39 32 2f 30 30 2d 2b 31 35 2d 2d 35 2c 31 39 2f 39 36 32 34 33 2c 3b 2f 35 31 35 33 35 31 39 45 4b 4e 5b 63 66 73 6c 73 75 71 74 7b 6f 74 7a 74 7b 78 6f 70 71 6e 67 6b 57 4c 3a 2c 1e 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 12 23 1e 1f 23 33 2c 35 36 3e
 41 50 53 50 4c 47 43 40 3f 3c 43 3e 42 3c 3d 36 31 3a 36 39 3d 3c 3c 35 32 33 39 3d 3d 43 41 48 4a 53 5b 63 5d 58 57 5a 58 61 59 54 5a 5a 67 64 5b 4d 48 3a 3a 39 36 2d 31 32 36 3a 2c 29 2e 2a 29 2c 2a 27 20 24 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 2e 33 31 27 29 33 2e 27 30 29 29 31 28 2c 36 2a 2a 32 2a 34 36 2f 30 29 31 29 35 2f 2e 2f 34 31 30 3a 31 39 3c 38 38 2f 3f 43 43 4b 49 52 5d 69 72 70 7b 75 78 71 72 78 72 73 69 79 6a 73 72 6c 66 6c 68 65 57 4e 42 33 2c 14 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 19 1c 28 1f 2c 2d 30 35 33 44 42 51 4e 4f 54 4e 46 4e 45 3c 3b 41 3c 42 44 36 36 37 40 37 3c 3a 39 3b 3b 3e 3a 36 3d 42 51 4e 50 59 5e 5d 5c 5f 59 5a 51 5c 5b 5a 64 68 5f 57 48 40 38 36 36 32 26 30 30 38 35 2b 2e 27 2b 29 2a 27 26 2a 29 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 27 32 3a 31 2a 2e 31 2d 2a 2f 2f 2f 2f 2e 29 32 2e 32 1f 31 2d 2e 31 35 2f 3b 31 23 35 2f 3a 31 33 34 34 34 36 36 3d 33 3d 47 41 5e 5c 61 6f 71 76 77 72 77 77 7b 76 6b 76 6c 6f 6d 6b 6a 71 70 68 6c 63 5e 54 45 36 28 18 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 14 1f 1f 20 29 2d 30 33 3e 46 54 52 54 5e 54 54 47 3f 40 3d 3f 3e 42 42 3b 3e 3d 3e 35 3c 30 37 3c 36 3a 37 3b 3b 43 48 50 52 5e 5d 54 5a 56 59 5c 57 54 5e 5b 5b 5f 5e 56 4c 3b 36 33 31 36 31 2f 2d 34 30 28 34 28 25 2d 25 23 27 1c 26 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 24 31 2d 2d 31 29 2c 2e 24 2d 31 2a 2d 2a 2a 27 2d 2d 2c 2c 2c 24 2e 35 2e 30 2d 2e 32 2f 32 32 36 31 2f 31 2d 32 36 39 44 4e 54 65 6a 6c 70 76 70 6a 70 6c 68 6b 68 65 6c 6a 66 64 6e 5b 5e 61 5e 6e 59 56 46 33 24 17 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1a 1b 24 20 21 2b 2f
 3b 3f 3f 50 50 52 52 53 56 50 40 3f 3d 39 36 41 3a 45 39 3b 3b 3d 3e 31 38 32 32 3a 3e 34 39 50 4b 50 56 60 5e 5a 51 51 54 52 50 56 59 63 56 59 48 41 34 2a 2f 30 2d 2c 31 2e 28 30 2f 31 27 30 23 21 26 27 29 21 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 24 23 2f 2d 2a 22 2c 27 1b 2b 2d 24 2f 29 20 23 25 2a 23 2b 36 1f 2b 2e 2e 24 2d 24 23 2a 27 30 33 28 2b 31 3a 3c 39 50 55 5f 60 65 72 67 6f 6c 6a 68 66 62 62 65 62 5e 67 67 57 5b 5a 63 63 61 5b 52 4c 3b 36 15 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0b 0e 17 23 26 2b 2c 33 31 38 43 4a 4f 5b 55 55 59 51 4c 40 3a 46 3b 36 3f 3d 37 3d 31 3a 3d 3b 37 38 35 3d 47 45 4a 3d 44 49 5a 5a 52 4f 55 57 51 50 55 51 4f 5c 56 55 48 3a 30 2c 2d 2f 2c 27 32 25 31 2e 25 2c 27 2d 23 28 25 27 27 1d 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1e 25 24 35 2c 28 29 28 26 24 2c 2c 30 22 29 1e 24 25 29 2c 28 25 29 27 25 2a 2c 28 29 2a 2e 2f 2b 2b 30 2c 33 4e 4b 5a 56 61 67 62 5e 62 68 68 66 61 5f 5e 60 55 5d 5c 5b 52 53 55 5a 53 5e 5a 47 4b 3d 29 1b 0b 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 15 1a 21 1e 22 28 2e 37 35 44 4d 4f 49 4d 54 5b 47 40 40 43 3d 3e 3c 3b 3f 3d 33 3b 37 36 3b 35 32 3e 3d 36 41 48 51 47 4d 53 51 52 51 49 49 46 4b 4f 51 50 45 43 42 34 29 2c 28 2f 2b 2c 2e 30 21 2c 25 27 2b 22 23 20 29 24 1b 21 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 23 1d 1c 1f 1e 1f 19 17 1e 1c 28 1d 1b 1f 25 1c 17 1c 22 24 22 25 1d 25 24 23 21 1c 1e 24 2e 26 29 2f 38 45 4d 4a 54 51 54 53 55 51 4e 4e 4d 4c 4a 4e 53 4a 49 53 52 4e 4f 50 4e 55 45 43 44 3e 37 28 19 08 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 13 14 21 21 21
 31 33 2d 34 3b 46 4c 4b 4b 4e 45 41 37 3a 3d 3a 37 38 3a 3a 39 38 35 2b 32 37 36 35 3e 32 39 43 4c 41 48 4e 40 44 44 42 4a 44 44 49 43 45 34 39 2e 26 25 24 25 29 2b 25 28 1f 24 25 18 22 24 24 20 1b 1a 1e 17 14 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 19 12 15 11 0c 17 13 16 13 15 16 10 0e 11 0f 0e 09 1e 18 11 18 15 15 0c 1c 1b 14 13 0e 1b 19 1b 24 27 2f 2f 34 35 38 3b 3f 3d 42 3b 45 36 38 39 36 3a 37 36 39 35 36 36 41 38 3d 3c 38 36 38 31 25 16 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 0b 20 23 24 24 27 2d 33 3f 43 3e 45 48 48 49 42 35 39 3b 41 39 34 41 37 39 35 37 33 35 3b 33 34 35 32 35 43 3f 3a 4a 45 4e 46 3d 44 46 40 40 44 39 38 2c 31 27 20 1e 23 28 1f 24 27 1c 25 1f 20 1b 20 22 1b 15 15 14 10 13 10 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 07 06 05 06 0d 0a 09 05 0a 11 08 11 0c 0e 08 0c 09 06 0f 0a 0c 0d 05 0a 11 0b 11 14 1a 19 22 25 25 29 24 27 2b 27 2a 28 2c 28 31 24 1f 2e 25 2a 25 24 2e 27 24 20 26 2b 23 21 25 19 1c 11 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 12 12 1a 2a 2b 28 2a 2f 38 33 38 42 45 41 3f 3f 3a 3a 3a 34 36 3d 3b 33 31 39 31 3e 3b 32 30 33 30 34 34 37 32 3f 40 41 3b 40 3e 3c 3d 3b 39 3a 2e 24 1d 1e 11 16 0d 17 19 1d 1c 14 15 16 11 08 12 0a 09 12 0c 0c 0b 0c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 0b 08 05 03 02 06 05 03 00 09 05 03 00 06 05 07 06 06 10 09 07 06 09 0b 0b 0b 15 16 13 17 1a 12 11 16 19 1d 1f 12 14 1a 11 0e 17 15 19 15 1a 1d 1b 15 15 1e 10 18 12 09 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 0e 20
 1d 22 20 26 26 22 2e 35 39 37 32 3a 38 36 30 38 3a 33 3c 36 32 39 2d 32 2d 2c 28 28 2e 1e 32 29 29 27 2f 38 2c 2c 27 29 31 2f 28 28 29 22 19 14 0d 05 0b 06 0a 09 06 08 08 01 06 0b 05 0b 06 05 05 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 07 00 06 05 0c 00 06 05 03 09 06 07 09 08 06 06 03 04 06 0b 05 06 06 05 04 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 18 18 22 20 1f 24 25 30 33 34 35 34 39 34 37 3a 2f 2d 2a 2d 2d 2a 2f 25 23 2b 20 16 18 1e 1f 1e 20 23 2d 26 26 21 27 23 25 20 20 24 22 21 1f 14 0e 06 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 18 18 1b 1b 22 1c 22 29 2c 29 2d 24 36 2b 30 28 26 24 26 2b 25 1f 21 20 18 15 14 0d 06 0e 0d 13 12 16 17 19 14 0e 1a 11 13 18 1a 1e 17 11 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 04 0b 13 14 1b 1b 20 1b 26 19 25 24 25 21 24 1a 17 1b 11 11 13 1a 09 0e 05 06 06 03 01 06 09 03 00 0a 05 0d 07 06 12 0f 0d 13 12 0a 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 06 19 13 0c 17 12 18 18 0d 13 0f 0d 0c 0a 07 0b 04 04 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0e 0d 08 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 03 0f 06 05 04 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 05 06 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
