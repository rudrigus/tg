 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 09 06 08 0a 12 10 07 1c 16 1a 19 19 18 22 2a 2d 21 18 1e 1e 1f 1b 2d 33 2f 34 29 1f 20 25 25 1d 25 25 20 1d 1f 1e 0b 14 0a 0a 0e 08 09 0e 0d 18 10 09 0a 03 07 06 05 07 00 06 05 09 0d 06 05 06 03 06 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 06 05 0e 05 0b 09 03 0b 07 0a 10 12 14 0f 15 17 15 17 23 1e 29 24 2d 30 28 29 32 20 2e 34 25 2c 2a 3a 3a 3a 3e 44 3c 3e 44 38 36 39 2d 34 2e 38 2b 2a 2c 26 20 1c 16 19 1a 24 24 33 3b 29 1a 1d 14 07 09 13 14 0f 0b 0d 10 0f 0c 14 06 0b 09 00 06 06 05 0b 06 06 0c 0c 06 05 03 00 06 05 03 02 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 05 03 04 07 0a 0b 07 06 09 10 01 06 0f 0a 08 09 05 14 12 1a 19 15 1f 20 22 24 29 2b 34 2e 3f 4b 44 43 44 3e 44 45 47 45 4a 4f 52 5a 58 56 66 64 64 5d 54 52 51 48 4f 46 42 4a 44 3f 3c 31 27 2c 27 2d 47 49 47 35 34 2b 1c 17 1d 15 1e 18 1b 0f 1a 1a 16 1e 14 12 0a 08 0e 06 09 06 05 07 0d 06 05 03 02 06 05 03 00 06 05 05 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 08 02 06 05 03 0a 06 05 03 09 06 0f 0b 0d 06 05 14 0e 0c 11 05 0f 14 15 17 24 30 25 27 2b 2a 3f 4d 4f 4f 60 5d 67 6d 64 6e 67 6c 65 63 69 6d 74 77 7b 7a 77 7b 82 81 84 85 7b 7a 70 6a 67 69 67 5a 5b 5e 57 51 4f 50 49 4e 55 53 55 4b 4a 50 40 2f 30 2f 36 33 2c 29 27 28 2e 24 1d 1a 1e 16 1c 0e 17 14 0c 17 0f 06 0d 08 09 0c 05 04 00 06 05 03 04 06 06 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 03 00 06 05 03 10 09 05 11 0f 0d 0d 12 08 0d 0d 0d 10 19 14 0d 18 1b 24 3e 49 4a 54 5f 59 5c 65 73 73 73 7c 83 85 85 8e 94 84 85 90 96 96 97 94 a0 a4 9d a8 a2 ac a5 a0 a6 af aa a7 a0 8a 88 7b 68 6b 62 60 68 64 71 6e 77 7a 7a 6f 74 6d 6f 61 5b 5c 56 53 54 4f 4a 45 3f 42 38 40 2e 2e 2b 31 2d 26 1c 1b 19 16 15 1a 0b 11 0c 05 03 06 08 08 03 03 06 05 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0b 05 06 08 06 0b 0c 04 09 0d 09 09 19 15 18 11 10 17 25 1d 27 1e 23 2b 29 3a 5a 6d 7b 7c 7e 7e 7d 86 85 99 ae b9 ba b8 ba a9 b1 9f 9f a8 a8 af b6 c0 be c7 c7 c1 c1 c4 be b1 b4 b5 ba bb b6 ae 94 88 7a 82 82 7a 70 74 7b 82 7c 97 90 95 96 8e 8a 88 88 84 85 86 83 73 76 72 6c 64 5f 5b 4e 5d 54 4b 41 4a 36 35 2b 27 0f 21 1e 16 16 0f 11 11 15 0b 0e 08 0e 06 05 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 06 05 07 0a 09 09 0e 14 0d 0e 17 14 11 1b 1e 29 27 2a 32 30 38 36 3e 40 4c 4e 6d 95 9d 90 9a 8c 99 94 96 a8 b5 c6 c2 bd b8 a4 a1 a1 a0 a6 a3 b2 b3 b9 bb c0 bd c2 bd bb b2 b1 b0 b4 b6 b7 b5 b0 a3 9a 95 95 8e 94 8b 8a 7e 8d 8c 8d 8f 98 94 98 94 a0 a7 a2 ad a9 a1 96 90 8f 83 87 85 7e 71 6d 5f 59 59 55 56 4a 50 4a 4b 40 2b 1c 22 1b 13 16 17 15 0e 0f 14 0e 10 12 0d 05 09 07 06 05 04 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 05 06 06 04 01 0c 08 10 0e 06 17 15 11 0e 1b 23 1f 27 34 3c 4f 5d 5d 64 62 5e 5f 67 6e 71 73 86 9e 9a a1 a0 a3 a5 aa b3 a7 b0 ae ad af ae a6 a6 ab ac b4 b6 be b8 c0 be bd ba b5 b2 a9 a8 a5 a5 ac a6 ad af ab ab ac a9 a0 a8 95 99 9e 90 9b 95 92 99 97 97 94 8f 91 92 9b 9f 9e a0 95 8e 8a 83 7d 76 74 6a 69 63 60 58 5c 56 51 52 55 50 50 52 45 3b 32 28 24 26 20 1c 19 1b 11 12 0c 06 0f 17 09 0d 06 06 06 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 06 0e 09 07 0a 11 12 1a 1b 13 21 27 2a 33 42 4e 5b 79 82 83 86 85 82 8b 8c 94 8b 88 9a 88 94 92 94 90 9f a7 a8 ae a7 b0 ae ab a7 b0 b2 bd bd c7 cb d0 d3 d3 d8 cd ca c1 bb ac ab ab a7 9a 9d 96 91 98 a2 a3 a2 ac aa a1 a4 9b 99 99 97 8e 94 8a 8f 8c 96 91 83 8c 89 88 86 86 82 81 7a 79 71 75 68 6e 5f 58 61 57 55 57 55 54 55 51 52 5c 67 60 4e 3c 2e 36 28 27 2a 21 26 1f 0f 1e 13 0c 07 09 05 0b 04 06 0c 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 04 0e 07 05 12 0b 16 15 23 29 28 2f 34 41 41 5a 69 77 81 8c 85 8f 85 7d 83 86 86 89 8c 94 8d 8f 91 8e 8e 94 92 8f 95 a3 b4 b9 b7 be c5 be cd d5 df e6 dd ee f1 f3 f8 f1 ee e7 da d6 c9 c2 c2 b1 ac a4 9d a3 99 a0 9a 95 9f 98 9a 98 99 93 91 89 80 88 85 82 7d 82 87 7e 86 81 80 82 7f 79 7a 79 72 72 6a 6a 64 61 64 5b 5c 61 62 57 4f 5b 51 56 5a 67 70 5b 5c 55 4b 4d 4a 43 35 3f 2b 2f 29 25 1d 12 1f 15 0e 11 0b 0f 10 0a 10 05 03 03 06 0a 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0b 08 09 0b 11 0e 0d 1b 16 2b 2f 3b 47 4f 59 5a 62 6e 80 89 88 80 7b 81 6e 77 7c 79 77 87 89 88 8c 89 8f 8d 88 8f 8f 93 93 a6 cc ce db db e1 e8 f0 f8 fa ff ff ff ff ff ff ff ff ff fc f0 e1 e2 d6 c4 be bb b0 ac ae a1 9b a0 a1 9c 94 8d 91 87 81 88 84 81 80 7a 6b 77 80 79 76 7c 75 7f 7f 81 7e 7e 7b 71 6e 67 6d 68 65 64 5b 60 65 5b 54 5a 55 5e 56 56 55 55 53 5a 5e 5c 62 51 65 5a 59 4f 46 30 33 2e 25 28 2c 27 2c 2a 1b 17 10 05 0a 08 0d 05 03 01 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 07 08 0a 08 14 1a 18 1f 26 30 32 40 45 52 6b 74 70 62 6f 72 74 79 71 76 79 72 77 77 7a 7d 7d 7c 8c 8b 8d 84 95 98 8b 90 98 96 97 ae d2 ec f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f4 e0 e5 d8 d5 d2 c1 be b4 ae a9 a6 96 93 93 8c 84 8e 84 84 8a 7e 84 77 7a 7c 77 6f 6f 77 7c 7b 82 82 7a 78 74 70 70 6c 6e 6c 6a 6b 67 5b 61 60 63 5e 57 58 4d 4e 53 5a 59 55 57 5c 5e 5f 6d 6f 75 76 6c 5a 50 41 38 39 3c 3d 3a 31 25 17 23 12 11 09 12 0a 0b 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 04 0a 06 0b 0e 0f 19 15 1e 22 30 3b 44 52 5b 5e 6a 72 80 76 6c 6d 6a 71 72 71 75 78 75 71 78 7a 7a 82 85 93 8a 90 94 91 9d 9f 98 97 9d a4 ab b3 da f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ee e6 e0 d0 cf c7 bc af aa 9b 9b 97 90 89 94 8b 8f 87 89 78 81 7f 7d 7c 77 80 7e 84 77 82 7c 78 7a 7b 80 6f 78 77 6f 72 72 69 6f 64 6d 64 63 61 64 66 5f 5d 5d 5c 5d 64 5e 5d 64 63 6f 7a 79 75 6c 5d 60 62 70 5d 4e 49 43 37 33 2d 1b 1c 11 14 10 0b 05 03 07 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 07 05 07 13 09 15 1c 25 32 3e 4b 50 64 68 69 6e 72 73 77 74 70 65 66 70 6b 6b 72 75 80 7a 77 81 80 8b 84 90 8f 8b 98 92 99 9a a5 a3 a7 a6 ad b1 b4 c4 dc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f0 ee d1 d1 c1 ba b5 9e 9c 9c 9e 95 99 97 8a 8f 83 89 8d 7f 83 82 84 84 82 81 85 80 81 89 85 84 7e 7a 83 80 83 7e 72 7e 71 72 71 71 66 6e 72 65 6d 6a 67 64 6a 60 56 59 5c 61 6c 70 6b 66 71 74 77 82 74 6e 6a 5c 55 44 3e 39 27 2b 1c 11 10 13 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 04 06 05 03 0c 09 10 13 19 19 26 38 43 58 64 7b 87 80 80 74 74 7b 7a 75 6f 64 63 64 67 65 64 72 74 7a 7d 78 7b 82 83 88 8d 95 9a 96 9f 9f a4 ac ae ab af c0 b9 c0 c9 db ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f3 df dd d5 c2 c0 a9 a7 a3 9f a3 a3 9e 9b 97 99 8c 8b 8c 8b 83 87 80 88 8d 85 83 87 87 8c 8e 87 8b 97 89 8c 88 82 80 79 7e 83 78 7f 7a 77 75 76 6d 70 69 5c 5b 65 52 5d 58 59 5b 5c 64 6b 6f 74 7a 6d 6d 6f 5f 5d 56 4b 3f 40 34 22 1c 18 13 19 0b 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 04 06 05 03 00 06 05 07 03 06 0b 0a 0f 10 1a 2a 2f 3b 44 54 66 82 7f 86 82 78 78 72 74 6e 6b 70 69 6b 6c 6f 65 6c 74 73 70 7d 7b 89 87 82 90 96 9b a5 a0 a7 b1 b6 b1 b9 ae af bd bb ba ce de f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f1 ec dc d7 b8 bf b9 b5 ba b3 a5 a4 a2 a1 99 90 9d 95 91 92 91 88 8c 91 8c 91 88 90 95 9e 95 98 9a 96 97 87 96 91 84 8c 87 8a 8d 84 84 79 71 75 74 5f 64 5d 65 5d 5c 54 59 5d 61 5e 61 68 69 5f 69 61 5f 63 5c 54 60 59 47 41 34 27 18 17 14 14 0d 0c 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0b 07 11 0b 15 12 1e 2c 2e 3e 50 50 5b 5d 67 76 75 75 63 66 67 67 73 60 6b 62 6a 66 7a 6a 76 71 80 7c 7b 86 82 8d 8f 99 9d 9d a2 a9 a6 b8 ae be b5 bc c9 c2 c7 d3 d1 dc e3 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f6 e6 d5 d8 c9 c7 c0 b9 b3 bd b0 ac a6 a5 9d 9b 9a 94 9a 93 95 8e 9b 92 96 9f a3 9e a8 a3 a1 a4 9a 9d 9e 9c 95 98 8b 8e 84 8d 85 80 83 76 75 6f 6c 61 60 6a 64 5c 57 60 5c 5a 60 59 50 65 61 59 57 56 51 5f 6f 72 64 58 40 2f 2e 30 23 20 14 0f 11 13 0a 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 08 09 00 0e 09 10 1f 19 24 26 30 3e 44 53 60 67 5c 56 56 6b 68 62 6e 6a 68 66 65 68 71 71 72 75 74 6e 74 7b 83 85 8a 89 8e 9c 9d a0 a5 a2 ac ad b4 b2 c2 b9 c4 c6 c0 d0 c8 dd de e7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e4 df d6 cc c7 c2 c5 be b6 ac ac a5 a4 9f 9d 99 a2 9c 9f 9e 9f 99 a5 a3 a6 b0 ae a9 a8 a6 a5 a5 99 9e 9e 9e 93 94 8c 7d 85 77 79 7b 74 6c 6b 63 5e 60 68 67 5e 5a 5b 5d 62 5a 64 62 5f 5d 54 5a 5a 62 77 73 6c 5d 4f 48 43 33 2c 1d 1e 10 10 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05
 03 04 06 05 07 0e 11 19 21 26 2e 3d 3e 4b 4e 5a 5f 5c 61 5a 60 63 64 59 5f 65 6c 74 6c 70 73 72 79 7c 85 7c 79 7d 86 87 8e 99 9f a5 aa ab ad b1 b3 b2 ba c4 c4 cb ce cc d4 d2 da db de e9 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f1 e5 dd d3 d2 c6 c3 c1 b6 bb a9 b2 a4 ac aa a0 a4 a1 a6 ad a9 aa ac b5 b9 b4 b3 b1 a6 a6 a6 a4 9c a5 9d 94 9b 84 8e 86 87 82 86 71 72 6e 6e 6a 69 63 65 60 65 62 5f 60 5f 62 5c 57 57 5a 54 52 60 64 64 67 66 60 58 54 48 3b 33 2d 22 1e 08 0d 0d 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 0c 0b 08 10 0d 1d 20 2a 2e 38 43 4d 52 57 5d 5f 61 64 65 65 67 64 68 67 6d 70 76 72 74 77 81 7e 81 82 87 8b 8c 92 92 8d 9f 9d b4 bf bd c4 c6 c4 c3 c7 cb d6 cb d5 d9 db e6 de df ea ed f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f2 ea e7 d5 d5 cb c6 bb bd c0 b5 b3 b0 aa a8 a6 ae b3 b0 b1 b6 bb b7 bb c1 b8 b6 ae ab ad ac a8 a2 a5 94 99 90 8b 8a 86 84 7c 7f 79 7a 6d 69 71 6e 66 6c 68 66 62 68 59 60 69 61 63 5a 5a 57 55 53 55 4d 5d 58 5b 68 65 4e 48 3b 32 2f 1e 19 0f 09 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 0e 0f 16 16 23 22 2c 36 47 56 60 54 52 54 60 5a 62 59 5d 64 61 67 68 6d 70 74 76 7f 82 80 85 84 84 89 91 97 a0 9d 9e a4 a8 b9 bf c5 d0 d6 dd da da db da d4 e4 e1 e4 e9 ea e7 f5 f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 eb eb de d6 d7 ca c9 c5 c4 c5 ba b8 b4 b5 b4 ab b5 af b5 b9 b5 bd b7 c2 b5 b5 b2 b6 b4 a5 ab aa a8 a2 9f 92 91 8c 8f 88 84 7c 75 81 73 73 74 6d 68 6a 66 65 61 60 62 5b 60 5c 57 58 5a 54 4e 4e 53 56 4c 46 51 55 59 60 4e 4d 3a 3a 31 21 1b 19 0c 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 09 06 09 0c 0f
 12 1c 22 21 24 37 3c 4c 57 64 61 59 58 57 56 5e 61 5e 68 6f 70 73 75 78 79 7f 79 83 85 84 86 96 9a 9f a0 ac a5 ab ab ba c2 c7 ce d7 d8 e6 e6 e5 ea e2 e8 e5 eb ef f6 f3 f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f3 ea e4 d8 d8 d3 cc d3 cc c5 bb b9 b5 be bc bb bc bd c5 c6 c5 bf c1 bf ba ba b3 b5 b1 a8 a8 9f a2 9d 95 98 90 8d 8c 8a 88 7f 7f 78 73 72 72 66 60 63 65 55 61 60 5b 5c 60 5d 5d 56 5b 4f 54 4d 50 52 4e 49 4b 4c 4d 55 50 4a 49 41 34 22 1d 17 0e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 04 06 06 0b 0a 13 17 17 1e 23 2d 35 48 5a 6a 65 63 58 50 53 55 5d 6b 66 65 6a 6b 71 7f 80 81 8a 8f 90 8c 93 97 93 9c a2 a4 b0 b4 ae b6 b7 c9 d2 d3 e7 e3 ed ef f9 eb f9 f8 f8 fa f1 f4 f0 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ef ec e3 e6 df db c9 d3 d1 c9 c5 c2 ce c8 c3 ca c4 c4 c8 cb ce c5 c4 c7 bb bd bf af b3 ab ae aa a2 96 93 96 8f 91 90 8f 7e 7c 7c 80 78 74 6f 71 6c 66 60 64 5b 5f 5d 5a 5b 50 5b 5a 57 5a 5e 54 4c 50 45 53 4a 49 49 52 49 43 46 3b 35 22 26 20 1e 0c 0c 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 12 11 14 1f 11 21 23 24 41 52 60 67 61 5a 5c 53 4e 59 58 66 69 66 70 6e 7a 72 84 88 89 90 8f 8b 95 93 9a a4 9f ad af b8 ba bc c0 c9 d0 ce dd e9 eb f4 f7 f9 fe fb fd ff ff f8 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f9 ed ee e5 e2 dd db d6 d7 d0 d0 cf ca cd d5 d6 ce ca ce d0 cc ca c9 ba b9 b8 c4 bf b7 b9 a2 ab a5 9c 90 9b 8a 94 8a 8a 87 7f 82 71 75 6e 71 6e 6b 70 60 61 61 5f 60 5f 62 59 60 5e 56 62 5d 5a 51 4b 4e 4d 51 4e 55 43 4f 49 44 3d 36 3b 2d 29 18 0b 03 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 03 01 06 0a 0c 0e 0c 15 1f 1f 15 25
 28 32 47 60 69 63 60 54 50 5a 54 5a 5b 5e 65 64 66 6f 73 83 89 8b 87 91 90 94 97 99 a1 a5 9f ad b1 b3 b5 c3 ca c9 d7 d9 e4 ec ee f6 f3 fe ff ff ff fa ff ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc f3 f3 f0 de e2 e2 d8 d4 da d2 d1 d9 d4 d7 ce cb d5 d2 d3 d1 c8 c9 c1 bb c3 c2 c1 b7 af b0 ac a6 a3 a2 9f 97 9b 94 80 88 80 7c 82 78 76 74 68 69 66 65 6a 63 5b 61 5e 65 64 61 59 57 60 60 5b 4f 52 52 4b 57 4a 4e 50 51 4b 4a 4b 46 3d 38 39 2d 1e 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 03 0b 05 0f 12 13 1f 2a 1a 27 2e 36 50 6e 81 83 66 54 5d 58 60 61 5b 64 6a 66 6d 79 79 82 89 85 93 9c 9c 9e 9e 9e a7 ad ab b4 b5 bb bb c1 d3 d3 d2 d1 e2 eb f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc fa ff ee f0 e8 e6 e0 dd e2 db d8 d9 dd e1 de e0 dd d1 d0 d4 d2 c6 ce cf c6 ca c4 b7 b9 ae a9 a7 a5 a2 a0 81 97 8d 8f 8a 85 85 82 80 7e 70 69 73 74 6b 6b 6f 63 6d 67 68 6d 6d 61 62 61 5b 59 4a 4d 53 5b 58 58 5c 58 52 55 5a 4e 4d 53 4f 44 3c 24 14 0c 05 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 05 07 08 0d 14 16 18 18 26 1d 27 33 42 60 78 87 89 72 5c 59 5a 5b 5f 67 64 6d 68 6f 74 7c 80 89 9a 92 9a a1 9e b2 a3 ad ac af b9 b7 bf c2 cf d0 dc e1 df eb f1 f5 f2 fc ff ff ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 f4 ef ef ea e5 df d9 df e2 df e4 e0 de da dc d8 d6 d0 cb cd d0 d0 cb c4 be be ba ae a6 b1 a3 a0 a9 97 9c 94 8e 87 89 84 89 8a 7e 7f 7b 71 71 7a 71 6d 70 6b 70 69 6d 64 62 62 5d 56 57 57 55 57 58 54 5d 57 5a 59 53 56 54 4f 4d 50 49 3c 27 0f 12 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 08 06 05 08 04 06 0e 11 0a 0e 07 12 1b 18 24 2d 32 4e 69
 85 86 80 78 60 57 5a 5d 67 6c 64 76 68 73 7a 82 83 85 98 9d a0 9e ad af ab a8 b2 b4 bd bc c1 c6 cc cf d8 de df e7 e8 f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff f7 f3 f4 ee eb e2 e4 e5 eb ea e7 ea e4 e0 e0 dd e6 de de db d4 d2 d1 d2 c7 c0 be ba bb b0 b0 b2 a3 ab a4 a0 a1 99 93 8b 92 88 89 82 7f 7a 7a 7b 84 7a 79 72 6b 69 74 6a 68 66 66 65 5e 50 58 55 5d 5e 5f 5e 5c 5c 5e 59 5c 59 56 5d 54 5a 48 40 30 10 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 0e 06 05 0e 0e 09 0a 12 12 13 17 20 23 29 36 40 57 80 89 88 81 6d 59 56 5d 5b 63 66 70 6e 75 75 7a 85 89 96 98 9c ae a7 ae ad b3 b4 b0 b4 bf c3 d0 d0 c9 d7 dc e1 eb e8 ed fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb f4 f1 eb e5 e9 eb ea e9 ee ed eb e8 e4 e2 e4 e0 e0 da da d4 d3 d6 cd cc cc c9 be ba b3 b7 b4 ac a4 a7 a7 a3 9f 9d 96 98 94 8c 88 8c 8a 88 7d 88 80 7a 84 76 74 7a 71 73 72 68 68 67 5a 62 5f 5b 58 64 63 5b 65 62 65 60 61 61 64 60 62 55 41 25 17 0c 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 12 0d 0c 0b 0a 0f 1b 0a 11 1d 14 22 2a 31 3a 4a 64 74 8b 92 7f 6b 5a 5f 5e 65 5e 75 6a 78 7d 82 88 8a 95 94 9d a0 ae ae b8 bc c0 b4 c5 be bf ce cc ce d8 e2 df df ea ed f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f2 f7 ea f0 f2 eb e9 f1 f4 ed eb ee ea ef df ea e4 e6 e7 e4 e1 e1 db d4 cf ce cc c1 c4 c2 bc bb b7 b7 b4 b9 a7 a6 a0 a5 9a 9c 99 93 8e 88 88 95 89 80 7f 7d 7e 74 7f 81 7a 72 75 68 68 67 5d 63 65 64 60 64 66 6b 67 6e 65 64 5b 65 6b 70 65 4d 30 15 13 0c 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 04 10 06 0e 19 1c 17 17 20 23 1d 2a 2f 39 48 6e 83 8c 8d 7a
 69 59 59 57 5e 65 72 73 71 81 88 89 97 9e 9f a6 a4 b6 b1 ba c6 ba c7 c3 c7 c9 c8 cb d4 d5 dd e5 e8 eb f0 f9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fb ef ef f0 ec f0 ec ef e6 ea f0 ec f1 f1 ef f1 ee ef ed e7 e8 e5 df e4 d6 de de d8 d8 c7 c5 c7 c6 c6 c3 b3 bd b8 b1 af b4 a7 a8 9f 97 99 92 9a 90 96 8d 8b 85 82 83 80 7f 84 81 78 73 70 64 66 5f 6c 67 65 72 6e 69 6d 69 6b 65 65 6c 64 6a 81 72 55 31 23 15 0d 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 09 0b 09 0f 10 1a 15 12 18 26 2d 3a 4b 5f 7c 85 7c 8a 74 62 54 52 5f 68 6b 6c 77 7f 84 8f 9b 99 aa a1 ac b0 c2 c5 cb c4 ce ce d4 d2 d6 d5 d0 e0 db e0 e8 f1 f9 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff f9 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f6 f8 ea e9 ee ed f2 f2 ec f4 f1 f4 f8 eb f0 f1 f0 f4 ef f5 ed e0 ec ed e4 e7 e0 e2 df df d8 d0 ce d2 c2 cb c6 c0 bf b3 b6 b6 b5 ad a1 a4 a1 a0 aa 9d 96 9a 8c 8f 97 8f 8f 86 87 89 7c 70 6d 65 6d 65 6d 6b 6a 72 74 6c 75 67 71 6f 6e 70 6d 70 7c 76 4f 39 20 19 14 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 0c 06 0c 06 0a 07 15 19 1b 22 25 1b 25 2b 3d 56 7f 8b 94 8e 8a 74 60 54 5e 64 64 6c 74 7d 8e 8a 95 a1 a9 ae b7 c5 c4 cd cb ce cc d0 dc dc df df da e0 e2 e5 e4 ee f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fe fd ff ff ff ff ff fd ff ff fb ff fe fb fc f8 fd f8 fb fd fb fe fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f4 ea ed ec f5 f2 f0 f2 f0 f3 f6 f6 f0 f5 f8 f7 f9 f2 f5 e9 ef f0 ed ed ea ee e5 e4 e6 e6 d9 d4 ce d2 d7 d6 cb c8 c6 bf bc b7 c0 b2 ad a9 b0 a8 a1 a5 a4 9a 9a 9b 99 91 91 91 83 85 82 79 73 6e 6c 71 76 6c 7b 73 76 73 6f 72 6e 75 6b 6f 6f 81 8c 73 54 38 1f 1f 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0c 08 0a 11 11 17 12 1c 1b 22 2d 2f 33 3c 5f 7d 8f 9a 9b 8f 73 5d 5b 5e
 64 66 6e 78 80 84 91 97 9f ae b1 c4 ca c9 de d9 d4 dd e4 de e2 e3 e9 ed eb e2 f1 e8 f4 f7 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f7 ff f9 ff ff ff fd fb ff fa f6 f6 fb f7 f8 f4 f8 f2 fa ee ea f1 f6 ee f4 e7 f4 f3 f2 f6 f8 f3 f9 fd ff fd fe fa ff ff ff f6 f8 ed e4 eb ed ec f3 ee ed eb f1 f0 f2 f8 ef f0 f6 f9 f6 f5 f1 ee f1 f2 f3 ed eb f4 ea e0 e3 e6 e3 e1 e1 d6 da d6 cd c8 cb c8 c0 c6 be b9 bd b2 b0 aa aa a3 ac a7 a2 a0 a2 95 97 98 8b 8d 84 81 75 77 76 6d 75 74 74 7a 78 76 7b 71 72 73 6d 79 84 91 8f 6e 50 41 30 1f 0e 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 08 0d 16 11 0e 14 13 1e 16 21 1f 35 34 4b 5e 5b 6c 83 90 96 95 83 65 58 5c 61 65 6a 74 79 88 93 a0 a7 ad bd be d1 d8 dc e0 e4 ef ef ea f3 ee f2 f5 eb f1 f1 f1 f9 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff fe fd fd fc ff ff ff ff ff ff f6 fb fb fa f7 f5 f3 f8 f3 ed f0 f2 ee ee ec ef e8 e8 e9 e7 e8 ec ed f0 f4 f9 ee f8 fa fd f7 fc fc f5 ee e9 e6 e4 eb e7 ea f3 f7 ef f0 f8 f3 f6 fa f9 f5 f2 f6 f3 f3 ef ed f3 fc f0 ef ee e8 e2 e8 ef f4 ee e4 e2 dc cb ce d0 cc c3 c7 c1 c1 bd b8 b3 b3 af b1 b4 af ab ad a5 9c 99 92 92 8c 88 81 79 7b 74 6e 85 7e 81 76 77 74 7e 78 78 72 79 76 82 9b 96 7b 66 4e 34 23 14 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 07 05 12 15 1d 19 16 1e 1b 1c 23 31 3a 55 67 80 8a 86 83 8b 91 9c 92 6f 5b 61 59 66 73 77 7a 85 96 9b aa ba bd cc d1 d7 e6 e6 f2 fa f8 f8 fe ff fa f9 ff f6 fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fc ff ff ff fe f7 ff fd f7 fd fa fe ff ef f9 ef f0 ec e9 f1 ea e9 e8 ea e0 dd ea eb e5 e1 dc e7 eb ee ee f5 f2 ee f6 fa ed eb e8 e8 e9 f2 f1 ed f4 ec ec f2 f7 ff f5 f7 f7 f3 f3 f5 f9 f9 f8 f4 f1 fd f0 ee ef f6 fd ff ff ff fb ef e4 da d8 d3 d0 c5 c9 c8 c3 c2 c8 c7 c4 bf ba b8 b5 b7 b0 b0 a5 9c 9f 92 95 8b 89 89 86 7f 87 7f 86 7a 80 81 79 74 75 76 72 75 73 7d 92 a2 9f 8b 6a 5e 44 35 23 11 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 0f 11 20 1f 15 18 1e 22 21 31 44 5e 78 93 95 a2 9a 87 84 84 7a 74 5d 5e 60 65 65
 75 73 82 8e 97 a0 b6 c4 cc d9 df e6 e7 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff ff ff ff ff ff fd f8 f7 fe f9 f6 f8 f4 f3 e9 f0 e6 e8 e3 eb e4 df de e1 de e1 e0 e6 e4 e9 e8 e4 e4 ed ef e9 e5 ee e1 e0 ef e3 e7 f0 f5 f3 f1 f3 f6 f9 fb f4 f5 f2 f2 f4 f6 f1 f5 f4 ef f5 f0 f1 f6 fd ff ff ff ff ff f8 ea db da d5 d6 d5 cd d1 ce c6 cb c4 c7 c4 cb bc be bb bb b0 af a5 a2 a3 9c 94 90 89 88 89 7c 86 7f 83 7b 7e 7e 80 72 7a 76 75 73 75 75 83 9a aa a8 8c 63 45 3f 25 21 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 1d 18 23 23 1e 24 20 35 3b 52 70 8c 96 9b a8 a4 a0 88 7f 68 65 65 61 64 6c 6f 73 78 81 8f 91 a0 a7 b7 c4 d7 e3 e4 ef ef ef fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff ff f9 ff f6 fc fe ff fe ff ff fc fa ec ef ec ef ec e9 e2 e4 e1 e0 e4 de dc da da df de e0 e6 e4 e6 e5 e7 e5 e2 e0 e8 e4 ef eb e3 e9 e6 f3 f0 ee fa fb f6 f7 fa f4 f1 f4 f2 f3 f8 ed f5 ef fb ff ff ff ff ff ff ed e0 df e7 d4 d6 da cf d7 d7 d2 ce ca c7 c9 c9 c5 be c2 b5 b2 b5 a9 9d a0 8d 93 92 8f 8f 84 85 7f 78 75 7e 7b 72 7d 78 7d 74 75 72 6a 68 74 89 a6 ab 94 6f 53 3d 29 1a 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0b 0b 0b 1e 26 22 25 34 39 37 3d 4f 6e 86 92 9c a3 a8 aa a4 9f 85 76 6b 65 5f 67 68 66 77 81 80 89 91 95 a5 b6 c4 cf d9 e5 e7 ee f8 fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fa fa f1 eb f0 ec e6 eb eb e3 e1 d8 e0 dc e2 dc db e0 d9 e6 d9 e2 ea e4 e0 e7 e8 e6 e9 e5 ec e3 ed eb f1 f4 ef fb fa f0 f9 f9 fb f6 f7 f0 f1 f4 ee f4 ff ff ff ff ff ff ff f3 e4 e0 e1 dc e2 d8 d0 db df db c9 cc ce d1 c6 bc c0 b9 c1 af a9 a9 a8 a0 9e 9a 96 94 8e 85 84 7e 82 83 7b 7b 7c 7a 7d 77 75 73 6f 6d 68 72 6d 84 9f a9 90 78 54 44 2f 21 18 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 07 11 14 20 22 35 42 4e 5b 55 5e 71 8c 98 a6 9a a8 b8 b0 91 83 6a 5e 6e 60 69 7b 74 79 7c 7c
 8c 8f 95 99 ad b6 c7 d7 df e6 ec f3 f9 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f5 f0 ea ed e9 e4 e4 e0 e2 e4 e0 e3 dd e0 dd e0 d7 e1 df e0 dd e5 e3 ed eb e9 ef f6 ee ee f5 f1 f6 f7 f1 f4 f9 f5 f3 f5 f0 f5 f3 f6 f4 fc ff ff ff ff ff f6 e5 e7 e5 e9 eb dc e5 e3 dc dd de d8 ce ca c4 c9 c3 c1 b6 be b3 aa a8 a5 99 9b 9e 97 91 8d 87 83 8a 7e 7e 78 77 78 79 7c 75 7a 6e 67 72 70 74 75 77 90 b5 a6 89 68 4b 3f 27 14 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 0a 0a 1d 22 28 32 45 5e 61 72 7d 85 8e 8e 98 a5 b1 b0 a3 8b 79 6b 69 69 68 78 76 75 7c 86 82 86 8b 9a 9e a6 b7 b0 c4 d3 dc e0 ee ee f7 fa f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f0 ec ee e4 e4 e1 df d8 e1 db dd dd dd df e0 e4 e2 d9 e0 e4 e1 e7 e5 eb f0 ea f1 f2 ee ed f1 f5 ed f3 eb f0 ec fa f4 f6 ee f5 fc fe ff ff ff f3 f1 ee ed e2 e9 e4 e1 e1 e0 d7 dc d7 cd ce c6 c5 c5 bf bc b7 aa ac a7 9e 9e 99 96 90 90 90 8d 80 7c 80 81 81 77 75 7c 7a 6e 73 7c 6c 6e 71 71 6b 72 72 85 af a6 92 70 52 44 37 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 0a 12 1d 29 3a 50 51 5d 61 77 89 a3 a5 97 88 99 90 9c 91 8b 78 73 6d 71 79 7c 79 7c 8a 83 86 8d 86 95 a3 a5 a5 b0 c1 c4 d5 e5 dd e9 eb f3 f8 f9 f3 f8 fa ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f8 f1 e3 e7 e1 e9 e2 da df de dd dc c5 dc e0 e1 e9 ea e1 ec e4 e2 e1 e8 e9 ee e9 ee f6 ee f5 ee f3 ee ec ec f1 f7 f3 f5 f2 fa fc f7 f0 eb f2 e9 e9 e6 e3 ec e6 e5 db d7 d6 da d6 d1 c2 bd b9 bf b4 b5 b1 a5 a2 a3 a1 99 98 92 8e 84 85 7f 7c 77 7c 74 7f 79 7f 74 7e 6c 74 75 76 77 72 72 75 78 8b a9 b1 98 75 5b 45 30 25 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 0d 0b 1d 2b 39 4b 5d 65 75 74 88 9e b5 bc 8f 84 78 7f 76 7f 7a 76 6e 70 75 73 7d 80 85 91 8d 84 93 99
 9a a0 a4 a8 b3 b9 c7 c8 d7 e0 e1 eb eb fa e7 f3 fa f9 fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 e6 e4 e4 dc de de dd dc e7 de df da e1 df de e3 e8 ea ea e7 e5 f0 eb f2 f2 ee f0 f2 ed eb f5 f7 eb f1 ec f3 f4 f6 f1 f2 ef f4 ea ed f0 e7 e9 e9 e3 df da dd d7 d0 d5 cc c3 c3 c1 bb b2 af ad a8 a6 9d 9b 96 93 8d 8a 83 7f 7d 74 7b 78 7b 78 77 70 79 74 7b 72 78 6c 7a 70 75 6e 73 87 b2 ae 9a 76 61 41 37 23 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 0e 1b 2e 3c 4b 56 58 75 7e 8f a0 a9 bb b1 91 7c 7a 73 79 81 7b 75 75 72 79 75 7d 7a 83 92 8a 91 95 96 9f a4 a4 ab bb b3 c8 c8 d1 db e2 de ea ed f4 ee f5 f6 ef f3 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e9 ea e3 df e6 dc e4 de d8 e0 de e3 e2 da e3 ed ed e9 e9 ed ef e9 ee e6 f0 f2 f3 f6 f2 f5 f2 ef f3 f5 fb f1 f4 f3 f4 f2 f3 e7 e4 e0 e8 eb ec db e3 d5 d4 cb d7 c5 c7 c0 b6 b9 aa a3 a5 a6 a4 9e a7 93 92 8b 85 86 84 7e 7c 75 74 72 7a 75 79 70 75 7c 76 75 71 75 6f 66 69 6e 6e 80 af b1 97 82 63 4b 31 23 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 13 25 37 49 63 69 77 81 97 a1 a6 ae b6 9c 83 83 73 7c 7c 7d 7b 82 7e 7e 84 84 88 84 85 95 95 94 a0 9a a3 aa aa b0 ad b8 c4 cd d0 e0 dc e2 e5 e7 ed ee f0 ed f4 f5 f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ea e5 e4 de e4 e3 e2 e0 ec e5 e4 de e6 e7 e8 eb ea d8 ea e5 ee f5 eb f5 f8 f4 f6 f0 f0 f9 fa f6 f2 f6 f0 f2 ef f8 f1 e6 f5 eb e4 eb e7 e8 db df d4 ce ca cb c0 bd b9 b8 b9 af a9 a4 a7 9c 99 94 94 8b 8c 82 79 7e 7b 74 7e 76 7c 76 7b 7b 77 7a 82 76 74 74 70 69 6e 64 74 79 8a ae b3 a0 7b 6c 56 3d 2a 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 14 25 33 40 57 6d 75 8c 99 a6 a4 a4 ab a7 94 7d 7b 75 7e 80 88 81 87 7e 84 8d 8b 8d 91 91 9b 9f a3 a3 a8
 aa a6 a9 b4 b9 bf cb cc cd d1 d0 e1 e5 e0 ee e5 ec ed f1 f1 f9 fc f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 ed e5 e4 e8 e3 db e2 e2 e5 ea e5 e1 e4 e4 e7 ed e4 f0 ec eb ef f7 ef fa ee f0 fb f4 f3 f6 f4 fa fc fa f4 ef f1 f2 eb f0 ea e9 e7 ee dd da da cf cf cc c8 c5 ae b6 b9 ae b0 ad a4 a1 9b 91 8c 8b 85 7d 84 79 7f 77 71 76 84 77 7d 7d 7d 80 7e 6d 7b 71 70 6f 69 6b 65 72 89 b4 ba a2 88 6e 55 46 2a 11 09 03 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0b 13 2a 36 47 5f 78 8b 9a ae b1 9c 96 96 94 80 74 78 77 73 79 7a 84 81 84 87 95 8f 90 94 9a 9f 9a a8 a3 a5 b0 b2 b1 bb b9 bc c4 c8 c8 d0 d4 d8 d8 dc dd e5 ee e7 ec ec f1 f7 f2 f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 ef ec e3 e1 e3 e5 df e1 e3 e3 e6 e8 eb eb ec ea ee ef f0 e6 f6 f7 f1 f7 f4 f5 f3 f5 fc f7 fe f7 f8 f7 f0 f8 ee e6 e8 e9 e4 de e1 dc da d8 d0 cc cd c3 c3 b0 b1 a7 a5 af aa a5 9d 91 91 83 78 84 7b 80 77 7a 7e 7f 76 78 83 7e 75 7a 73 76 79 6e 6a 6a 6b 65 6b 64 6b 8b b6 b0 9e 84 66 53 3d 29 1a 09 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 10 1f 25 42 53 66 84 96 a5 b8 a9 84 84 7f 87 7e 73 6f 73 73 77 80 82 7e 8a 92 93 94 88 9d 9e a6 a5 a3 aa af b2 b1 b6 bc be b9 ca c5 c6 cf d3 d1 d9 dc de e3 e8 e4 eb e7 ee f1 f5 f6 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fd e6 ec e8 e4 e4 e6 e7 e4 eb e8 e6 ed f0 ed ef ef ef ec ef f5 f5 f8 fd f8 f5 f3 f1 f4 ef f3 f6 f5 f3 ee ef ed f1 e8 e5 e2 e4 e4 da d5 dc c0 c9 c6 c2 bf b9 af b0 b1 b0 a2 a4 9c 8d 8b 84 7b 81 84 83 7b 7b 7f 83 79 7c 7a 77 80 78 7c 74 7a 74 6a 6e 67 68 69 65 68 87 a8 ba a8 8e 71 5b 3a 2d 15 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 09 14 13 25 28 4b 60 73 90 a0 b8 b0 8b 81 77 78 7a 79 6e 79 6e 7d 72 7a 7f 7a 82 8e 8d 97 93 9e 95 b0 b4 af b8 bb
 ad b6 c0 bd c3 c1 c7 bb c7 d9 d4 d2 db d7 de de e6 ec e8 f0 e6 ec fe fc f6 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 eb ef e8 e8 e3 e2 e4 e7 e5 f0 e6 ed f4 ed ee eb f7 f1 f2 f4 ec f4 f7 ff f1 fd fd f4 fb f9 f8 f6 f5 ec e9 e5 ea e8 e1 dc df da cd d0 ce ca c4 bf bc b9 b6 af b3 ae a8 a3 92 90 93 8a 84 86 85 7c 87 7d 80 79 7b 7e 80 80 7f 7c 76 7a 74 6e 6e 69 64 66 66 68 68 81 a8 b2 a6 8d 6a 53 3e 23 19 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 11 0d 1f 29 39 4c 5c 77 94 b4 bc a5 85 77 76 76 76 74 73 77 7a 71 78 75 79 84 7c 85 82 8f 8e 98 96 9c 9b a4 b0 ae bc bc c0 c3 c4 c5 c4 c6 ce c8 cb d5 d7 d8 db da e0 df e9 e7 ee f8 f0 f4 fd fa fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff fe fc fc f3 fe fa fc f9 fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 eb e2 e6 e7 eb e9 ed ed eb ec f2 ee fa f5 f1 f0 f3 f7 ee f7 f6 f8 f7 fe f8 f6 fa f4 f2 f2 f6 ed eb eb eb e1 df d4 e5 d8 d0 ce c7 c6 c7 bc be b6 b5 b1 ab aa ad a2 9a 95 92 8f 83 83 85 87 83 80 86 7f 7c 7b 7e 82 80 7e 7d 73 78 6f 75 6e 6a 63 63 5e 68 7c a0 ac a3 8b 6f 4f 30 18 0d 0d 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 09 15 1e 27 3e 4a 5d 7c 91 b9 b3 9c 85 7a 75 77 7e 74 73 7e 76 73 72 76 77 76 7c 78 87 8f 92 93 94 a0 9e a2 ac ab b5 b4 c0 bb c1 cc cb c7 c6 df d1 d5 d9 d3 d2 df e1 df e8 e5 ea ef f6 ef f7 f5 f3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff fd f5 f5 f4 f0 f3 fb f2 fe f9 fc ff f9 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ec ed e5 e9 ea e5 e1 ee ed ed ee ef ef f5 f2 f1 f2 f0 f3 f8 f3 f5 f5 f2 f6 ea f1 f8 f2 f0 e9 e9 e8 df e0 e7 e0 e4 e1 d8 d1 cc c6 ca ca bd b8 b9 b1 b7 a5 a5 a6 a2 a0 93 9a 94 80 8b 81 8d 8a 7c 80 86 7e 7d 84 84 85 83 7c 78 76 6f 66 6b 65 67 6b 66 64 75 9a a1 a4 83 67 46 24 1f 12 0b 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 09 1d 27 30 44 4d 69 82 a0 b5 b4 96 82 83 7d 80 7d 7e 72 82 7f 7e 73 80 7f 7b 7c 7b 88 8f 8e 99 9c 9c a1 a4 a1 a7
 b7 af b7 bf bb c2 c1 c1 cd cb d2 d3 d5 df de db e5 db dd eb ec ee f4 f7 f4 fe fd ff ff ff ff ff ff ff ff ff e4 fd ff f9 ff fa f5 fa fc f1 f8 f9 fa f3 f4 f3 f4 f8 ff fc fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ec ec eb ee e6 ea ee ec eb eb ef f1 e7 ea f0 fc f9 f1 f8 e9 ee f9 f8 f3 f2 fb f3 ec ef e9 ed e4 e4 e1 e1 e5 da da d9 cf cd d1 c8 c4 c3 c8 c2 b3 ba ae af ae af a3 9b 92 96 8e 92 90 86 87 83 8d 8f 8d 97 85 89 84 87 7f 81 7a 6f 71 70 6f 65 6b 61 6b 7a 8a 9d 97 84 5d 40 2b 18 09 08 0a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 0c 12 2b 3c 4b 59 76 8a 97 b9 b9 9e 81 83 83 7f 80 7e 7f 86 85 80 82 7e 80 79 7d 81 83 8e 92 90 92 9e a3 a6 a9 b1 b5 b1 b5 bb c3 bb c0 c7 cf d2 d0 d2 d1 d5 d5 dd e0 e0 e4 ee ec f5 ee ef f9 fc ff ff fd ff ff fd ff fe fe ff fd ff fa f1 f5 f0 f5 f4 f9 f6 ee f4 ed ef f9 ef fb f2 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f3 e7 e5 e9 ea e8 f1 e7 f0 e8 eb f6 e9 fc ed f5 f4 f2 ef ee f6 f6 fa f9 f2 ee ee ed ef eb e9 e9 eb e0 e3 e0 d8 dc d6 d3 ce d0 c6 ca c5 c4 c2 c1 b2 b4 b0 ac a8 9e 9a 9a 93 90 8e 90 8c 8c 8d 8e 8e 8c 8e 82 90 83 89 82 87 7f 75 6e 71 67 62 6b 66 69 6a 83 99 91 7e 56 3d 22 18 0a 0b 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 11 26 35 4b 4f 5c 69 80 96 ab ba a5 84 79 74 7d 82 80 7f 8a 84 83 86 84 85 7f 7d 82 87 89 92 91 93 98 99 a6 ad ae b7 b1 b3 b8 bc bb c6 ca ca cb c8 d2 d3 d8 db df e1 e4 e9 e8 eb f2 f5 f6 fb fe ff fa ff ff ff fc ff fc f6 ff f5 ef f5 f3 f5 e9 f5 ee f5 ee ed ed f3 ee f7 f0 f0 f5 fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 ee ef e0 e9 df e9 ea ec eb ee ea ea f3 eb ef f1 f1 f2 f2 f1 f1 ef e8 ec eb f5 ee eb e3 e5 e0 e5 ea db e1 dc d5 d1 d5 cf cc c9 c8 c9 b9 bf be b4 b3 b2 ad ae a8 9c 99 92 97 93 93 92 89 96 92 8b 8b 8a 8c 91 89 8c 81 7a 85 75 7a 6f 72 62 63 61 62 6b 7f 8b 89 6c 4b 34 15 0c 0f 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 05 06 13 23 3e 4d 63 6d 75 89 9a ab bf a2 83 76 7b 79 7e 7a 8a 87 88 84 8a 8b 88 80 89 87 8d 8c 89 92 98 94 a0 a4 af a8
 b1 b8 bb bb c2 c8 c4 c9 d0 d5 d3 da dc df e2 e0 e3 df e9 ee e8 ee ed f5 f6 f8 fb ff ff ff ff fc ff ff f5 f4 ea eb f3 f3 ee ed ec f0 f2 f1 f4 f5 f2 ea f6 ef f1 f5 ff fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f4 ea eb e7 e3 e8 ea e6 e9 e8 eb ea e8 ef ee f0 f6 f4 f8 f3 f5 ec f3 ee ed f1 ee ed e8 e5 e5 e1 de e5 e1 e1 d9 dc d5 d7 d1 ce ca c7 c7 c6 be be b8 b2 ad aa a7 a4 9a 9d 9e 8f 96 92 97 8a 93 96 8c 90 8e 91 8c 85 8a 7a 80 7e 79 72 76 6a 60 68 64 68 6a 77 84 88 6d 52 36 28 19 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 07 10 13 1f 29 3d 4b 6c 77 7a 7f 9c a3 b3 a4 77 6e 72 76 77 7a 81 85 87 8c 82 86 86 90 89 8e 8c 95 96 95 9b 9f a4 a5 ad b0 b3 bc ba be c5 c5 c9 cb cf d5 d1 d0 dc e0 e3 e0 dc e6 ee ee f4 f1 f5 f6 ff f8 ff ff fb fd f8 ff ff f9 f7 f3 f3 f2 f0 e8 ec e5 eb f3 ef f5 ea f5 ed ef f1 f2 fa f4 ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f4 eb e3 e8 de e4 e7 e6 e1 e4 e2 e8 ef eb eb ec ed ea ee f6 e6 f0 f0 e8 ef ef e2 e2 e3 e5 e0 e8 df de d5 d9 e2 dd d6 cd d2 d4 cd cd c5 cb c9 c0 bf b8 ae ae ad a7 a3 a2 95 92 98 92 95 99 94 95 8c 8e 94 99 96 8e 87 82 8c 80 76 77 6f 6d 6a 6e 64 68 6d 7b 8b 85 69 44 2c 24 1a 0d 0b 07 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0e 1e 37 39 59 6d 87 8a 85 83 8b 98 89 6f 64 6e 6f 76 7d 79 7e 87 88 88 92 8d 83 92 90 8f 95 8f 9d 99 a0 a6 9f ad ae bb b1 c3 c0 c7 c4 c6 c4 d3 d2 d4 d9 d9 df e4 e7 e6 e7 f2 ea f2 f7 f6 f4 f4 f6 ff ff fb ff f9 fc f3 f0 f3 f3 f7 f1 ef e8 ec ea f4 f2 f3 ed f6 ee ed e8 f1 e9 f9 f8 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 eb e1 e9 e5 dd df de de e4 e1 e5 e5 e8 ed eb e8 ef ed ed e5 e8 ed e9 e6 e6 ea ea e5 e5 e2 e5 e2 e0 db db d8 da db d5 ce cf c6 d0 c9 c5 c5 bb be b6 ae b1 a7 ac a4 a1 9e a1 9b 93 9b a0 93 9c 9a 91 8d 90 97 8b 83 8b 85 80 76 75 6d 70 6f 6f 69 68 60 6b 84 8d 81 61 37 32 21 29 18 10 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0b 18 28 39 4b 5b 77 84 90 82 75 6f 77 70 61 66 6c 75 75 76 7f 7c 85 86 8b 88 8d 82 84 8a 91 96 95 9b 98 9f 9d a4 a8 ac
 b8 bd b7 c1 c9 cb c6 cd d0 d9 d6 d8 e3 df e9 e2 e9 e1 f0 f5 f7 f5 f9 f7 f4 f6 fa fe ed f2 f0 f1 f3 f4 f7 f6 ef e7 eb e6 ea e9 e3 f1 ee ea f0 ea f2 f0 f8 f1 ef f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 e3 de de e5 e1 e1 e1 e2 e1 de e6 e8 ea e9 e3 e1 ec ea ea e4 eb ee ea ed e5 ec e8 de e2 db e2 de de da d8 d8 dd e0 d2 d3 cd c7 ce d1 c6 c6 b7 bb b3 b5 af ae b0 ae a4 9e a2 95 93 9a 9e a2 a1 98 8f 8d 96 90 87 92 8b 87 86 7b 75 70 68 71 72 64 65 6e 6b 83 93 7e 60 4b 3a 3c 31 22 10 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 07 12 12 2d 3c 4f 5f 7a 8b 98 85 71 6a 6a 5f 5e 66 6a 70 6c 71 75 7f 85 87 88 8a 86 87 88 88 95 92 96 99 9c 9f a5 ab a9 af b3 ba b2 b9 c1 c8 c9 cc cd d6 db da dd e6 dc ec eb e5 f2 f5 f2 f9 f6 f6 f3 f3 fa f6 f7 f0 f4 f0 ea e9 ea eb ea e8 ee e7 ec e9 ee f4 f1 eb e9 ee f3 ef f6 f5 f9 fd ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 dd e1 d8 dd e3 de e0 e7 df eb e8 e3 e9 e9 e3 e7 eb e7 e2 e7 e4 e8 e3 e8 e4 e8 ea e3 df e0 e1 e3 d6 d8 d5 e1 d4 d7 c8 cc ce cb c9 c4 c2 c1 ba af b4 b6 ac b0 ae a6 a9 9a a0 99 a0 9d 97 9c 9b 9d 9e 94 94 98 8c 8a 8f 83 86 76 75 7b 6f 70 65 6b 70 6a 7a 8d 92 81 66 54 4e 45 3b 20 16 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1e 26 40 55 66 73 8b 99 8e 74 5f 59 5a 5a 64 64 65 66 6b 73 7c 83 82 87 8a 87 90 91 94 91 93 96 97 9a a5 ab a1 9e ae b2 b2 b6 b6 bb c9 c1 ce d1 cb d8 d3 d5 de dd df ea e5 f3 ef f1 f0 f2 ec f3 f8 f5 f6 f2 ef f3 eb f0 ee ee e8 e6 f1 e8 ec f3 ec e9 eb ec ec ef f2 f4 f3 fa f8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff bf ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb dc e0 d3 de d7 df dc df d9 e8 e1 e0 e0 dc e5 e4 e1 e4 e4 e5 e7 db e0 dd e1 dc e6 e3 e0 db db d4 d6 d8 d0 d3 cc ce d9 c8 cc c5 c8 c5 bf c5 b9 b7 b3 b3 ac af a4 ab a0 a4 9a 97 99 9a 9e 97 99 9e 9b 9a 97 93 8d 8c 8a 90 82 84 78 78 6b 75 6b 6d 66 6e 70 7c 8e 92 87 71 5b 58 46 34 27 1d 0f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 11 1e 31 3f 55 6f 82 8b 9a 98 79 5e 50 5e 58 64 6e 62 6e 72 6b 76 70 82 8e 84 97 91 88 92 99 9b 9a 9a a1 a2 a4 a7 a7 ad
 b2 b2 b6 b4 c8 bf c5 ce c8 d5 d5 d4 de e2 e1 ec e9 ea ef ed f3 f5 f3 eb f7 f0 ef f6 ef ed f2 f1 ef ef ed eb e7 e5 e7 e7 f0 ef ef ef ed e9 ec ee e8 f0 f7 fe ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 e1 e4 d6 d5 d5 db df da dc e1 e5 dc db dc e3 e2 e0 e5 e5 db de e8 e3 e2 e8 e3 dd e1 dc de d8 de d2 d7 ce d3 d2 d3 d5 d8 c5 d1 c8 bf c0 c8 c4 ba bc b9 b5 ae ac b0 b2 a1 a5 a3 a1 9b a0 a1 95 9b 9d 9b 98 95 9d 8e 94 86 88 7c 7e 7b 73 70 6a 6a 67 69 6e 69 7e a1 93 8e 79 6b 5d 4b 4a 36 22 18 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0e 17 18 2b 3d 56 6f 7b 94 a2 99 7c 61 5b 5a 5d 62 63 63 62 6e 71 7f 77 88 84 8e 97 8f 95 9a 9d 9a 99 9b a0 a4 a1 a8 9c b5 b4 b3 b2 b7 c0 bd c6 c1 ce cf d4 d0 df df e5 e9 eb eb f0 ed f3 f6 f8 f1 f7 f7 f5 f9 f3 ef e6 ef ed ea e7 f0 e8 ec ea f4 f6 ef ef e9 e4 f0 e9 ec f6 f3 ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 f2 f6 fe f8 ff ff ff ff ff ff ff ed e7 e8 fa ff ff ff ff ff ff ff ff ff e8 de d0 d9 d6 df d7 db e0 da de da d9 e2 e3 e1 df e4 e3 e8 e2 d9 e1 e0 e0 e3 e3 dd d7 d5 d9 d4 cc d1 d2 d1 d3 d4 cb c9 d5 c5 c7 c9 bf bc c1 bd be be ad ae ae a6 aa a5 ad a3 9f a3 a0 9a 9a a5 9e 91 9b 99 96 97 8f 86 8a 8c 89 84 79 7c 73 6d 6c 6d 64 68 70 81 95 99 8f 89 70 65 53 3c 32 2b 13 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1e 2d 48 55 72 84 8b 9d 9f 77 5c 59 5f 5c 5a 63 6a 67 6f 6d 7b 77 7a 88 82 8e 8f 98 a4 9c a4 a2 9d a1 a0 ab a5 a7 ad ae ad b8 bf c2 bd c6 c8 cd c6 d2 d5 d7 de e0 ee eb e5 e5 ea f2 f3 f0 ec ed f5 f9 eb ed ea e9 e9 ed ea eb e6 e5 e3 e6 ea ed ea e7 eb ea e9 eb eb f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec d7 dd d6 d7 d2 d8 dc f3 ff ff ff ff eb d1 c3 c5 d6 f4 ff ff ff ff ff ff ff fd e5 d6 cc ca da d5 d6 df e2 db dd e2 de e4 d9 da dc e1 e4 de e0 d3 d7 e1 de da d9 d4 d9 d6 d3 cf d0 d0 cc d3 cb c6 d0 ce c4 c3 c1 c8 b3 c1 ba b4 b3 b3 b5 b3 ad ae a8 a8 a6 a0 a9 a0 99 96 9a 96 a5 97 96 97 8e 93 90 8f 8c 8c 85 7b 7f 7c 77 71 73 62 63 68 6b 81 92 a3 98 8a 76 69 52 47 34 22 16 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 1a 22 2d 40 58 76 89 95 a8 9b 77 5b 50 5f 60 60 6c 60 6e 6e 6b 78 7f 79 80 86 94 98 97 9e 98 a5 a6 a0 9d 94 a6 a4 ae b4
 ba b7 b7 bc c5 c7 cc c5 cf d0 cb e2 dd d7 e4 e9 e7 e9 ed ed f3 f2 ed f2 f8 f1 f6 f1 ec ec f0 f0 ed ec e3 e8 e6 ed f4 f4 f3 eb ed e8 f1 ef ef f0 fb f7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff df d0 b8 bd b1 af af b2 b3 c5 ea ff ff ff da bf b5 ab c1 d2 e8 fb ff ff ff ff ff ff d5 d4 c7 cc d4 d5 d9 d7 dc de da de d5 df e6 e1 de df e2 dd da d8 d3 dc d6 d4 d1 d7 d8 d2 d9 cb d0 ce ca c6 cd be ce c1 c5 bf c0 c0 b5 ba b8 b2 ab af a5 af a7 a6 a5 aa ad a6 a3 a6 9f 9e 97 92 9d 8f 99 8b 88 93 91 91 85 90 85 8d 82 7d 76 7b 6b 63 66 61 5a 6b 8c 94 9e 84 7f 65 5f 51 3a 36 1b 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 1c 22 32 4b 5b 7c 8f 9a a0 90 6e 5f 54 62 61 5d 67 64 68 74 6c 72 7a 7c 7f 8a 8f 97 9f a1 a3 aa aa a4 ad ad ad a9 b2 a5 b0 b9 b5 b2 c9 c2 c8 d3 d8 c8 d8 d9 dd d8 e0 de e4 ed e8 f8 f6 f5 f9 f8 f4 f8 f5 eb f3 ef ef e9 e7 e9 f0 e9 ed f0 ee ed f7 eb f1 ea f3 f3 ed f8 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e4 d9 ce b7 ad a3 a3 a1 9b 9a ac d0 ef ec f0 b9 b5 aa 9f ad be cd ed f8 ff ff ff ff f6 cf d0 c1 cc d0 cd cd d3 da e3 e3 e2 d7 da d8 d6 da dc d6 d7 dc d3 d0 d5 da de d4 d5 d1 d4 d3 c9 cf ce cb c6 c3 c4 c2 bf bc b2 be b5 b3 bc b0 b6 b4 a7 af a5 a7 a4 ab ac a0 a6 a0 9f 9c 95 9b a0 9b 9a 93 94 87 8f 8c 92 99 84 89 89 7f 7e 76 74 6b 69 64 6b 56 63 7b 8e 94 98 7f 76 56 4a 45 2d 20 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 14 1e 28 45 5a 70 94 a8 a5 84 69 54 5b 59 60 5d 68 6a 6d 70 73 69 72 74 84 8f 8d 8b 9a a4 a5 a9 aa a9 a9 af ab b7 b4 b2 b6 b4 b9 bb c9 cb cc d3 d3 cd d2 d7 db dd de e4 e0 ef ec f0 f6 f5 f3 f8 f7 f0 f4 fa f8 f0 e8 ef ea e7 ea e8 e7 ef ed ec ee f0 f9 f4 f7 f9 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f0 e8 da ca ca bc ad 9b 9f 96 8b 8c 9f b2 c2 c7 c1 ab 9c a5 94 a4 b5 c9 d5 e8 e4 f5 ff ff f7 d0 c9 c4 cd ce d7 ce ca d4 cd dc da d4 dd d6 d5 dc d4 d3 da d2 cf d2 d9 ce d2 da cf d1 cf d1 c3 c9 cc c1 c0 bb c1 b6 c2 bf b5 be b6 ad b5 b0 b3 ae a8 a9 a5 a8 a8 a7 a0 a3 aa a0 9b 99 95 95 93 95 95 91 96 8f 91 8a 8e 87 8f 8a 83 7a 74 6c 70 65 69 5c 59 57 5e 75 93 9a 92 84 76 5b 4f 4b 28 23 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 10 19 2d 3c 5a 75 8d 9d 9b 82 6d 5b 5a 63 63 64 5f 69 6d 6c 70 79 6f 76 84 88 8f 90 8e 9e a3 ae b0 b5 b4 b5 b4 b1 bb b2
 bc b5 be c5 c4 c9 cb ce c9 d3 d7 dc e0 df e7 e0 ef ec e7 fa f4 f4 ff f7 ff fb f9 f3 f5 f0 f2 f7 ec eb ec eb f2 f2 f1 f3 f1 eb f5 f3 f5 f8 fc fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 d0 d2 b4 a8 a0 9a 94 90 89 84 6a 69 7c 7d 8c 8f 88 89 7e 8b 86 8f ae c3 ce d2 d1 e4 ff ff ee cd c1 c4 ca ca c9 d3 cf d7 d1 d2 d8 d5 dc d5 d9 d7 de d1 e2 d8 ce d0 cc d1 cf c8 cb c8 c8 d3 c2 be c0 bf c1 c2 c3 b7 c0 b3 b3 b7 b5 b0 af b2 ae a8 a5 ad a9 a5 a7 a4 9e a0 a4 99 9e 99 97 95 99 98 94 93 91 85 8e 89 89 8d 88 81 88 80 75 71 71 62 65 61 61 5e 62 6c 88 9a 8b 83 77 65 56 42 39 1f 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 22 2c 44 5b 77 8e a2 9c 79 66 60 5b 5d 5a 66 70 6b 69 73 6f 76 77 7b 7b 8c 8c 89 8f a0 a5 ae ad b3 b0 b3 b3 ba bf bf ba bb bf cc d0 ca cd d5 d7 d4 d0 d5 db df e9 e1 eb f0 f4 f4 f5 f4 fa f8 fa ff f4 f6 f4 f1 f7 f1 ef ee ef f1 ef ef f9 f7 f9 f1 ee f7 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fd fb ff ff ff ff ff ff ff ff e5 cb b7 a4 88 7e 74 5f 6b 65 5b 60 60 57 56 60 65 65 6c 66 61 5c 6f 78 8d a0 ab c1 c5 ca f5 ff e7 cd c7 bd ca c9 cb d3 c8 ce d5 ce d5 dc d3 db d1 d3 d8 ca d4 d0 cb c9 cc ca cb d1 c5 cb bf c6 be bf bd bb c2 bd b0 bd b6 bb b4 ac b0 aa af ad b5 a3 a9 ac a3 9c a1 9a a1 98 95 95 94 9e 97 9b 92 90 90 8e 88 8c 8a 88 8b 8c 8f 84 89 7c 7c 71 72 66 64 62 5a 55 63 75 8e 98 96 85 80 64 5f 40 3a 2e 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0c 16 2a 44 61 7b 91 a1 a2 7d 65 62 5b 60 5d 66 69 6f 6c 67 71 72 7c 78 7d 8a 89 93 97 95 9d ad a8 b1 b8 bd bc b8 b7 b6 c7 bc c7 c5 d2 c4 d3 d3 d5 e0 df dd e0 de e0 ed ea ef f2 f2 f6 f6 fa f9 ff ff f6 fc f5 f4 f5 f6 f1 f1 f1 f6 f6 f8 f9 ed f5 f5 ff fa f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fe ff ff ff ff ff ff ff ff ff f8 cf af 98 82 66 60 5b 56 4c 53 4c 4b 44 45 4b 4b 4d 4f 4d 48 48 57 59 58 65 7c 8b 95 aa bb df ff ee d2 ca be c0 c5 ca c9 c9 d2 d8 c9 d1 d6 cf cc cc ca d4 cf cf cb cb c3 cc c4 ca c1 c4 c3 c3 be bf b6 b4 b2 b4 b3 b8 b3 b2 b5 af af ae a4 ad a5 a7 a1 a0 a1 a3 9f a2 97 a2 98 95 9d 9d 93 95 94 91 8c 8f 90 93 8e 8d 8a 88 89 89 8b 86 7c 7d 71 6f 6c 5f 5e 5d 5b 5e 64 84 9e 96 89 7e 5f 57 3d 3f 20 14 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0b 17 1a 29 44 56 72 8f a2 9b 81 6b 63 65 6a 6c 6d 68 6c 71 74 77 74 7a 7b 7c 80 84 8b 99 9c ab ae b4 b3 c2 be ba c2 c2 bb
 bd bf c5 c7 c5 d8 cb d4 d9 dc d8 df db e0 e4 e6 e5 e8 ee f2 fc fa f6 f6 fb fb f6 fb f6 ef ed f3 f4 f0 ed f0 f4 f5 f7 f5 fb f9 f8 ff ff ff ff ff ff ff ff ff ff ff f8 ff ff f9 fe f5 f4 f4 fd f5 ff ff ff ff ff ff e7 b4 94 7b 59 55 4c 43 48 41 48 42 44 41 3d 3f 47 40 4b 43 42 3c 49 4b 4b 50 5f 67 73 91 a3 d0 fa e6 cc b9 b7 c3 bf c5 c7 cb ca ca d4 cd cb cf d2 cc d2 d0 c1 c8 ca c4 c4 c4 be c6 bc c1 b9 b9 ba bf b6 b4 ae b0 b6 b0 b0 a9 b2 af a8 ae a8 a1 9f 9f a0 9d 9f 99 9a 94 9b 96 95 98 9d 99 95 8f 98 8b 90 86 84 87 83 8c 86 89 87 8f 8a 84 75 75 71 70 6f 66 66 60 5b 61 75 8b a0 97 8a 75 6a 58 4c 3b 23 0c 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 12 16 2a 37 5e 6b 85 a5 a4 89 6e 5d 5f 66 6c 6c 6c 6b 6d 70 7b 78 76 77 7c 86 87 8f 90 9a a0 af b3 b4 c1 c0 c1 c4 c6 c1 c1 c1 cc c3 d3 cb d0 d6 dc d7 de db e1 dc db e7 e6 ed eb f2 f1 f8 f9 fd f2 f4 f6 fc fa f9 f3 f6 f4 ee f6 fa fb fe ee fe ff fe ff ff ff ff fe ff ff ff ff ff ff fe ff ff fa fb fc fa f3 ee f8 f5 ff ff ff ff ff ff d0 99 78 5c 4a 3f 44 50 48 3c 3d 37 35 41 38 33 42 3c 36 39 43 43 40 44 48 4a 48 52 64 75 93 b9 e4 e4 ca b9 be b7 ba cb c5 cb cb d5 ce d5 cf cd cd c9 cd ca c7 c8 c4 bf c1 c0 bd c5 b7 be bc be b9 b8 b7 b0 a7 b2 a6 af ae a4 b2 a5 a1 a8 a5 a0 9d a0 98 9d 9e 94 9c 90 91 95 97 93 98 8d 93 8f 94 8a 8e 8a 8f 8c 8b 8c 8f 84 86 8b 7d 84 7d 7d 72 64 6e 68 68 61 5c 60 71 8c a3 93 85 81 68 57 51 41 25 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 12 10 20 38 4c 61 81 a0 a0 95 7a 69 68 64 6a 65 6b 74 6c 6c 73 7b 79 77 7a 78 81 8e 91 96 a6 a6 ad ac b7 bf b9 bb c8 c8 ca c4 c9 ce d4 cf d8 d5 d7 e1 d5 d8 df e0 e2 e2 e9 f0 f1 fb ff ff f6 f6 f5 f6 f4 fa fc f7 f9 f9 fd f3 f4 f9 fb fe f8 f8 fb ff ff ff fc ff ff ff ff ff ff ff ff ff ff ff f7 f4 f7 ed ef ec ea e7 ff ff ff ff ff e7 ba 84 5c 4e 48 3e 3d 3a 33 3e 33 2c 35 31 28 27 2b 30 2f 36 2c 30 34 3e 41 47 49 4e 54 64 74 a9 d7 e4 cb c0 b2 bc ba c3 c5 c1 c7 c7 c8 d0 c8 cb c6 c6 cb c5 c6 c0 bb ca bf bb bc bc b3 b4 b3 b2 ad ad a9 b0 af ac a7 a0 9e a5 ad 98 a0 a3 9b 9c 9e 97 95 99 90 95 93 90 90 8f 98 8f 97 91 8a 87 84 84 8a 84 85 86 80 8d 81 82 8a 87 85 86 74 7f 7e 6e 6a 62 5e 5b 5b 62 70 94 93 a0 8c 7b 6c 61 4b 36 27 13 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0d 19 1c 35 45 68 83 99 a8 90 7a 68 65 6c 6b 6d 6e 6e 71 75 71 6e 7b 81 78 81 86 82 94 90 a1 a5 a5 af ae bd c1 bf bf c9
 c4 c6 cb cb d1 d2 d0 d6 d8 d3 d7 da dc e1 e2 e1 e4 e2 f7 ff ff ff fe ef f0 f9 ef ec f6 f8 f0 f4 f6 ef f7 f4 f5 f7 fb f9 fe fd ff ff ff fd ff ff fb fe fe fc ff fe f7 eb f4 ee f4 ea ef e8 e7 e9 f8 ff ff ff da bc 96 6e 4b 42 3a 30 32 33 25 31 23 2b 25 28 2a 28 1f 24 1b 25 25 2d 2f 32 3a 42 3e 41 46 5a 63 99 cf db c4 bd b4 bb bf be c1 bf c7 c7 cb c6 c9 c2 c4 c9 c0 c1 b6 b7 b9 b6 be b6 b4 b7 b1 aa a8 af a5 ad a2 a7 a4 a4 a7 a3 a5 96 a4 99 98 9e 91 9a 95 8f 94 91 8a 8f 8d 90 8d 8d 92 85 88 8c 8c 86 89 8a 89 82 81 82 80 86 8d 84 8e 8a 83 7e 80 79 70 67 66 5c 56 57 58 55 6a 90 9a 95 8c 7d 6f 5d 47 33 1e 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 12 0f 1e 35 46 61 7f 96 a5 9e 84 73 64 65 6a 70 6d 75 72 6d 7a 7a 78 7e 84 86 88 93 94 98 a4 9b a9 ad b7 b9 c0 bc c4 c5 c9 cc c5 cf d2 d0 d4 d5 d5 d5 da d5 db db db e5 e4 e4 f5 ff ff ff ff ec f2 e5 f1 e8 f3 f1 f2 f4 f8 f3 f7 fa f2 fa fe fb ff fe ff ff fe ff f7 fb fd f4 f3 f5 f3 fa f2 f3 f5 e5 eb ea e4 e0 e6 e3 f0 ff ff ff dc 9f 77 57 45 3c 38 2c 2e 2a 2a 2c 24 25 1a 19 21 20 1f 28 1f 23 27 29 27 28 2e 36 36 39 43 52 6b 89 c6 d9 c0 ba b3 c1 ba bc c5 c4 c3 ca c9 c7 c5 ca c2 bd b9 c4 b9 b5 b5 ba bc b1 af ba b0 b0 ac ac b0 a9 9f a1 a7 a5 9c 9d 9d 9a 97 9e 9a 9b 95 96 8b 8b 96 91 8b 93 8c 8b 87 87 8e 87 8c 8d 8a 86 8c 81 88 84 88 8b 84 8e 85 87 84 8c 85 82 80 79 70 68 62 60 59 5a 59 56 65 89 9b 9a 8c 81 6e 5f 4f 42 1d 16 08 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 15 21 2d 43 62 75 9e a0 9d 8f 75 67 6b 6d 69 75 73 70 75 75 79 77 7b 80 83 8f 8b 93 9a 98 a1 ab b0 b3 bf b9 bd bf c2 cb cd c8 ce cc d2 d2 ca cf d4 d0 d5 d8 df db e3 dc d9 eb f4 f7 f6 ef e5 ed ee e7 ed ef ed f5 f0 f0 fa f5 fa ec f9 fe f7 ff ff ff ff ff fe ff fc f9 f6 fa f8 f3 ee f5 ee ef f0 e9 eb e6 e4 e0 e3 e9 ff ff ff e2 90 69 53 3c 2e 25 22 1f 24 20 23 24 1f 15 18 1b 1f 1d 1b 1c 1c 1d 1d 28 28 26 2f 2a 34 41 48 62 83 bf d6 bf af b0 b9 b9 b8 c6 bb c1 c6 bf c6 c1 c7 c8 c2 ba b2 b6 b8 ac ae aa b2 ab af ac a6 aa a3 a9 ab a4 a3 a4 a5 a0 9f 9b 9b a0 9a 95 97 91 93 95 88 91 86 87 8b 86 85 89 89 8c 85 8a 93 84 81 85 88 8a 81 83 8a 87 8d 8f 8e 8c 87 84 7c 78 74 75 71 5d 61 61 5c 60 61 5d 7e 9b 9b 8e 86 71 60 48 31 24 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 15 1d 30 4c 5b 77 88 a3 a4 86 71 6a 6e 66 6a 6f 6f 73 6f 79 7a 82 7f 7d 86 8e 8e 9c 96 98 a6 aa a9 af b8 bb c1 c1 c3
 cb c4 cc c4 c5 cf cb d2 d3 d2 d5 d5 db d4 da dd d9 db e1 e0 e3 ea e6 e5 e0 e3 eb e6 e2 ef ee ec eb f1 f5 f5 f4 f5 fa f7 ff f5 f5 fc f8 f8 f4 f9 f0 f5 f5 f5 f1 f0 f3 e0 ec eb de e7 de e2 e6 df df e9 ff ff d9 81 5e 4b 34 29 20 1b 22 1e 1a 19 1e 1c 19 18 14 17 16 1f 09 13 18 13 1d 1f 16 1d 25 29 30 44 59 7f b5 cf b6 af af ae b1 b7 c3 c4 c1 bf c1 bb bf ba b7 b9 bb b4 af b5 b0 ab ab ae af ab ae a8 a8 a8 a5 a1 9f 99 a0 a2 9d 99 a2 9f 98 93 95 8e 88 8d 8a 83 92 89 80 86 83 85 81 86 8a 85 85 84 7e 85 80 83 8c 89 87 87 7e 86 91 89 8f 84 81 81 71 76 65 66 67 63 5d 4f 5d 5e 62 6f 95 98 90 7f 6c 5e 4c 3d 29 13 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 09 0f 28 34 49 5e 76 88 a3 aa 94 7d 73 6e 67 6c 72 71 7b 75 7d 7f 7a 84 7f 84 8a 89 94 9a 99 a1 ab a8 b1 bf b5 c3 ca c5 c6 c6 ca c9 c9 cb d0 cf d0 cc d2 d5 d0 d2 ce d7 e0 d4 db d7 da df e4 df e2 df de e5 ec e9 e8 e5 ed f4 ed f5 ec ec f2 ed f6 f3 f1 fc f3 f7 f2 ee f3 f5 f5 f4 e6 e8 e7 e6 e1 e3 e5 e1 e4 e2 d0 d4 db df fc ff d2 82 5a 3e 2a 29 25 19 1e 14 19 14 0e 0e 0f 10 04 15 0f 11 16 0f 0e 14 17 22 25 21 1d 23 24 38 5e 7f bb c6 b5 ab ab ae b0 c1 bc c0 c3 c3 be c8 c0 c4 c1 bb bd b5 b3 af aa b3 a8 ad a9 aa a2 ad b1 a8 a7 a5 9a 9b 9f 98 a0 96 8d a0 a0 94 9d 90 90 88 8e 90 85 89 85 7d 84 83 84 83 86 78 7f 87 7d 84 88 7f 86 80 86 89 86 8d 90 8d 8a 82 7b 7c 71 6a 6f 64 67 5d 55 64 56 5a 5d 73 93 94 95 83 70 61 50 36 2c 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 27 31 4a 5f 74 8e 9c a8 a0 7d 71 6e 6d 6f 77 7a 78 73 7d 80 81 81 87 8a 8d 97 98 a0 95 9b 9d a3 ad b7 bc bd bf c2 cb c5 c9 c7 c9 c7 c9 cb cf ce cb ce cc d4 d0 cd ce c9 d2 d3 d4 d4 d9 db d5 dc e2 d3 dd e2 da ee ec e8 e8 f3 ec ef f2 ee f6 f2 f7 f3 ed ef ec f6 eb e3 eb e4 ec ec e6 db e5 e0 e1 db de dc d5 d2 d9 d9 e4 ef ae 79 5a 37 26 21 19 0d 16 0d 14 10 0a 0f 0d 13 0f 0e 0b 12 07 15 13 16 12 19 19 1e 1c 22 29 3b 57 7e b2 bf b0 ae ae b6 b4 b4 c3 bb be ca c7 c2 bf c0 c2 b8 b8 b1 b3 b7 b0 b2 b2 b5 a0 ac 9e 99 9e a2 a0 a5 9f a1 9d 9d 9a 9a 9c 97 9f 96 96 95 93 90 91 8a 89 89 85 84 84 7d 85 7f 84 89 85 8e 83 7e 81 89 80 8f 89 89 8c 96 90 92 83 82 7a 7b 70 6d 6b 5a 5d 62 56 5c 63 5a 5e 6c 89 92 91 84 70 64 4b 37 1d 11 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 0c 0e 1e 2f 49 61 71 8a 9c a3 a4 7d 6f 6a 69 73 78 79 78 7b 78 7e 85 84 8a 92 8b 93 98 9c 9d 9e a0 aa ae b0 b0 ad bd b2
 c4 c1 bb c4 c5 c5 ca c7 c6 c9 c4 c0 c3 c7 c3 c5 cf cb c9 c6 d3 ce d6 d3 dd dc d1 d6 d5 d5 d6 d7 d9 d9 e0 ef ea e9 ec e7 e7 ea ea f7 ec e3 e9 ea e8 e9 ee e4 e1 e2 e2 de dc e0 db e0 d5 d9 d7 d4 ce c9 e0 d8 b2 78 57 2b 28 19 15 0e 16 16 0b 0e 08 0c 06 09 08 0e 0a 0d 08 0d 0b 11 14 08 0d 10 18 20 29 28 56 7b b4 b7 ae a9 b0 b1 b5 b3 bc c4 c1 c1 c0 bb c0 b6 c1 b3 b1 b7 b2 a9 ac ab a8 a6 a4 a4 9f 98 97 9d 98 9d 9e 9d 96 97 95 95 a1 96 9c 92 91 96 96 94 9b 8f 90 8d 89 8b 87 82 83 81 7e 83 7a 7d 7c 7d 85 74 80 7e 8a 8e 8c 92 8c 81 7f 7f 7c 75 71 65 69 64 61 62 61 5a 53 55 61 65 85 94 91 83 6a 59 4a 2b 1f 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 07 1b 1c 31 45 61 78 94 a1 a0 9d 84 70 71 6f 70 76 7c 7e 81 7d 87 85 87 81 90 8a 93 8e 97 99 9d a2 a3 a6 ad ae b4 c2 bf bf bb bc bb c1 bf bc c0 c0 bd bb c6 be be bf c4 c9 cb bc c9 be c9 cf cd d5 d2 cb cc d7 d3 d4 d3 de d8 dd e0 e3 df e6 e4 e2 e4 e7 e5 eb ed e2 e9 e2 da e6 df dd e0 e4 dc da dd d8 d5 d3 d8 d9 d0 c6 d0 cc c5 b0 76 5a 2e 16 0f 0b 17 0d 07 08 0e 11 0b 06 06 08 05 06 05 0a 0c 11 06 06 0f 10 0f 17 11 1d 2a 4d 87 ad b2 b1 b9 af b8 b8 b8 c8 c2 c6 c4 c7 c1 bc be b6 b9 b7 b3 b2 a8 a6 a7 9e 98 93 a1 98 99 8e 8f 8e 8e 98 99 95 9d 93 90 8e 8e 95 8d 8b 8b 90 8e 8e 8d 9b 92 90 96 8f 98 86 8d 84 7f 7f 7b 7b 80 83 84 8c 7d 89 8a 8a 8f 87 87 84 7a 75 74 76 6d 62 66 5f 5d 5e 5c 53 5f 5e 71 80 94 8c 86 65 5e 49 31 20 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 0c 0c 25 2e 45 62 7c 8e 99 a7 9f 7d 70 74 6c 77 7a 7f 80 79 7d 84 82 8b 92 8f 94 95 94 96 a3 a1 a0 a2 ac ac a8 b9 b6 b4 b3 b6 be b9 bf bd c0 c5 bd bb c2 bb ba ba bb bb bd c5 c4 c5 c4 c8 ce c6 ce c5 ce cd d3 cf cd d5 cd d9 d5 d9 e1 d5 d6 dc e7 e0 e2 e7 e6 e4 e1 de e5 de db e1 e3 df da d8 de d4 d3 d2 cd d4 d3 d0 d1 cd c4 c2 a2 7c 54 27 14 15 06 09 0a 0c 0e 0c 06 0b 0b 0f 0a 0c 07 06 0d 09 09 0a 07 04 0e 1c 1a 12 1a 26 4d 86 b3 b6 b9 c1 ba b9 bd bf c5 c2 c2 c7 c4 bc bd bd b7 b3 b0 af a6 a6 9d 98 95 94 99 94 92 88 8e 86 8b 92 8c 94 8d 8c 96 8e 87 94 93 8d 87 91 8b 8a 85 84 89 92 93 91 92 92 91 8b 84 86 85 83 76 87 7f 82 87 8f 91 8f 93 86 88 85 82 76 77 6e 65 69 68 5f 5e 5a 65 60 5f 5f 66 6a 80 98 95 89 6e 5a 49 35 29 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 16 1b 2f 47 65 73 8c a3 a7 97 79 73 6a 6f 6d 75 7e 82 7d 86 83 85 8f 8f 8b 94 95 8b 90 a0 9a a1 a2 a5 ac b1 ad b6 b6
 be b5 b5 bb ba b9 b3 bb b8 bd bc c1 b5 bb b5 ba bd b7 b6 bf c3 c0 c2 c7 c5 bd c8 cc ca cb d3 c5 cf cc cc d9 d3 d0 d0 d5 d4 d6 dd da d7 da db d9 d9 dc d5 d7 d8 dd d8 d6 d4 cf d5 d7 d1 d1 c8 c5 c1 c9 bb bb a2 78 4d 1d 13 0a 06 05 03 0a 06 05 03 06 06 0a 07 00 06 0a 07 08 0b 05 0c 0e 10 12 0d 0e 13 25 44 8a b7 bd c6 c7 c6 c7 c1 d0 cb c6 c2 c0 b8 bf bc bc b4 b0 af a1 a0 a4 95 95 8f 84 92 91 92 81 87 8f 82 8d 7c 85 86 88 85 8d 88 8b 8d 86 88 84 8c 8c 83 87 8a 8d 8f 8e 90 94 93 91 8a 83 83 7e 7a 7f 88 8a 86 8f 8e 8b 8c 80 89 7e 7c 6e 71 71 65 69 5e 61 62 65 5f 64 5f 60 61 69 81 94 8d 8a 6d 5c 48 31 1b 06 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0e 0a 23 34 3f 5f 6f 86 9f 9a 91 79 70 74 75 74 7d 7c 7d 85 85 85 8b 8b 92 94 91 95 9a 96 9b 9b a0 9f a6 b7 a6 ad b6 ac b5 b1 b5 b4 b7 b3 ba be bc b3 b9 b1 b8 af b5 b8 b5 b5 b6 bb c0 ba ba b5 c4 c3 bb c2 be c2 c1 cb cc c9 c9 cd cc c6 c7 d4 d3 d0 d8 dc d3 d6 d6 d4 d3 d3 cd d7 d2 d0 d6 cf d3 ca d7 d2 cb c5 c9 bf c4 c1 b5 ac a3 86 4f 1f 11 0d 06 05 03 0c 06 05 04 00 06 05 05 05 06 05 03 01 06 05 03 06 08 05 14 12 11 18 3c 87 b5 c3 d1 ca c9 cf c4 c6 cb c3 c2 bd b6 af b8 b4 ab b0 a3 aa 99 9d 90 8f 8a 8e 8e 83 83 86 83 88 83 8b 87 81 87 84 7e 82 85 8b 8a 81 8a 79 82 86 7f 84 80 8b 89 90 93 99 9b 93 96 8a 92 8e 8c 8e 91 8f 88 9b 85 8c 7d 84 88 82 84 71 6f 6d 6c 69 64 61 61 58 61 64 60 60 68 72 77 8c 8b 7e 6b 5d 40 2d 1b 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 09 17 1d 2b 46 5a 71 8b 9d 9a 8b 75 6e 6f 72 6b 7b 7e 82 84 85 87 8a 8e 8b 8f 90 95 96 8f 97 97 9c 9d 9e aa a6 a2 ab af b0 ae b8 b8 af b3 b0 ba c1 b1 b2 b1 ad a7 b4 b5 b9 b2 b3 b6 b5 af b6 ba b9 bd be bc c0 c2 c4 c3 c7 c6 c4 c9 ce c7 cb ca d1 cf d6 c8 d2 ce ce d2 ce d0 cd ce cb d4 d5 cf d0 c7 c9 c8 c5 c7 bb be c3 bd b7 af 9e 71 49 1f 08 10 0d 0a 05 00 06 05 07 07 06 05 06 07 06 0a 04 02 06 09 05 0b 0e 19 0e 10 08 1a 32 80 b7 c3 c6 c8 bb c2 b8 ba c1 b7 b1 b0 ab b8 a6 a7 a6 9d 9d 9e 9e 99 96 92 8d 8a 88 87 86 8c 87 7c 7e 81 81 7a 7c 83 75 7b 80 7b 8a 7c 79 82 85 80 7f 86 83 84 8a 8c 8d 99 9e a0 a1 97 9a 8f 8e 8f 85 8a 90 8d 8f 8f 7e 8f 80 7c 7b 7c 77 70 64 6a 66 68 67 5f 62 65 67 64 69 71 81 8e 8b 83 66 60 43 2e 20 0a 0f 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0c 15 19 3b 48 5a 74 84 96 94 83 72 6d 70 72 75 79 7d 7c 81 86 8f 8d 90 95 8f 8e 92 90 98 99 95 99 a0 9d a5 a0 a5 a7 af
 ad a9 af b1 ac b4 b3 ab b3 af b0 ae af ac a9 ad a9 a6 b5 b3 b3 ae b0 b2 bb b9 c0 b9 c0 c2 b1 bf c2 c1 b9 c5 bc c1 c1 c6 d1 c6 cd c5 cb c0 cf d0 cc cd d0 c5 ca c7 c7 cd c8 c6 bd bf be bf bd b7 b8 b0 a6 a9 a0 7c 4f 23 09 07 06 05 03 01 06 05 03 0b 06 05 06 00 06 05 03 05 06 05 03 08 06 14 0e 07 07 12 35 72 ac b5 b7 b5 b4 b0 aa b5 a9 a7 a3 af a4 a1 a9 a0 9b 9a 9b 90 91 94 8f 8d 87 90 8d 8a 83 86 84 87 81 88 86 84 7e 82 7e 82 83 82 7d 82 86 7e 77 81 80 85 8c 8a 87 97 8a 95 90 95 9b 8d 88 89 89 8b 85 7e 84 86 8a 8b 8b 82 81 7a 76 71 79 6a 6d 67 65 64 6a 63 62 6b 68 65 66 65 77 8b 8e 84 69 59 45 2c 11 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0b 12 1b 33 43 54 77 89 94 93 7b 70 6d 6d 6b 6c 78 7a 75 80 86 85 89 90 91 90 99 95 8e 97 95 99 96 93 93 9b a5 99 a2 a8 a8 a4 ad ad aa ad b3 a6 ac a4 af af a6 ad ab a9 aa a9 ad b0 b1 ae b1 b5 bb ab b6 b8 bd b3 b6 be b4 b7 b7 c4 c2 c1 bd c4 c3 b8 bc bb cb c1 c3 c1 cd c6 c6 c3 bd c0 c2 c2 bd bf bd c4 b8 c1 ba b1 ab aa aa 9d 96 78 51 1f 05 01 07 05 03 00 06 05 03 02 06 05 03 00 06 05 03 01 06 05 06 00 06 08 0e 07 07 10 2f 7a a3 ae b3 ac a8 ae a0 a2 9e a4 a0 a4 9d 99 96 8f 9a 91 92 91 8f 8f 97 87 8a 84 83 84 85 89 84 7f 81 7f 84 8e 86 8a 84 84 80 86 85 7e 82 87 80 83 87 88 85 85 8f 8a 8f 87 85 86 89 81 8b 8b 82 7d 7e 79 79 7a 83 82 87 84 7b 78 74 78 6f 74 70 68 5f 64 65 60 67 63 58 60 63 6f 73 76 85 7a 69 5b 35 25 1b 02 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 25 2a 47 59 72 8b 8f 8c 74 72 6f 6f 6a 6f 6a 7b 7b 80 85 89 8b 8d 93 95 97 9e a2 98 96 99 9e 99 95 96 9e 9f a8 ad a9 a6 a5 ad ae ab a0 ac a7 ac ac b0 aa a9 a9 ac b1 af a1 a8 ae b2 b5 b3 ba b5 b2 b4 b3 ac b5 b9 b5 b9 ba c2 be b4 bd bc c5 bf bc b3 c3 c8 be c3 c4 ba bf bd bc b7 b7 c2 b1 b9 b5 ad af b4 b0 ab b0 ab a3 9e 92 77 59 24 0c 00 06 05 03 00 06 07 03 00 06 05 03 03 06 05 03 02 06 05 03 00 06 0d 0f 0e 14 0d 28 61 97 a3 a4 a0 9e a0 97 9c 96 9b 92 93 9b 95 89 8d 8b 90 8e 8b 87 95 80 84 8a 8a 86 80 86 7a 7a 7f 7e 83 7f 85 7e 83 82 75 7d 7a 78 80 85 83 8a 7b 7d 85 89 84 85 88 80 83 80 80 8c 84 88 7c 81 7d 81 80 73 7d 7d 89 81 84 80 80 7c 7a 65 74 6a 69 6f 65 62 67 66 66 65 5e 60 65 6a 7b 85 83 6e 5b 3a 26 1d 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 0e 1c 32 49 65 72 89 91 8a 77 6c 67 6f 6a 74 77 74 7a 7f 7f 87 86 91 95 92 9c 9a a1 9d 94 9c 9e 95 99 a6 9f a1 a1 a7
 a6 aa ab a9 ab a6 a5 a6 ac ae ae aa aa a9 a7 a6 a8 aa a9 b1 b1 b1 b6 b1 ae b3 ac a8 b1 a9 ab b0 b2 b7 b7 b8 af b3 b7 b1 bf b6 b9 bb b5 b8 b9 ae bd ac b7 bc b3 b6 b7 b2 b5 b9 b0 b0 ae a7 a5 a3 9e 9e a5 98 93 7b 5b 24 03 04 06 05 06 00 06 07 03 00 06 05 03 0b 06 05 03 00 06 05 09 08 06 0e 0a 0b 0b 12 25 5e 91 93 9a 95 8f 8c 94 90 94 8d 8e 92 88 8f 91 8b 93 88 8a 86 87 88 83 84 80 88 77 82 7d 7e 7d 7e 7d 81 81 85 7e 75 7c 70 7d 84 80 79 82 7d 80 76 83 77 7d 7b 81 7a 83 86 7d 8a 85 80 85 7e 74 78 72 72 73 7f 7e 80 80 84 80 81 7e 84 7b 7f 73 77 71 6d 6a 5f 65 68 67 6b 65 64 6d 75 81 81 68 55 40 37 1c 0d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 11 2a 30 46 53 71 84 87 86 77 6e 6e 64 68 69 75 70 77 82 79 7e 85 86 92 8f 8f 9b 9c 9e a5 9f 9e 98 94 9b 98 9e 9e a3 9c 9b 9f a3 a5 a5 a4 a2 99 a0 a1 ab 9e a7 b0 a7 ab aa aa b0 af ad af ae ae a6 ae aa ad ae ae ab b9 a9 a9 aa ac ad b3 b6 b2 bb b4 b2 b2 ba ac b2 b3 b1 a7 af a9 b0 a7 b4 ad a9 a8 ab a1 b1 a1 9f a0 95 95 90 84 72 60 26 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 05 09 09 14 26 55 85 89 8c 89 89 8d 8f 88 89 89 87 8a 8a 8e 86 8a 83 83 86 83 85 84 7c 80 82 7e 80 81 78 7e 7a 7f 83 76 7f 7b 83 7e 77 73 77 75 79 7a 79 81 72 72 70 7f 80 7a 7c 75 7d 82 84 86 82 7f 82 6f 71 6a 74 73 70 79 78 84 7d 75 7e 75 7a 83 85 85 8a 83 7b 73 64 5b 67 60 68 5f 67 64 6d 6f 80 76 69 60 3e 33 19 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 09 05 0f 17 1a 2d 41 5f 74 8f 8c 83 76 72 67 6a 6f 73 72 7d 71 76 74 81 81 8d 8b 93 97 9c 9d 9e a2 a0 ab a1 99 a4 9c a1 9e 9d a8 a3 9a a3 a3 a2 a6 a7 a5 ac a7 ad ac ad b0 ae b6 b2 a5 b3 ab a7 aa a9 ad a7 a2 ae aa ac a8 a8 ae a2 a8 ab b0 a8 b1 ad ae b7 a7 ac aa a3 b0 ab a6 af a8 a9 a5 a6 a4 a5 a3 a3 a7 98 9b 9d 96 94 97 90 8a 89 87 75 5f 35 06 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 0e 06 14 20 58 81 7c 8c 8d 81 88 82 87 87 87 89 82 85 82 85 82 8a 86 85 87 80 78 8b 79 7f 82 81 84 75 7b 7f 74 78 7a 7e 80 7c 80 77 78 78 7b 85 7d 78 7f 72 79 7f 84 7f 87 87 84 81 80 81 7c 79 74 76 75 70 6f 71 72 6c 6e 73 77 7f 7c 80 76 7a 7b 84 8d 90 8b 7d 74 67 62 61 6a 6b 64 6b 62 63 6d 81 7d 6d 58 3f 33 1f 16 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 14 1f 34 42 63 6f 83 90 77 6e 6d 67 74 6c 70 70 70 7d 72 73 7d 86 85 92 90 92 9d 98 9d a1 a6 ae a4 a7 a7 99 a1 a6 9c
 a6 a2 a2 a1 a4 a0 a5 a7 a3 b4 ad b2 b4 b9 b5 b6 ae b4 a9 ad a9 ab a9 a7 a9 a0 a2 a5 9f 9f a6 a9 9e a5 a4 a7 a9 a9 a5 a7 b2 a0 ad a7 a4 a8 9f a0 a6 a9 9d 9d a3 9f 9b a1 9b 98 9b 92 96 9b 95 99 8d 8f 8f 84 79 74 66 2b 0d 04 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0a 02 07 10 24 5b 7f 83 7f 7b 79 7c 81 84 86 84 7c 8c 83 88 8d 89 84 8d 81 8b 85 80 7b 7e 7a 80 7f 7a 77 76 7d 7b 79 76 79 7a 7c 7b 75 7b 79 7d 7e 73 7e 7e 72 7e 81 82 84 86 80 84 7f 7d 7d 7a 7e 7b 75 75 6d 6a 74 68 68 6a 70 81 74 70 74 76 7c 80 81 8d 8d 82 75 73 67 60 65 63 61 64 63 62 68 74 82 7d 72 5d 48 2c 27 09 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0b 14 21 32 48 52 75 81 89 70 70 71 65 6e 6a 6b 76 72 79 74 75 76 7b 88 8d 8d 92 91 94 99 96 9f 9f a5 a4 9c 9e 98 9f 98 a0 a1 a6 9f 9d a0 a7 aa b6 bd b5 b7 b9 b0 b2 b4 a9 ab a6 a2 9c a2 a3 a7 a3 9f 9e 9b 97 97 a0 9d a3 a0 9e a5 a2 a1 a4 a2 a2 a6 9e a0 9e 9f 9f a3 a0 9a 98 99 93 97 9a 9c 9b 8a 96 92 90 92 87 87 85 8b 81 88 7c 72 65 2b 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 03 0a 09 16 4d 73 7d 7d 7f 70 7c 73 7f 85 84 7e 82 7f 83 85 87 7c 7c 86 7e 7f 82 76 76 79 71 74 78 73 7a 7d 79 76 78 75 71 77 76 78 75 7a 7c 73 7d 77 7c 81 82 7a 82 79 7b 7d 7b 6e 6c 69 7e 73 74 78 6a 69 6c 68 6f 6f 6f 6f 71 65 67 6b 67 76 74 7e 93 85 85 7b 66 60 61 5e 64 6b 60 70 61 69 72 82 8a 6a 5e 4d 35 1c 0f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 14 1e 2a 42 5c 72 83 7d 70 66 68 6d 69 6d 69 74 70 74 77 77 76 7d 7c 85 85 86 90 88 93 95 9b a5 a4 a7 a5 9d 9f 9e 9c 9f 9c 9c a4 a1 ad ae b5 b5 b0 b4 ae ae af ab a5 a4 a2 a9 a9 9f 9e a1 96 a8 9b 9d 9d 9b 9b 94 9c 95 9a a2 9c a3 9f 99 9f a0 9d a1 9b 9c 95 96 99 97 8d 93 93 92 90 8e 88 8b 92 8b 8c 84 8a 8d 87 7b 83 81 7e 7e 7a 6a 35 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 10 1c 4a 6c 77 78 79 6f 78 77 78 77 78 84 86 81 7f 7e 82 7e 84 7a 77 6e 7b 7f 72 76 75 71 6e 6a 73 6d 79 79 7a 78 75 76 79 7b 6d 74 7d 79 75 84 7d 78 7f 87 76 7f 81 75 72 6b 70 7b 6f 70 6b 6a 6a 6b 6b 71 6c 62 69 6e 71 6f 65 73 63 6f 71 82 84 88 87 7c 75 68 69 5a 5d 64 6a 69 64 66 6b 85 84 71 65 45 3c 27 15 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 09 0e 1d 34 41 5b 72 83 74 75 6b 6b 6b 6c 73 6a 6a 75 75 75 74 78 7f 82 85 80 88 8a 87 8c 8f 95 98 9c a6 a3 a8 9a 9e a2
 9f 9f a1 a5 ae a3 b5 b1 b3 ad ab a8 a4 ad 99 a1 9f 9e a6 99 9b a2 a3 95 9b 99 96 94 98 a0 95 9d 99 97 96 a0 9a 9b a1 9f 9d 97 9d 93 94 92 94 91 95 86 91 8b 8a 91 8b 94 90 8c 8b 89 7a 7f 86 86 7e 86 87 77 7c 77 6e 34 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 03 06 0a 15 3b 68 7c 77 76 6d 77 7a 76 7c 7d 7f 84 7e 78 85 83 7c 7a 72 75 73 75 77 76 73 71 75 6c 76 74 74 76 7a 79 78 7a 79 77 78 7a 79 81 83 89 85 8b 7f 78 81 75 7b 73 6a 6d 6c 78 76 77 75 70 71 6d 6c 65 6b 70 5f 72 68 69 6a 6a 5f 69 68 77 79 84 88 87 72 63 60 63 63 63 64 60 6a 5d 64 69 7c 83 77 62 55 42 2f 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0d 18 2a 3c 54 70 74 73 6f 63 66 67 66 69 6b 6a 6a 6c 67 62 6a 75 7c 87 82 81 80 80 82 85 89 8f 8e 9f 9d 95 a1 9c 9e a0 a0 a9 a5 a3 ad ad ab b2 a0 a5 a0 9a 95 92 9e 92 97 93 95 91 98 99 91 94 8f 96 94 9b 92 8c 92 97 95 95 91 9a 8c 88 96 93 91 99 94 92 87 8e 8e 86 86 85 87 7e 8a 82 7b 83 82 82 7c 85 86 86 84 8c 8f 86 7e 74 6f 61 30 0c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 09 0d 3e 74 77 74 73 6f 74 73 72 74 79 72 7e 7b 77 78 6f 75 75 73 6f 6b 72 71 6f 73 74 74 72 75 68 6f 79 7a 78 70 76 78 70 71 7e 76 7e 7e 7d 79 82 73 74 77 71 70 6f 72 6f 6d 67 77 6c 71 72 6a 69 67 6c 69 5f 68 67 70 6e 5f 69 5c 6a 6b 70 83 7d 7c 78 6e 69 65 65 6a 6a 68 62 5f 67 65 6e 7b 84 78 65 54 3b 2c 15 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 12 21 2b 42 55 72 7f 74 71 66 68 6a 6b 6d 69 69 6a 65 74 68 6a 70 72 77 78 84 80 7e 83 8a 8a 8e 8c 95 96 9a 9f 9f 9a 9e a1 a3 a2 af ac a3 a0 9f 99 9b 94 91 93 8a 92 8e 90 92 91 90 92 9a 97 90 8d 91 95 8a 8b 90 99 95 93 94 93 8f 90 8a 98 92 8f 87 8d 85 87 89 84 8a 7d 80 84 84 81 7c 84 7f 81 84 84 83 82 87 84 8d 8d 7e 7f 71 6d 69 3d 0d 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 0a 04 06 07 12 3b 68 73 71 74 6a 73 68 77 74 74 74 71 72 7b 6d 71 6a 6d 69 6b 69 6a 6e 6e 73 75 6e 73 6e 67 6e 6f 73 7b 72 73 7e 78 7b 7b 81 84 87 78 79 7f 73 6d 72 6e 73 6f 68 6b 5f 6c 66 70 6d 6c 73 6b 65 67 67 66 67 63 62 65 64 65 66 66 74 75 7b 79 76 6e 66 64 68 70 66 6b 62 5e 65 65 67 64 80 7f 70 6b 50 46 2c 1c 0e 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 0a 16 15 22 49 58 66 7d 77 65 70 65 68 6a 6e 67 6a 6b 65 66 6d 6d 73 77 76 72 7f 7b 7c 76 85 85 86 89 8b 94 94 91 9b 9e
 9c a2 a2 a2 a9 9f 9f a4 93 96 94 8c 8e 91 95 94 90 8a 93 91 91 8c 89 8f 8d 8c 94 8c 84 90 88 91 90 87 8d 8d 87 8a 88 89 88 88 84 87 89 83 7c 7d 7f 81 82 7e 7d 7a 7e 75 7d 7e 7f 84 80 8e 8b 90 95 89 82 76 73 6b 60 38 0d 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 06 15 3a 5c 6c 66 69 62 73 64 71 72 68 76 71 72 6a 71 6e 67 6d 66 60 66 6b 64 69 69 6b 6a 74 75 6b 66 71 75 83 76 76 74 79 78 7b 84 7e 86 75 74 73 69 74 68 67 68 6d 6e 66 64 6e 69 6c 6b 6e 6a 71 62 69 6a 6e 66 69 63 67 5e 66 6a 68 67 6b 76 7e 72 69 66 68 71 6e 6b 6a 71 65 6a 5c 5e 63 75 8f 7a 6d 52 4a 37 22 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0b 12 1b 26 42 56 61 76 6f 70 6b 6a 64 69 66 65 6a 67 62 67 68 68 6f 77 77 6f 76 7a 7b 80 84 84 78 77 86 84 8d 93 92 91 9d 97 a6 98 a0 9b 9e 93 88 8d 85 85 8e 8b 8b 8e 88 86 92 8e 91 8a 90 85 8a 8f 93 87 8c 88 8b 96 8e 90 83 91 8a 85 81 83 83 85 7e 83 79 82 80 84 7f 7b 80 81 7a 74 7c 7c 78 7b 7b 82 84 8f 85 84 90 83 76 74 65 67 5a 3a 08 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 10 29 61 5f 62 6b 60 6e 69 60 65 6c 6e 76 6d 6f 65 67 6d 64 61 62 5e 66 61 6d 68 6b 70 74 72 6f 70 6e 6c 73 7b 71 79 79 74 79 81 76 75 74 74 75 6b 6e 71 6c 67 6b 69 64 6b 66 66 6c 6c 71 70 69 68 65 66 5e 62 63 62 69 60 60 5b 64 60 6a 74 6a 67 67 64 68 69 6a 69 71 6b 63 65 64 62 61 75 83 7e 6f 5b 49 33 21 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 26 2f 41 4e 61 71 6c 63 60 6d 60 65 6a 66 6a 6f 62 67 5e 64 68 6c 71 73 72 71 74 74 7e 7b 7e 82 78 84 86 8a 8d 92 91 96 9a 94 9b a1 95 94 8d 8e 86 82 8b 8b 8a 8c 83 8e 85 8d 83 8e 90 8e 93 8f 83 87 86 8b 85 82 8a 8e 85 81 7a 7c 84 7a 85 84 7e 79 7b 7a 7b 7e 82 7f 7a 73 78 79 79 79 77 76 7d 84 87 7e 8a 8a 80 77 73 6e 68 67 5f 3e 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 2b 5d 6a 62 60 5e 64 62 61 60 65 64 69 76 73 5b 65 66 60 62 5d 5d 5a 63 5d 66 6c 71 73 76 70 73 6f 72 72 73 7b 78 77 75 7c 7f 7a 78 74 6e 67 65 6c 67 66 63 5f 66 6c 65 68 69 6a 65 6a 66 71 65 69 6f 69 61 5c 58 64 64 6a 61 61 62 6a 6a 68 66 5e 6a 69 69 60 67 68 69 6a 63 65 58 64 72 80 7e 6f 65 46 3b 1c 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 21 32 42 56 6f 79 6b 60 6a 68 69 6f 65 71 64 6a 6a 68 6d 6c 6d 6b 70 75 75 77 70 74 73 79 7e 81 83 88 87 89 89 89
 95 94 92 9d 8d 90 97 8b 8b 87 84 85 85 89 85 87 8c 86 8b 88 88 87 93 8c 8e 85 85 84 8e 83 84 84 89 84 85 8b 88 7b 7b 76 80 78 7b 74 75 79 72 75 80 74 7c 78 7c 70 7d 82 72 73 7b 85 84 84 79 80 74 72 6b 60 66 62 60 3c 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0d 28 56 65 63 69 60 65 60 69 67 64 68 5a 65 66 70 60 6a 60 65 61 5a 62 67 65 68 76 6d 79 7d 72 6e 6e 73 6c 73 70 74 71 79 78 78 75 70 74 76 71 6f 63 65 60 67 63 5b 6a 65 68 5c 65 69 6d 6f 6d 66 6f 69 61 62 65 68 6a 5e 63 64 63 73 64 6c 68 61 6a 6c 64 69 60 60 66 6e 6d 6e 5e 5c 66 76 7d 7b 72 60 46 3d 27 14 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0d 15 19 37 39 55 6d 6b 67 69 69 65 6c 66 66 6c 6a 64 67 6c 5f 6a 6d 72 6e 72 72 78 75 80 75 7b 77 71 7e 80 80 84 82 87 8f 91 95 91 8c 8d 87 8b 87 89 8b 85 7f 88 81 84 8e 87 8a 82 87 83 86 80 8b 86 82 88 7b 81 85 85 85 81 7d 7a 7d 73 7b 7c 7c 7a 75 74 75 71 74 75 77 71 74 74 74 79 77 7d 77 7e 85 84 72 70 70 74 6e 6e 6b 61 67 5f 66 3c 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 03 27 4b 62 5f 6c 61 66 64 66 60 59 61 64 61 67 62 63 62 61 60 56 5b 5e 5d 61 5d 70 6a 75 75 6e 74 75 73 76 6e 75 74 73 6c 70 73 70 70 69 6d 6b 69 62 66 61 58 5e 5f 69 5c 60 5e 64 60 62 69 68 64 66 66 66 66 64 5e 62 60 5a 65 64 6b 5d 5d 67 58 5f 67 62 60 5f 60 63 5c 5f 61 62 62 5e 6f 75 79 75 64 4b 3f 22 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1b 20 28 3b 55 61 69 6d 66 69 63 5f 6c 6a 6a 6c 68 71 5f 69 6e 6d 6e 6f 71 71 70 6e 75 76 7b 79 7d 81 81 78 85 85 88 8b 86 90 8b 88 84 7b 86 86 82 79 84 7e 7f 84 81 87 82 83 87 82 87 84 8b 8b 8a 7c 85 80 7e 85 84 7b 7e 79 81 7a 79 70 74 78 6c 76 71 6a 75 70 76 6e 70 72 76 7a 78 72 82 7a 81 7b 7f 76 75 79 68 6e 66 59 68 57 5d 5d 42 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0e 21 4d 64 60 63 5a 60 59 63 59 59 59 63 5d 62 5a 60 62 63 62 5a 5d 5f 63 62 64 66 64 68 70 6b 6d 67 6a 6f 71 6f 66 75 6d 67 6c 5c 6c 61 66 62 65 66 65 59 52 66 5d 5f 59 60 65 62 66 5e 6a 67 63 66 61 63 5e 5f 60 5a 59 65 62 61 65 62 68 60 62 5f 66 5c 64 5e 63 5e 5c 60 59 59 5b 5b 68 7d 7e 72 61 4f 39 2a 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 09 13 27 33 43 54 61 68 61 5e 6e 67 63 6b 61 6a 68 73 6f 6d 6c 69 64 6b 6b 70 75 70 7d 76 75 76 7d 74 7a 7e 79 82 7b 85
 85 84 85 8b 87 87 88 80 7b 83 85 82 83 7e 80 84 7d 77 7e 88 7e 84 8a 78 85 7f 84 7e 80 78 7c 81 7b 7c 7b 76 71 74 73 78 73 6d 71 74 6b 7c 71 75 76 6e 71 75 6f 77 75 7a 76 81 7b 71 70 6f 6a 63 5c 60 66 5c 5f 61 59 3e 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 4d 5e 69 64 59 62 60 5b 5a 58 58 5e 5c 63 56 5e 59 60 5d 5e 64 54 62 64 63 66 61 67 65 68 6e 72 71 6c 69 69 6e 69 66 66 6a 6a 6f 5c 66 68 60 62 5f 65 60 5f 63 63 5b 60 60 63 66 5f 67 61 5c 60 68 66 5f 5e 57 61 5e 61 61 62 66 60 5e 65 5a 5b 5c 5a 63 5e 5d 56 5b 51 65 5c 60 5d 6b 70 76 78 68 4a 3b 23 11 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 12 0f 24 3b 3a 56 68 6b 62 5e 5f 68 63 67 66 62 67 68 66 64 68 6b 68 74 69 69 75 70 6f 76 77 79 81 7e 80 7e 7e 7a 7d 8a 89 8d 88 82 87 87 85 79 8f 82 78 81 83 80 83 86 78 7f 83 84 80 81 85 82 84 7a 77 7c 7a 7c 7b 7b 78 78 70 77 75 74 6e 6d 73 7a 6d 74 73 70 69 72 71 6c 72 6e 73 78 72 7c 7d 74 75 6d 6f 6d 69 66 67 62 59 64 57 59 5c 3e 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 1e 49 56 5f 5d 5b 61 54 5a 59 5d 5b 62 5a 54 58 5a 53 5f 5a 5f 5e 63 5c 59 66 63 68 6a 68 6d 6a 65 68 60 66 5f 5f 66 61 67 66 5e 62 5d 67 61 53 58 62 61 60 5e 57 60 63 55 5e 65 62 65 60 62 5f 60 61 62 62 57 60 5e 5d 62 66 64 63 60 64 5d 5d 63 65 59 5c 64 5a 66 63 59 64 65 5b 5e 59 70 73 74 65 4f 3c 25 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 20 2b 36 4f 59 67 69 5c 58 57 63 61 69 5f 67 65 5d 6d 6c 69 6e 63 75 6c 6c 6b 76 7a 79 7e 7a 72 7a 7a 7f 7a 7c 83 7b 85 88 7f 85 88 7e 7a 7a 7b 7e 79 7c 7c 7f 7d 7a 78 85 7a 81 7f 82 85 80 81 7a 78 78 75 75 7a 73 78 73 72 77 66 70 70 6c 6e 6b 65 70 6c 70 6b 73 70 71 6d 70 68 6f 7b 82 88 76 72 69 6e 69 62 5a 5f 60 5b 5b 5a 60 5d 3a 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 18 44 5f 64 64 5e 5b 53 59 5b 54 56 5f 59 5e 5a 5c 63 5b 54 5e 62 61 5c 61 62 64 64 6c 6b 6d 6a 6b 68 64 67 60 5e 64 60 5d 5e 5e 67 59 62 62 59 56 5d 5d 5d 60 59 5b 5d 5d 63 65 59 5a 5f 65 61 60 62 58 58 59 59 59 55 5d 5e 5d 62 54 5c 63 60 5c 5b 58 66 58 61 68 5d 5e 5c 5e 53 5f 59 5d 72 6a 60 45 2e 27 11 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 16 17 26 36 44 5d 69 66 60 64 5e 60 59 6a 65 6f 61 65 6b 60 6a 67 69 6d 6e 6e 71 75 74 79 83 78 7b 81 7f 7b 85 7b 87 82
 82 86 7f 81 86 88 7a 84 7a 75 7e 7d 7c 7a 7b 7a 75 7e 82 75 7e 83 81 7c 77 7a 79 7a 7c 7a 77 75 72 76 72 6e 6a 6b 68 68 6a 6e 66 6c 71 6e 65 70 72 6c 6e 72 6b 77 7f 7a 78 67 71 6d 69 60 60 5e 61 5b 5a 6e 59 58 5d 3a 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 07 05 03 12 3c 56 5e 61 62 59 5b 60 5d 5e 59 5e 53 5a 53 61 5a 5e 5d 5d 5f 64 5f 61 60 64 66 6d 6b 6a 6a 67 6e 64 68 60 5a 5e 5d 5d 63 5b 64 5a 58 67 61 5a 57 59 5f 57 66 65 58 5b 5d 68 5c 60 62 5c 5d 63 63 58 5c 61 5f 5b 5b 56 5f 64 5c 67 59 63 60 5a 60 57 67 63 66 5e 5d 5d 64 56 5e 5b 63 63 62 6d 5d 3f 2e 20 0f 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0a 10 17 25 3e 4f 5f 64 62 55 58 67 61 64 61 5c 64 68 62 69 5b 61 6e 67 6e 6a 64 71 74 7a 81 7b 77 84 76 82 7f 7a 7e 85 85 81 85 82 82 83 76 75 7a 82 7b 78 7d 7b 74 79 7a 75 7d 78 84 7b 7a 7d 75 7b 72 7b 76 6f 79 74 74 76 6d 6d 71 6b 71 6a 6d 70 67 64 6d 65 70 6c 67 65 65 69 78 73 7a 81 78 6f 6c 6a 65 61 5f 59 65 5c 59 5d 60 52 51 54 45 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 12 47 59 5e 5f 5d 5b 59 62 59 5c 5b 64 58 5d 57 5d 65 5e 60 5f 5f 67 5c 67 6a 66 61 6a 66 61 6b 62 6a 64 5c 60 5f 60 64 5e 61 58 60 5c 5b 5f 56 58 5e 60 59 5d 60 5e 5f 60 61 61 5d 5b 62 63 5f 5c 56 5e 59 5f 58 5c 56 66 5a 64 5f 59 5e 61 5f 5c 5e 5d 61 62 59 5e 5d 5b 65 53 56 57 55 5d 62 61 54 42 2c 1f 0d 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 13 20 37 40 4d 61 65 63 5b 5a 59 62 5b 63 64 5a 6c 64 5d 64 61 6b 6d 6f 6c 66 73 76 75 7a 81 84 73 7e 7b 7d 73 7b 8c 84 83 87 85 7d 7a 7b 7c 71 7b 78 74 75 76 7a 7a 74 77 74 7e 79 77 7c 6f 78 79 7b 77 75 6a 64 6d 6d 70 6d 69 71 67 64 70 67 65 6a 64 64 6d 60 6b 6e 6f 6e 71 75 75 78 76 6f 63 65 65 63 62 5d 59 53 57 58 57 52 4c 50 50 3b 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 31 54 5c 5f 5e 5b 54 57 5c 64 61 5e 60 5b 54 5e 5b 5c 60 5b 5e 5e 60 65 63 69 5f 64 61 61 5d 67 5c 5c 5f 5b 56 54 56 54 53 60 52 5a 59 5f 55 5a 60 54 57 5c 55 5c 58 5b 5e 5d 5b 5b 61 56 55 5d 5a 60 64 5b 5c 5f 5c 62 5a 61 5d 63 5b 5d 56 5b 5d 60 61 65 63 59 5a 5f 5a 5d 5e 5b 55 59 57 5a 4e 3b 28 1c 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 15 1e 2c 3d 4f 60 64 61 5f 59 5d 5c 4f 5a 5b 62 66 60 62 64 64 66 65 6b 6b 6a 72 72 73 7b 7a 79 70 73 6b 7b 7a 7d 89 7b
 7e 81 7c 75 82 72 7d 79 77 84 6f 75 80 7c 7d 72 75 79 77 7a 75 70 76 6e 74 72 75 7a 70 74 6f 66 6f 6c 6c 6e 69 68 69 63 70 6b 6c 6c 6e 68 65 65 6a 74 74 74 73 69 65 68 63 5e 6b 5a 5b 58 55 57 62 5b 56 4f 5b 51 5d 3d 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 0c 33 4b 62 59 5b 58 59 5e 69 57 62 63 66 5b 60 59 5d 63 5f 65 5f 61 67 5d 5b 63 64 5b 64 63 5f 5e 5d 5e 62 5e 5d 59 5e 59 53 5b 56 59 61 5c 5d 56 5a 63 5d 58 5a 5c 5b 5c 61 55 63 5c 57 58 51 58 58 61 5d 5e 59 59 58 56 61 58 5f 5c 60 6b 5f 60 60 54 63 5d 63 5f 5f 62 5d 5e 5b 54 59 55 52 4e 41 35 27 1a 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 1a 1f 32 42 54 60 65 5a 5b 58 5b 58 5d 5f 61 57 62 5f 69 68 61 66 66 65 6b 64 63 70 79 6f 7b 75 78 6e 6e 74 73 71 7c 79 7d 81 7d 7a 73 79 70 75 7a 77 7c 78 79 77 77 74 78 7d 7e 74 72 71 6a 72 6f 6f 73 71 71 6a 6b 68 6b 6e 6d 6e 65 67 6b 6a 6c 64 73 6c 64 6a 6a 67 6f 63 76 6d 7b 6e 66 60 61 5e 5c 59 5c 5c 5b 5e 5c 60 59 54 50 52 50 2f 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 36 55 59 61 61 5a 53 5d 62 5b 5c 62 56 65 59 5f 64 59 62 63 5b 63 5e 66 5f 62 61 60 68 63 5e 61 5f 5f 5a 59 5f 58 61 5a 56 5a 5c 57 5a 5f 52 50 5d 58 57 5d 58 5a 5f 5e 5a 66 62 5d 5d 58 59 53 5c 5e 59 63 5e 58 61 68 5a 5f 5c 64 56 5b 59 60 63 5f 5d 5e 68 64 5a 5b 5b 5b 5d 55 55 47 47 46 35 2e 28 2a 0e 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 08 1a 2c 34 45 61 5e 5c 51 52 59 52 4f 5c 5b 60 63 62 5f 5d 67 5e 57 66 64 62 6c 66 67 6a 6c 69 68 68 6b 6b 72 71 67 71 79 78 74 76 78 72 77 6f 79 72 73 79 77 75 75 7a 74 78 70 6e 71 6e 74 6d 64 6b 67 65 67 63 6b 6b 6d 67 61 65 65 67 64 61 64 6c 5f 68 68 61 6a 67 6d 73 6d 69 6f 67 5f 60 5d 59 58 5c 55 57 53 53 51 51 56 56 54 50 54 51 3c 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 36 49 5e 56 51 52 4c 5c 5b 5d 5f 5f 5e 52 57 59 5c 63 5a 57 56 54 5e 60 5d 5f 5b 5a 5a 5c 58 58 5b 5b 57 50 5a 5d 55 59 5c 52 58 55 4f 5d 55 5d 5c 5c 5a 58 5b 5d 54 65 59 57 5b 55 5a 54 4e 57 54 5e 5a 5f 62 64 5e 60 59 56 5b 5c 5e 5b 5b 5f 58 54 55 5a 5d 61 57 5d 58 5a 52 55 50 48 42 3c 31 26 1e 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 10 14 1f 32 48 5d 5e 56 56 59 54 62 59 5b 60 5a 5e 6b 5f 61 5e 5a 59 62 5e 6d 69 64 65 65 69 63 6a 61 64 5d 66 64 71 73 6d
 72 76 77 74 7a 6e 77 6d 70 77 6f 72 76 72 6f 76 73 70 77 6d 78 70 6b 65 6a 6a 66 6c 64 6b 6d 6e 68 65 66 68 68 64 64 66 67 66 66 66 65 62 64 65 6c 73 6e 64 5e 60 56 56 53 56 60 56 52 59 4d 49 49 51 50 4d 5e 4b 56 3d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 09 2b 54 55 50 50 5b 52 63 5b 59 5b 57 59 5f 58 50 58 50 5b 5f 5a 5d 5e 5b 56 5d 60 58 60 60 54 5d 5d 51 5a 5b 5b 52 58 52 56 52 55 53 58 59 58 55 56 5a 59 5a 53 5e 61 5f 57 5e 5a 60 57 50 4f 58 55 52 5d 60 60 5f 57 61 5b 5b 5b 5d 58 5c 59 5a 58 59 5c 54 60 5f 5c 5d 59 53 57 4e 4e 46 42 3b 2d 28 23 1a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 1a 1b 29 3b 54 55 65 58 5a 5c 5f 57 57 51 5c 5b 60 67 60 62 65 64 5a 5a 63 65 61 5e 64 5d 60 6f 64 60 6a 68 6d 67 6c 70 72 6a 6f 74 6d 76 74 6f 70 6d 70 76 6f 76 6e 74 75 78 71 6f 6e 64 6d 6b 68 69 68 62 68 65 5e 63 67 62 5c 67 68 62 5f 65 64 6a 6b 64 69 67 6f 64 69 6f 6d 70 63 5d 5f 56 5a 60 51 59 54 58 53 51 50 5c 53 49 54 4e 4c 4b 41 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 05 08 27 49 5c 5c 59 53 53 5c 59 54 5b 61 62 63 5b 56 58 5f 57 59 56 57 5a 5e 64 56 5b 5f 5a 5f 4f 5d 5a 5a 5d 58 5d 59 54 53 56 5a 58 57 5c 5f 56 5c 5b 60 56 57 64 59 5d 56 5c 57 5f 5f 56 57 59 5a 65 60 5d 63 68 5e 5c 5e 56 5b 5f 5a 5a 5b 5b 5d 5a 5c 5f 5f 61 64 5d 5f 5a 55 53 52 51 4e 3b 38 30 20 1e 15 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 09 17 2c 36 51 62 66 64 59 5d 5e 55 5c 57 63 5f 65 67 63 66 66 60 5a 61 5f 61 64 63 5b 5e 60 63 67 62 67 66 69 62 65 6c 67 63 75 6d 69 70 76 6b 72 77 76 6a 69 70 70 6b 6d 73 68 66 6c 6a 68 67 6b 67 63 62 64 64 66 65 5f 61 65 61 65 64 60 60 65 64 60 5d 64 68 61 6f 6a 70 69 62 4f 56 5b 52 54 57 4f 54 53 49 53 57 5a 49 4d 4f 48 5a 4c 47 39 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 03 00 25 4d 52 59 56 5b 5a 60 5d 57 5b 5d 58 5b 58 5f 5d 5a 63 5e 55 57 52 59 5d 59 5f 60 59 55 5f 5c 5e 59 54 5c 51 55 56 51 58 53 52 4c 52 5e 59 5c 5c 4d 53 56 5a 60 50 54 55 56 4e 60 4e 55 4f 53 63 66 63 60 64 60 5a 59 4e 58 55 5e 59 5a 5c 5a 5d 5b 59 58 5c 5f 5a 5a 53 56 54 56 50 4f 39 30 28 21 1e 10 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 13 25 2f 3d 54 55 60 5e 60 59 5d 5f 5b 5d 5e 60 63 66 64 63 5b 61 65 67 61 61 5f 5f 5e 66 61 66 65 65 65 69 65 66 65 60 6a
 65 64 6b 68 67 6d 6a 6e 6f 6e 6d 67 6e 72 70 74 70 62 65 6f 63 6c 67 5b 69 59 66 5b 62 61 5e 5d 65 61 61 63 57 5c 69 5f 5e 6a 68 70 64 6c 66 5e 6b 61 60 5e 5d 5c 59 51 4d 50 4d 4f 57 4d 54 54 52 51 50 4d 50 4b 50 37 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 25 48 5b 59 50 54 58 60 53 53 55 58 62 5b 5d 54 5f 5f 56 53 5a 63 57 5c 4d 5a 54 5c 58 58 60 50 55 56 59 5d 57 5a 55 55 4f 5b 52 57 58 55 58 4f 55 55 58 5f 52 5b 56 5b 56 5b 56 50 56 55 52 5a 65 66 6c 65 5c 5d 51 5a 59 58 5a 58 5e 54 60 4b 53 5f 57 50 5d 57 4b 59 5e 4c 53 52 50 47 37 3c 2c 21 18 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 0f 28 2b 49 59 62 5f 5a 61 58 61 56 5c 5f 5b 65 62 5e 62 63 65 5b 61 67 60 60 61 61 62 5f 64 66 64 64 62 68 64 61 66 66 64 66 6b 6a 64 6f 6f 76 6d 6f 6e 70 6f 6d 6e 64 67 69 74 6f 6a 63 65 62 6e 62 64 67 5e 5e 65 61 65 5d 64 66 64 63 65 64 63 65 66 70 6b 6d 6f 62 63 68 5b 58 56 58 5d 50 4f 52 55 52 50 52 4d 4d 50 4a 4e 4d 4a 4a 49 50 36 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 19 43 55 59 56 54 54 5f 5b 5b 5d 5d 5c 63 55 5a 58 58 5c 55 57 56 56 58 56 60 58 58 5b 54 5a 5d 5b 53 55 56 52 57 55 59 55 5a 5c 56 59 55 52 59 5a 50 5b 52 61 57 57 5b 54 57 4f 52 59 59 5b 56 65 68 70 70 64 5f 4e 59 56 5a 52 58 53 56 51 55 57 5a 59 5b 57 5d 5c 60 61 56 59 4f 53 48 3d 30 20 20 21 12 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 12 1a 26 30 40 54 61 6b 5f 5e 55 61 60 66 57 60 60 64 69 67 65 62 60 60 65 65 65 60 61 65 65 5f 65 63 66 6b 65 67 66 5f 61 62 60 60 67 63 64 6f 64 6b 6f 74 72 6a 6a 6c 6f 69 6c 66 6a 66 60 64 65 69 5e 56 60 5d 5b 55 5e 63 64 65 5d 64 61 6b 5a 6a 68 64 67 68 67 6a 69 67 65 5d 5e 51 51 50 50 53 4f 4c 54 4c 4d 57 4c 49 4a 4f 51 4d 4a 4e 44 37 08 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 21 47 54 51 55 54 50 55 55 58 5b 5f 63 5f 5b 55 56 5a 58 5a 59 5e 5b 5d 53 5e 54 5f 5e 50 5b 55 58 59 5a 55 55 59 54 53 56 4d 5a 57 5d 54 57 57 56 57 5d 55 55 4c 50 57 55 54 50 55 55 51 52 56 5e 6a 66 5f 5d 57 58 51 5e 56 59 58 57 5e 52 5b 5c 55 56 58 59 58 5b 5a 5a 55 54 50 4d 4a 3f 32 24 20 1c 10 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 18 15 22 32 42 54 5d 6d 5e 5d 5e 5d 64 5d 61 66 56 5b 62 60 5f 65 68 64 5b 62 5e 58 6b 5d 62 5e 62 65 64 69 66 65 6a 61 5d 61
 5d 6a 64 64 5c 65 63 5e 68 65 66 6e 6e 5f 6e 6a 65 6b 69 70 64 63 65 61 61 66 5a 56 60 5d 5a 5e 5f 5b 65 64 5e 65 64 60 69 64 6b 71 61 6d 66 66 59 50 59 5a 4a 55 55 4a 51 51 54 54 4e 52 4b 4b 4e 49 4c 4e 43 4c 4d 3b 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 1e 46 58 57 58 52 56 4b 4e 55 57 62 62 5e 5f 64 59 5d 53 5f 53 5b 4f 60 55 59 52 5d 60 57 62 59 56 5e 4b 58 5b 54 5b 4f 5b 57 56 58 5e 55 55 56 58 5b 57 59 4f 53 51 54 54 5e 4f 47 4b 52 57 60 5e 62 67 5f 5d 55 50 55 55 53 5b 5f 53 52 4f 54 55 57 54 5d 55 52 59 58 55 58 52 50 42 47 34 33 20 1b 15 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 14 19 25 2f 45 5f 64 70 64 60 62 68 5b 5e 61 5a 60 63 62 5f 68 5d 69 5e 5c 5b 5d 65 66 62 65 64 58 6b 63 5f 69 64 62 60 65 67 5f 69 62 60 64 64 6a 66 61 64 66 65 66 72 68 6a 63 67 67 64 62 60 61 5b 65 60 58 62 5f 5c 60 62 5f 67 5b 5b 59 63 62 6b 70 6c 6f 73 60 64 63 54 5a 59 59 4e 4f 4a 4d 51 54 4d 54 49 59 4e 53 4e 4f 53 51 51 50 4c 47 32 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 49 54 58 54 52 54 53 53 4c 56 55 5c 62 58 59 52 54 5a 57 55 62 56 61 5b 59 5e 5e 5b 5a 54 5c 56 55 4d 52 5a 55 53 5d 51 5e 62 58 57 5b 58 5a 5b 54 54 5a 55 55 58 55 4e 4e 50 56 51 59 54 5d 63 6b 68 5f 5d 53 51 52 57 55 57 5f 50 5d 55 52 5b 53 5a 59 53 5f 5b 61 5b 5e 5b 4f 4b 43 3b 2c 1f 1e 14 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 14 2f 35 4b 60 62 70 66 68 65 64 60 66 64 63 66 64 66 6c 6a 5d 61 60 59 67 66 62 61 5e 62 63 61 64 68 5a 5d 60 67 61 67 60 5e 60 62 64 5e 5e 62 68 65 6a 62 63 69 65 67 66 62 69 66 64 61 5e 69 56 5f 60 58 60 5c 54 61 63 5f 61 65 61 5b 62 66 68 69 63 6d 6d 70 66 62 5d 55 53 51 5c 53 56 54 58 52 4b 57 4b 48 51 5b 55 51 4b 4d 46 47 4e 4a 35 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 18 45 52 5c 54 53 4c 4f 57 4f 54 4f 59 56 61 60 5f 5c 50 55 54 57 5a 54 55 58 5c 5e 5a 53 57 52 50 52 60 56 5b 58 56 52 55 4c 5a 56 51 60 4a 58 55 53 57 55 53 52 4f 4a 53 52 50 55 58 57 5b 60 6c 64 5d 5a 58 4e 4d 5a 53 51 54 5b 55 52 52 55 5a 4e 59 5a 56 5b 58 5a 58 59 59 4d 4d 42 2f 30 1e 24 10 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0b 0a 1e 1d 2b 44 58 61 6c 71 67 5d 5b 64 5c 5a 66 5f 5f 5b 67 64 5d 64 5e 60 63 5d 64 59 5f 5f 58 62 60 64 65 60 62 66 62 63 5f
 66 5f 5c 5c 5b 5f 61 64 5e 66 5d 6a 62 60 63 66 60 5f 64 61 61 5d 64 63 67 61 56 5d 5d 5f 60 60 5e 59 53 66 63 5f 64 6a 76 5f 74 64 5d 62 58 5e 52 4f 54 50 49 53 4e 4c 55 4c 50 4f 4e 4e 46 4e 50 50 46 4a 42 4a 42 36 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 3f 53 50 4d 4b 4a 53 4e 53 52 53 55 54 56 60 59 59 59 5e 50 58 5a 5a 50 51 58 5b 56 55 55 5c 5f 58 54 4f 56 55 50 57 53 56 52 4e 52 54 50 54 57 54 50 53 55 4e 48 51 50 4b 50 4d 4e 5f 55 59 65 64 61 54 49 51 4b 52 4e 54 50 57 4d 5d 47 53 52 53 57 5d 55 5c 54 59 5a 56 50 49 4c 47 2e 22 1a 19 0f 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 12 1d 1e 2f 3f 56 64 79 70 69 63 64 5c 64 5c 66 5b 64 5d 61 66 65 59 61 61 64 64 5e 5a 55 5c 5d 5d 65 61 5f 5c 62 63 64 64 64 5e 64 55 61 63 5a 65 62 63 60 5f 64 61 60 69 65 5b 61 60 5f 5d 5c 5c 62 5c 5f 65 5f 5e 5c 54 5c 5e 5f 64 64 62 65 6a 66 70 6e 69 68 5d 65 63 5b 59 59 4e 58 56 49 52 54 4a 4c 4c 4d 44 4f 4e 54 4a 49 4c 4a 48 4e 49 3a 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 15 3f 58 59 56 50 51 54 51 46 45 4e 4d 59 5a 57 58 56 56 52 53 56 5a 5d 58 5e 52 5a 52 5e 56 54 53 58 58 56 55 4a 51 5b 53 54 57 53 58 56 4b 4e 4e 53 55 53 4c 50 52 51 4f 52 4e 4e 50 54 62 60 6a 61 5b 55 58 59 53 4f 57 55 51 4f 5b 57 4a 51 52 58 5b 57 5d 5b 52 54 58 51 4f 49 4a 3f 38 2a 1f 11 0d 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 12 1d 16 28 3d 50 5e 75 6f 6d 5c 60 63 62 63 60 5d 5b 61 57 5e 5c 58 5f 5d 5d 5f 5f 5f 5b 56 5f 5f 5f 66 63 5f 60 61 5b 5e 5c 60 60 63 58 56 5b 5b 58 57 61 5c 60 63 67 60 5c 5f 61 62 61 5e 5f 62 5d 5c 5e 60 5a 55 59 62 5f 63 5d 60 61 65 6a 72 73 72 6d 6d 67 5e 5f 57 55 59 54 55 51 4d 51 53 54 4b 4e 4d 4a 47 52 4e 4b 47 4a 4a 44 44 47 43 35 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 37 51 5e 50 4e 47 48 4b 52 4d 52 4f 54 4d 52 5a 59 52 5a 57 5b 57 5a 58 5a 52 5a 51 59 5d 58 50 57 5d 58 57 54 4f 4e 54 52 55 51 57 4d 5a 53 4e 53 50 50 51 47 51 52 51 4f 4c 4c 4e 52 55 62 64 56 53 56 55 63 51 59 4e 4f 4c 5a 59 5d 57 4d 52 4d 55 56 55 5f 59 5f 5a 55 59 48 47 42 30 20 16 14 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 06 06 1c 18 2b 40 49 62 6e 80 69 65 63 59 55 52 5a 60 60 62 5b 63 55 5f 54 5b 56 59 62 5a 5d 59 59 60 61 5c 5f 67 68 64 60 67 5e
 5c 5b 59 56 5b 53 5a 5e 5a 5b 5d 58 56 5f 5a 61 64 5f 58 60 5a 5c 62 61 64 5e 5e 53 57 5d 5d 58 5b 58 59 64 66 70 66 6f 6c 67 62 63 5a 5d 50 58 58 54 51 54 49 52 4c 4d 48 45 50 4c 53 49 4e 50 45 48 52 49 41 49 48 40 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 42 53 51 57 52 4c 4e 50 4b 4d 4f 53 53 56 4e 55 53 59 5f 5d 5d 5f 53 5a 5e 4f 5f 57 5a 5a 57 59 5c 55 55 55 57 4c 50 4d 4f 51 4f 55 4e 52 4f 53 52 4f 4f 4a 4b 51 4d 46 51 51 4e 59 53 53 57 56 55 58 56 4c 4d 4e 4e 48 4f 56 4f 51 4e 4d 50 59 4c 52 54 5f 4f 60 5f 55 56 50 4b 49 38 24 18 16 0f 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0c 0f 18 20 25 36 43 5a 6f 7c 7b 68 5f 5c 56 5c 5b 5b 5d 5b 61 59 5a 59 5f 67 5a 5f 5f 58 5e 59 58 63 5e 5e 5f 61 63 64 63 5c 61 62 5f 62 5b 5e 59 5d 62 56 5e 5a 5a 5f 60 55 5e 62 5a 67 5e 56 5b 5d 5e 62 69 59 64 5b 5b 5f 61 63 69 65 67 62 69 6d 6d 69 67 61 60 57 56 58 5b 5c 56 56 56 50 4f 4a 44 4f 4a 41 50 4a 49 4a 47 49 42 4f 54 49 45 4c 34 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 34 52 50 51 4b 46 50 4f 4b 50 54 52 58 50 59 5e 55 5e 51 55 54 59 5e 57 5b 56 58 56 57 52 54 4e 51 4e 4f 5a 58 57 5a 54 58 51 55 59 4a 4c 4d 4a 49 53 4d 50 4c 50 4f 4d 4c 4f 4c 54 4a 4d 53 59 54 5b 54 50 53 4a 50 51 53 5a 53 4f 51 52 50 59 54 5b 5b 59 54 57 57 5a 5f 53 52 49 40 24 1e 11 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 06 11 0e 1e 1f 37 42 57 6c 74 72 6e 5d 54 54 5a 5f 62 62 65 60 5f 53 62 55 61 52 59 60 63 54 56 5a 54 5d 5e 5f 5e 5b 5a 5e 5a 61 5b 60 5e 5a 5c 56 5b 54 63 59 4f 5a 59 5d 55 60 5e 5f 5c 64 5d 63 63 62 5b 5f 67 65 63 5d 5f 63 5c 5e 68 68 6f 73 6a 6c 71 61 66 5e 5b 58 5f 60 54 57 4c 51 55 56 52 50 54 54 5a 4e 4a 4f 49 4a 4b 45 46 4a 44 3b 46 34 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 35 4f 5a 4e 54 47 52 52 4f 48 50 53 4c 4f 53 5c 5c 52 5a 5a 5c 57 61 58 5c 56 5a 57 5c 52 55 5e 54 52 58 55 4b 54 53 52 52 53 54 4e 5d 57 4e 53 52 4c 50 57 48 4d 51 52 55 54 58 52 4c 4c 54 5c 55 54 54 50 47 4c 4f 52 4c 4c 5a 55 5e 56 5e 56 58 5c 5b 56 5a 57 5b 5b 5a 56 50 3e 3a 2d 1c 15 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 10 15 18 26 29 44 49 5a 76 7a 70 60 5c 53 52 5a 5d 5e 5e 57 5f 4f 4a 52 53 59 5b 4e 59 55 53 52 54 5a 5d 5b 5e 66 54 52 57 5c
 55 60 56 59 5b 5e 58 5d 5a 5b 4f 5d 54 4c 5c 59 5a 5d 5b 5e 61 58 64 62 67 5d 61 61 5a 5e 65 5e 5d 5f 62 6e 65 6c 69 65 70 59 5d 5e 60 5f 5b 60 5c 51 54 51 50 56 54 4e 51 46 4d 4b 47 4b 4f 48 48 46 4c 48 47 3d 48 35 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 4c 4e 55 4d 43 4a 4b 49 50 52 44 51 54 4e 51 4f 5c 5a 59 5e 5f 58 59 59 50 5e 54 58 57 55 56 57 53 5a 4e 50 50 52 4b 51 49 55 54 4e 50 4c 54 58 4f 50 4a 4e 40 4e 4b 4a 4d 4b 4c 5b 4e 51 5e 4f 55 51 51 4c 51 4d 59 50 4f 59 53 51 57 54 55 58 5e 57 5d 54 5a 5c 58 5a 54 47 4c 32 29 18 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 17 15 20 2a 32 47 4d 6c 7b 73 60 52 50 5a 51 5e 57 5c 53 58 5a 57 58 54 5a 5f 58 4f 55 61 57 55 5d 54 5c 5b 60 5f 5e 62 5d 5d 55 57 59 4f 56 52 57 5a 5a 55 58 55 5a 4c 57 5b 50 5a 59 58 63 5a 66 63 69 65 64 5d 60 60 5d 58 5f 62 6d 65 65 6a 69 65 67 6a 5d 59 5e 58 59 5c 52 55 55 52 4f 4d 4b 51 55 56 50 49 4d 44 4e 4d 50 4d 3e 45 44 42 3b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 2b 50 4f 49 54 46 53 51 48 4f 4e 4f 52 4d 50 56 56 5c 57 52 57 55 5f 52 58 5b 5d 53 5c 50 58 55 51 4a 56 4e 54 53 57 53 55 54 4b 4f 4a 47 49 4d 4a 50 51 4d 49 50 51 4e 54 4c 49 54 51 51 54 56 53 58 56 4f 47 50 47 4b 59 4d 54 54 50 5f 5b 55 53 55 59 56 55 52 55 5c 56 59 47 41 34 20 13 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0d 13 18 1d 26 35 3f 47 65 75 70 6f 59 54 55 58 53 5d 59 5e 57 5c 5a 5a 57 53 53 5f 5c 51 57 4c 52 59 59 5c 60 62 56 59 5b 5c 5d 62 5e 58 57 53 5d 5a 56 61 5d 56 53 57 53 4f 53 5c 58 5f 5a 62 6a 66 6e 5f 61 63 69 5f 61 61 5b 67 61 71 6d 6d 66 6d 65 6c 62 67 64 5e 61 5f 52 5d 5a 4c 50 51 52 53 4d 50 57 55 4d 51 4e 4d 4a 49 4a 4b 49 4b 46 35 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 29 50 4e 4b 4e 45 4f 51 56 48 52 55 54 51 58 61 59 5a 60 58 57 5f 5c 59 5d 59 50 5f 5c 54 58 5c 5a 52 55 55 52 51 50 4d 53 52 55 53 5b 52 4b 58 4f 53 51 4c 49 44 4f 4d 4e 53 4e 4f 56 4e 52 58 57 58 56 55 55 58 57 60 5e 4e 51 49 5d 60 61 5f 62 52 5c 5d 5c 62 54 5a 55 4d 4b 3a 2c 1e 0c 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 16 13 17 29 28 32 48 57 67 6f 63 5e 53 4f 58 50 51 5b 59 4e 5c 57 59 55 56 58 54 53 54 52 51 54 4e 4e 51 58 62 52 51 50 57
 60 62 59 55 5c 52 57 59 57 5a 4f 5a 59 52 55 54 4c 59 52 5e 54 61 63 60 62 5b 61 65 57 5c 5f 61 59 5e 5b 5f 6b 6d 5d 6b 64 6a 68 64 64 61 5a 4c 5f 52 54 59 53 52 52 55 52 51 43 44 48 49 4c 4f 50 49 48 42 46 49 42 3b 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 44 5a 55 4e 4c 50 4d 46 51 4d 51 54 52 4e 55 4c 57 59 5a 5b 5b 57 54 5c 52 5b 55 58 5a 55 54 53 53 4d 52 50 59 59 51 4d 50 4a 55 51 4e 4e 51 50 4e 4c 48 47 4a 44 4f 4f 4f 4c 4d 52 4e 4a 48 52 5d 57 5d 54 56 4f 51 56 53 53 55 5c 5d 5e 62 51 56 59 5d 5c 5f 55 57 56 58 43 37 24 17 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 08 16 1c 25 2e 35 4c 64 75 6c 5c 58 4c 56 54 51 54 4b 58 51 55 5a 54 5c 57 56 55 5e 51 54 54 50 4a 56 4e 58 58 5b 61 58 53 5c 51 5a 5a 59 57 58 5c 5d 54 52 53 52 55 56 56 51 57 57 5a 55 5b 5a 60 59 5f 5d 5d 5d 5d 5a 60 65 64 6e 6a 66 63 6d 69 6d 6b 59 5e 5e 58 5e 54 4e 50 59 53 55 4e 52 4b 57 53 4b 4b 4e 52 49 4a 4d 51 44 43 3d 47 38 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 4f 55 4d 4c 47 45 4b 4f 4b 4a 4c 4e 56 50 54 57 59 59 5b 59 5d 58 59 57 51 53 60 54 55 59 55 58 53 51 5e 55 51 50 53 51 52 4e 56 4a 4a 4d 54 4f 51 4b 4d 54 50 53 52 51 4c 4a 51 48 4a 4f 57 4a 4c 4f 56 50 50 58 51 4e 51 50 53 60 5f 62 59 56 5e 50 5a 56 58 58 55 55 48 44 2a 1e 0b 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 11 1f 2a 31 37 4b 5d 71 6e 57 57 4e 52 4b 57 51 5b 4d 54 50 50 58 52 52 59 53 50 4f 54 56 55 5f 59 54 56 4d 5a 62 54 5b 5f 5c 58 53 51 51 56 4e 5e 54 56 5d 54 5a 51 52 57 5e 5a 58 5a 57 60 5b 5c 65 5d 63 61 55 63 64 5f 65 6d 65 6b 6e 69 6e 62 63 62 61 57 5a 59 5a 59 56 4c 54 5c 5c 4f 57 58 51 54 55 55 4f 53 43 4b 4d 46 43 4f 43 36 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 27 4e 4e 54 4a 42 4b 4f 50 52 58 4b 4b 52 58 59 59 61 5f 57 5f 56 58 53 5d 5b 59 4f 58 55 51 5d 4f 51 52 4e 4d 4f 54 55 4a 4f 4d 54 4a 4d 54 4b 59 53 53 4d 4c 48 51 53 56 58 4d 4b 48 49 4b 50 4d 50 5a 56 5a 4e 52 4f 4f 56 5f 56 60 5a 5e 56 5b 59 5f 5c 58 57 51 5e 55 4b 33 2f 20 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 18 16 1c 26 2e 47 56 6b 6f 5f 54 4e 53 4a 54 51 58 55 4b 4d 56 4e 58 56 5a 59 54 53 58 57 56 57 50 4e 4d 51 54 56 59
 55 5d 57 54 5b 59 58 56 5d 50 57 50 58 5c 52 50 5c 54 55 51 58 5a 54 5c 5e 58 52 52 5f 5a 58 64 67 66 61 69 5b 67 6b 65 6f 5f 66 61 63 54 53 55 59 5b 54 5c 53 51 55 49 57 54 4b 49 4c 5a 50 4e 4e 55 4b 4c 43 46 48 3a 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 43 53 56 4f 42 52 55 45 57 50 5a 55 53 55 4f 56 52 50 55 4f 52 52 54 57 4e 56 50 5b 57 58 53 4b 4d 52 4f 52 50 50 4f 4e 51 51 4d 4e 49 49 52 52 4d 50 4a 4c 53 54 57 51 50 49 48 51 49 50 50 55 4f 55 52 47 47 4c 50 49 50 58 55 5c 5c 5e 55 55 59 5a 57 55 51 5c 55 52 40 34 24 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0e 13 20 1e 27 3a 51 5f 70 5e 59 47 48 51 54 52 5b 56 50 55 54 55 52 52 56 56 56 50 5b 55 4e 55 4c 51 55 54 5b 57 4b 52 58 52 4b 55 52 52 4f 51 55 59 4d 51 50 4d 57 54 53 51 51 55 51 5d 4c 55 51 56 55 59 5a 5b 65 63 60 68 5f 6b 69 68 63 6c 60 65 62 53 54 56 57 56 59 4c 46 51 4f 52 52 4e 54 4e 4e 46 52 54 54 4f 4a 45 44 45 49 42 36 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 47 4c 52 4e 49 53 4a 4f 49 53 4c 53 52 57 56 51 57 5f 59 5e 59 5f 55 56 51 50 55 52 4c 52 57 55 53 54 50 4c 47 55 4c 54 4d 4c 50 52 4e 4c 50 51 4a 45 46 49 51 54 50 54 4a 4d 45 4b 4a 51 47 45 4e 4f 49 4e 4b 51 56 55 59 52 59 5f 66 61 5f 56 5a 5b 55 58 58 52 55 45 37 23 1b 11 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 16 18 24 21 2f 4d 65 6f 61 59 54 49 45 4c 53 53 50 4e 4b 50 56 54 52 59 54 53 4c 49 56 52 52 53 4b 4d 55 58 54 53 58 54 53 54 54 5a 51 5c 54 58 51 52 55 55 50 4e 56 51 57 50 52 58 52 5a 52 55 54 4b 4d 5f 56 5e 5e 59 5b 66 62 60 62 55 62 65 63 60 5a 5f 51 59 57 4e 55 5a 50 51 57 4e 52 4b 57 54 4a 4f 4b 4c 4a 50 4e 53 4c 47 4b 3f 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 4a 4d 5a 56 53 51 4e 52 4a 55 53 54 55 4e 54 57 56 5d 55 51 5d 55 52 59 51 55 4f 5c 4b 5c 5b 55 58 55 51 52 49 4f 4d 54 4e 52 51 4b 4b 51 54 50 49 4f 4d 55 55 53 4e 4b 4a 45 46 4d 45 51 4b 4e 4d 52 4a 4f 50 4e 51 4a 58 59 55 66 62 5f 5c 5c 5d 56 5c 5a 4f 5d 49 48 37 23 19 0d 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 02 11 13 1b 2d 31 3c 54 69 68 62 51 4b 51 4b 53 5e 50 51 56 51 50 54 57 56 51 49 51 4d 55 5b 59 50 56 52 50 4f 50 54
 52 57 58 55 53 55 56 57 52 55 55 5b 5b 56 53 4c 5a 53 4f 57 50 51 49 4e 4e 51 4f 58 4d 51 55 59 5f 5f 55 5a 54 52 52 5a 66 5b 5e 63 5f 4f 5d 5e 5a 59 55 5b 4f 55 5c 54 4e 58 57 57 51 54 4e 51 50 57 54 46 50 4b 51 42 15 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 16 44 54 55 51 48 4e 52 53 52 54 4d 50 52 4f 59 56 58 5d 5d 5d 56 53 56 59 4a 55 5f 52 57 4e 4d 56 49 4d 55 4b 59 58 57 54 56 53 57 57 4e 46 56 54 4b 50 49 55 55 51 45 53 4e 48 51 49 48 49 48 49 4e 51 4a 4f 50 55 50 53 54 5a 58 5a 6a 59 54 53 5d 5f 5b 5b 4f 50 4d 40 38 23 12 0b 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 07 10 10 1e 2b 3b 55 6f 6b 59 4b 4f 46 4d 4a 51 49 55 4c 55 5b 55 53 52 4c 49 4e 4b 55 54 4f 40 46 51 54 4f 4e 58 53 56 50 4f 51 57 4e 4c 52 52 55 4b 58 52 61 55 4e 4e 5c 4e 56 52 4f 56 57 56 4b 55 49 50 56 58 57 59 56 55 55 5a 5e 56 5d 59 5e 53 52 5b 5e 55 52 5c 5a 4f 55 58 5c 58 52 52 55 59 51 56 50 50 51 4b 50 4f 53 48 4b 3e 17 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 3b 59 4c 4c 4c 4f 56 54 56 55 4e 52 59 50 5b 59 50 5d 5d 5c 59 56 55 57 5b 52 56 50 52 4f 56 53 52 54 55 4a 4e 50 50 52 4f 53 50 4f 54 53 4d 50 4a 4a 4e 52 53 47 43 4a 48 4d 4c 46 47 4d 48 4c 50 50 45 48 4e 53 4f 51 4b 54 5a 5d 5c 54 51 55 5a 53 55 56 4e 54 4e 38 26 18 07 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 08 0b 18 22 29 2b 57 65 6a 5e 4d 4a 49 50 4e 4d 50 4e 50 4e 52 50 4e 4f 51 51 49 4b 4f 50 53 4f 54 54 47 52 4d 51 5d 54 4f 4f 4f 54 53 50 57 58 4f 57 48 60 55 54 57 52 4f 58 4f 4b 59 50 51 51 57 54 51 56 57 57 58 58 56 51 4e 4f 55 58 5d 5b 54 52 53 57 57 4f 58 4e 57 56 58 50 54 52 4f 5e 5e 5b 5c 5e 5a 52 50 50 52 4b 49 4e 4b 3f 19 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 47 50 5a 53 50 58 51 53 5a 56 55 54 5b 55 5a 54 5e 58 53 5c 5f 59 59 58 58 5d 57 5c 5e 52 53 4d 4f 4c 4a 4a 54 50 52 55 5a 58 5b 51 5a 5c 52 50 4b 4c 48 51 4e 42 4e 4b 48 45 47 4c 45 49 47 4b 4d 4f 57 4d 4f 4f 4c 48 50 64 52 59 58 5f 5a 55 5a 57 5a 52 4f 4b 46 2e 2b 12 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 10 1c 1e 28 30 40 5f 61 60 4f 4f 49 4c 53 51 51 51 44 4c 50 5d 4e 58 55 51 4c 49 53 50 4d 4e 52 50 51 4c 45 54
 55 47 4d 4d 4d 50 46 4a 53 50 56 5b 53 51 55 4d 55 54 4f 5c 52 50 58 49 56 52 4d 54 50 5b 60 5b 5c 56 59 54 50 58 56 59 59 53 4f 51 52 4d 54 4f 52 54 55 51 5b 5e 56 5c 57 61 63 66 5c 61 5d 58 5c 59 54 48 4f 51 4e 45 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 40 5f 51 57 43 4b 51 51 52 54 5a 58 56 5a 5b 59 5a 5e 61 5b 5d 59 57 5d 58 53 4f 50 55 50 56 53 4c 50 56 52 56 4d 53 53 59 53 55 54 4a 55 51 58 4c 4f 53 4b 53 49 4e 4f 49 48 47 44 48 4c 48 49 4e 53 4e 56 50 50 48 4a 57 59 5f 5e 5a 5d 54 56 52 50 53 5b 51 4a 41 2c 1b 0c 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0d 10 1b 21 2e 3a 47 55 56 4e 4b 4e 4d 4f 54 56 54 53 4e 4e 4d 48 53 50 4d 4b 43 43 52 46 4a 4d 49 48 49 4f 50 4c 4f 4a 49 44 48 47 4c 4a 4e 45 56 52 4c 4e 53 4e 55 4f 56 4a 50 56 5e 59 53 58 54 50 4c 58 56 52 58 4c 48 52 4f 4e 54 55 4e 4d 4d 4a 54 56 4f 50 4c 51 54 56 55 5b 54 56 57 5e 66 63 67 5e 63 5e 5d 5d 53 53 4c 58 47 19 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 3d 4f 5a 5b 54 50 58 4e 58 5a 57 55 53 59 56 56 5f 59 5c 58 57 61 57 5c 59 51 52 58 4d 59 52 4b 53 4f 51 50 4e 55 56 55 55 4b 4a 56 4d 4e 4a 52 4f 4a 57 55 47 51 4b 48 48 4b 44 42 4a 4c 4d 4e 50 44 45 53 4a 50 51 53 51 54 4d 5a 56 5e 5d 57 5c 58 59 5d 4f 4d 3c 23 14 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 11 1f 1e 20 3c 3f 49 51 4b 4c 4f 55 53 50 47 4f 4e 4d 50 4d 50 4a 56 49 4d 50 4d 48 47 52 50 50 54 44 51 52 4e 4d 4b 49 47 4b 47 49 4f 4c 53 4b 4b 4f 55 4e 4c 52 53 52 50 54 56 57 53 4f 52 51 56 56 59 56 55 54 49 4c 4d 53 59 57 5b 49 4b 47 46 4c 4d 4d 47 4a 51 54 4b 5f 55 53 59 54 55 54 6b 61 6a 60 5c 5c 5e 62 56 5d 52 4b 23 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 3f 4e 55 59 49 55 57 56 4c 50 55 59 57 57 5a 51 59 5f 5b 5b 55 63 5a 59 58 57 50 53 55 54 54 4c 50 54 58 54 45 5c 56 54 56 50 4a 5a 50 4b 4f 53 4a 4b 53 4a 48 4f 44 4b 4c 4b 47 46 4e 48 4b 4a 48 4e 45 41 53 58 51 52 55 5b 5a 5a 58 56 57 57 5c 52 5c 4f 50 43 37 20 13 08 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 08 10 1a 29 2b 48 49 46 51 50 4b 49 4f 4e 50 4e 4a 4c 48 46 56 51 51 4e 43 45 4d 49 54 4d 51 50 48 52 55 54
 54 4f 4b 4d 53 4d 49 50 4f 51 4d 4b 52 57 53 5d 53 54 4e 54 57 52 50 53 57 55 4c 50 56 5d 5e 4e 4e 47 42 54 4b 58 4f 55 52 4a 4a 48 49 49 4c 48 53 4f 4e 50 53 53 4c 4f 53 50 5a 5a 4c 5f 5d 5b 62 60 68 64 5e 5e 5d 54 1f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 3b 57 57 5a 4c 52 55 54 5a 59 52 5c 60 55 58 58 58 59 55 58 5c 64 51 65 52 5f 55 5b 55 5a 58 59 56 4c 54 58 54 53 52 51 50 54 4f 4f 51 51 58 4d 55 50 4a 50 4a 4d 3d 45 54 48 48 42 4c 4c 49 44 4b 4a 51 4f 49 4f 54 49 56 5f 4f 59 5b 56 58 4d 57 59 5c 50 49 3a 31 22 10 04 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 11 17 23 2f 37 3c 44 4a 4a 47 4a 51 4e 49 45 50 51 4c 44 46 4e 50 4e 4b 49 4e 50 4a 4b 51 42 49 47 46 4d 4c 52 4c 4b 45 44 45 50 54 44 54 4c 4c 57 51 55 56 50 58 54 47 5b 57 55 4c 4e 51 4a 4a 4f 4f 47 4d 4b 4c 4e 49 53 53 4d 51 47 47 50 51 4b 4b 4b 4e 49 55 4d 4b 4f 55 50 54 4e 53 51 59 50 58 5b 5c 54 53 64 68 67 66 53 1a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 3d 4f 5a 61 51 57 56 5a 53 5c 5c 61 58 56 56 54 5b 5f 5d 64 56 5f 5a 61 60 5c 5a 53 56 56 57 56 4c 56 51 51 58 55 53 54 5f 51 54 55 4e 51 50 4b 48 4d 53 55 4b 46 44 44 49 48 42 49 45 49 47 46 4b 48 52 4e 49 4d 54 56 57 4d 58 53 4d 5a 57 53 5b 56 55 4e 43 38 27 0f 16 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 1d 25 2f 31 45 45 46 42 4c 4b 53 53 4a 4d 46 53 4b 47 4b 56 4f 50 4e 4e 51 4d 4a 4b 4d 4b 49 4b 4b 4f 4a 51 4b 44 47 4b 51 4c 45 50 40 4e 4e 50 5c 57 55 51 55 51 48 50 54 4f 4c 4f 4d 4a 46 49 4e 53 55 51 49 4a 48 4a 52 4e 4a 4c 4a 4d 50 4c 41 4e 51 46 50 4f 4f 49 4a 50 53 54 56 5b 56 5f 4e 56 4e 59 5b 62 6b 73 76 5e 28 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 38 50 59 53 50 5e 5e 55 55 50 5d 59 54 5d 51 56 55 5c 5d 5e 5c 5c 5b 6a 5a 60 58 60 56 57 55 64 5c 5a 5e 4c 57 58 57 5b 5a 59 52 55 55 51 53 53 4b 4f 48 4d 4b 4d 4d 48 4b 43 48 4d 45 4a 45 48 4d 45 4e 47 4e 4d 5a 51 54 54 59 4f 5c 5d 57 59 4c 54 4b 49 40 30 21 15 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 15 1b 2a 33 44 43 4a 49 48 4a 50 4e 44 4c 54 4f 4c 51 49 47 4d 4c 4f 4a 50 48 4c 4f 4e 47 4c 4a 4e 4d
 52 47 4a 45 50 45 3f 4b 44 4a 51 4f 4e 56 4e 47 52 51 51 50 53 50 54 47 52 50 55 46 47 4b 45 50 47 49 46 4a 44 4b 4b 45 48 44 4a 4a 4e 4d 50 4b 4c 4d 51 48 55 4c 51 52 52 53 57 52 4f 56 57 58 50 59 5b 75 77 8c 79 64 2f 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 39 5e 56 55 54 57 56 54 5a 58 5e 5e 5b 5b 5c 5c 5f 5e 5a 60 5e 5c 5d 60 60 64 61 5a 62 60 5f 5f 60 55 50 5b 56 5c 5a 54 55 54 53 54 56 59 58 50 48 4e 50 50 50 53 48 4b 55 51 4d 41 43 48 49 47 4b 48 4d 4c 52 63 52 4e 4f 57 56 5d 4f 5b 54 4e 59 4d 55 42 3c 22 1c 0e 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 10 16 24 2e 3e 44 3f 4f 4a 44 51 4e 4c 49 46 52 48 48 4c 53 4e 4d 4b 4b 50 4d 4a 4d 47 49 42 45 47 52 46 47 4a 44 47 49 41 50 48 4c 50 4e 4b 41 54 4b 4b 4a 4b 51 51 48 4c 4d 49 4d 47 48 3e 47 54 4f 4d 4b 41 43 55 4d 4f 45 48 4f 52 51 4b 47 4d 4b 50 4f 4c 50 4e 4a 51 50 4e 4e 52 4d 52 56 5a 59 54 4f 5e 67 72 71 77 64 20 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 32 56 57 57 54 5a 5b 53 5c 55 57 5f 59 59 5a 54 51 5e 5d 5c 50 63 55 63 59 5d 5a 59 54 5d 61 5b 5c 5e 5b 54 4f 5a 4d 4f 5f 51 4e 58 53 54 52 53 54 48 4d 46 4d 50 52 49 48 4e 4a 4a 43 43 44 49 4c 4f 4d 4d 50 47 55 4e 52 5a 54 52 54 54 5b 4f 4e 52 4b 45 33 22 1e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 11 21 2b 47 44 44 4e 40 4d 49 4c 47 47 4b 48 4f 55 45 4d 4a 4c 51 47 4e 4a 46 4b 4c 48 4d 4e 4f 48 4e 47 3f 47 41 43 48 44 4e 46 48 4e 49 4c 4c 4e 53 51 52 45 51 48 48 4f 4c 4a 49 42 4d 46 4a 4a 3f 4e 4e 4a 48 4f 43 43 47 49 4d 54 43 4a 48 4c 47 49 4d 49 4c 4a 54 4f 45 52 54 55 58 51 52 52 50 60 59 5e 68 66 52 29 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 32 52 53 55 5a 5a 56 57 52 61 57 5b 57 59 58 56 5a 5c 5f 5b 5c 5e 5a 57 5d 5b 56 5b 53 63 59 5a 59 57 56 56 57 4d 4f 56 59 5c 52 54 51 56 51 49 57 46 51 54 47 4f 48 4e 48 4c 45 45 46 4d 45 46 49 50 4c 53 4d 4c 4f 52 53 57 56 59 4a 50 4a 4c 50 48 4d 3b 2d 20 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 18 22 2d 42 47 46 4a 48 49 45 4c 4b 49 4d 53 4f 44 4f 4f 49 50 50 52 59 4d 4f 4e 4f 45 4b 4b 48
 44 4a 49 4f 4b 4b 47 48 48 4a 45 4a 4f 47 49 4c 52 54 4e 4f 4d 4f 55 48 56 4d 4f 4a 42 47 48 4e 4d 42 47 4b 4a 4f 49 48 50 4b 49 52 50 46 48 4a 4f 4b 4e 4b 4c 4a 56 4e 4e 4f 57 56 55 4f 4f 46 54 53 56 5a 55 58 54 50 29 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 30 4c 57 59 58 57 57 4c 5e 57 65 60 58 5f 61 59 5e 60 58 63 5e 5b 5f 5b 5c 5b 5a 5c 57 57 59 58 56 5b 59 5b 54 4b 5a 50 59 62 60 5d 55 59 55 57 4f 52 50 47 4e 51 49 52 4a 49 4d 4d 4f 49 49 51 4d 4f 4d 4f 51 56 4b 56 59 52 5b 54 4e 56 56 58 53 4b 4d 3c 25 22 0d 0b 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 20 2d 36 3e 44 4a 47 4b 4a 45 42 44 50 4a 43 49 4a 4d 51 4f 4b 4c 4e 4c 4f 4d 4f 48 4d 4d 48 49 4a 3d 47 46 49 42 43 44 42 3f 41 43 4f 48 4d 4a 4a 4c 4c 4d 4b 4c 4b 4d 4f 56 4b 3f 3b 48 49 41 45 48 45 49 47 50 49 4e 4d 49 4d 47 4c 4e 4b 4e 48 48 4b 4b 4f 4c 4b 4a 52 55 52 4b 57 50 51 4d 4e 47 4b 48 4c 45 4a 2c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2b 4c 59 5f 56 5a 5b 5b 5b 5a 57 56 57 60 56 57 62 60 5d 59 57 60 58 5f 5c 53 5a 53 52 57 56 52 53 51 53 56 58 59 53 54 5d 5f 5e 5e 5b 54 54 54 4b 51 45 47 49 4f 48 53 46 4c 4c 47 48 4a 51 52 4f 4e 4e 53 52 50 56 5d 56 57 57 5c 55 53 52 50 58 4e 40 34 1d 12 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 11 2b 31 3e 3e 40 45 4c 4b 49 4d 42 45 50 45 44 4f 4c 4f 48 4d 45 44 52 50 45 52 48 4b 47 4b 49 45 3e 44 46 47 36 46 40 53 40 41 4b 53 47 45 43 49 45 4e 50 46 4b 47 4d 4e 55 39 48 43 4c 4c 40 40 42 50 44 44 46 4b 53 4d 49 4e 4c 51 44 4f 50 46 49 50 43 50 49 4c 50 4d 4f 52 51 4b 52 50 4d 4c 47 47 44 43 51 4a 23 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 23 4a 58 57 48 59 51 50 5b 5c 57 59 50 54 5a 59 5f 59 5f 63 5d 56 51 5b 54 5b 60 5b 5c 5a 5c 54 61 51 56 59 54 56 55 58 5b 60 69 66 51 4d 4c 44 4f 43 50 4c 48 4f 53 4e 46 45 40 49 45 4c 4e 4a 50 4f 50 53 4b 4f 51 4d 56 5a 57 5f 4d 52 52 4f 52 44 42 35 16 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1c 1d 2b 38 46 42 48 4a 4b 4a 48 45 50 51 4b 48 4e 48 4f 51 4d 51 4e 4d 4c 4d 4e 40 41 41 4b
 45 49 47 45 45 47 44 51 43 43 4c 49 41 47 49 4d 4b 4e 45 55 4e 51 4a 43 4e 4b 48 4c 49 49 4b 4b 4a 46 3d 48 3f 47 4e 49 4c 48 4b 4d 46 4e 49 4d 4a 4d 51 52 49 56 4d 4a 4c 48 55 4d 53 48 4f 4a 4b 49 4f 47 52 4c 4b 50 2e 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2d 56 50 54 4e 56 56 4f 54 56 56 5d 55 56 57 5a 5d 5a 54 5f 59 60 56 59 59 59 57 5e 59 5a 5b 58 57 54 52 56 53 52 54 5c 59 5f 64 64 5a 55 54 48 4a 41 4f 47 44 47 46 4f 50 4d 50 4d 4b 4b 4f 4a 4d 56 55 55 4f 51 53 57 50 56 59 57 54 56 4b 4f 51 42 34 29 16 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 13 12 26 37 3d 3d 46 51 4d 46 49 46 47 45 4e 50 47 4f 53 49 49 49 50 4d 55 48 4a 46 44 4b 44 46 4e 49 44 44 3d 3e 4c 43 49 44 49 44 48 4d 46 4f 49 47 48 46 4f 4b 4d 4d 46 44 4f 4d 49 4d 46 4a 4a 46 4a 4b 42 44 47 50 4b 4d 4f 42 4b 48 47 50 4c 4d 4f 41 4f 4f 52 42 4d 52 4c 52 4b 4a 4c 44 4f 4d 47 46 4b 54 4e 2b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 24 45 4c 54 50 55 52 4f 4f 5a 4f 5a 59 5d 57 5a 62 5d 5a 5f 5e 5a 54 5b 5b 5f 5e 5a 59 5b 5a 54 52 55 57 58 53 52 52 54 58 5d 5d 5d 52 4d 55 4f 4c 49 4e 46 47 4c 49 47 51 49 4b 47 4c 4f 47 51 53 4f 54 50 54 51 55 55 53 5f 5a 5c 4f 4c 52 4f 45 45 35 26 08 10 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0a 19 1d 2f 3f 3e 4b 46 3f 48 44 42 4f 42 4c 3c 41 4c 45 57 4f 4f 46 49 47 46 4a 42 46 43 48 3e 4e 3f 49 3f 3b 3e 40 40 44 49 41 45 43 3c 4f 46 4b 4d 4f 44 4b 48 4d 4b 4b 40 51 40 44 45 48 42 43 4d 47 50 40 43 4a 47 49 43 42 41 46 4a 45 51 47 4c 48 47 4e 47 47 49 4c 53 50 4c 45 4a 50 4d 4e 4a 48 49 4a 55 3e 2b 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 4a 44 5b 47 4f 49 4a 53 50 54 57 57 51 58 54 55 58 53 61 5d 5d 5a 57 5f 56 59 59 5a 5a 5a 51 53 50 52 5d 56 50 57 5f 51 56 5b 5b 52 4e 4f 49 49 48 52 4b 45 48 46 4c 4a 4d 54 4f 4a 4d 59 4f 55 54 53 53 48 51 50 4f 57 54 4a 5a 47 4c 55 4e 47 3a 28 20 0f 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 14 1e 2c 3c 3c 46 4a 41 49 43 43 4b 46 51 40 4a 49 48 50 50 48 45 52 4a 43 46 45 50 49 4e
 3d 44 43 44 48 46 3b 45 4a 44 4b 45 45 49 4b 4a 4a 45 47 49 4c 4b 47 53 51 49 48 44 4b 4a 4c 40 47 4a 43 4b 3e 43 46 49 4d 43 44 3f 49 47 45 49 4e 4b 4e 4c 48 52 52 48 4a 52 4f 4c 4a 52 54 52 46 49 4b 4c 4f 4d 4b 47 2f 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 49 4d 4c 4a 50 53 51 52 52 5a 57 5b 57 52 5d 52 57 56 5a 56 59 57 60 58 58 54 54 5e 5c 52 57 56 4e 55 57 52 4b 54 56 61 5e 58 53 50 4c 55 56 4e 4a 43 4b 4a 49 49 50 4c 4a 50 46 47 51 53 49 4f 58 4a 57 55 5b 53 56 56 5b 51 57 50 50 55 48 45 38 26 1e 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 24 3a 44 40 45 43 43 46 47 45 38 3e 48 4b 48 48 40 4a 49 50 48 54 4a 4e 4d 4b 4a 41 45 48 42 43 48 42 3c 45 3f 3f 41 48 47 3f 47 4a 48 45 4e 44 46 4c 4f 4c 4b 4b 49 47 45 43 4b 47 4f 48 41 40 44 46 4c 46 49 43 4a 47 46 48 47 46 4d 45 4c 53 4b 4c 4d 4d 4b 4c 4e 55 4c 4e 4d 48 4e 45 44 45 49 42 41 47 27 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 40 49 4e 4e 4c 56 47 50 52 4b 5f 57 52 50 5c 57 56 56 56 58 5a 53 55 55 5c 55 51 5c 5b 56 58 52 55 53 5b 53 56 4d 57 58 4f 51 54 4f 44 49 4a 44 46 51 50 4c 46 47 4e 49 47 53 4d 44 46 54 51 55 4e 54 57 48 55 51 52 54 5d 56 5c 4d 50 44 41 46 27 19 0f 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0d 13 14 2d 39 46 41 3d 40 48 49 3f 4a 47 4a 41 4d 4a 43 46 4d 52 49 49 50 51 46 46 45 3f 44 40 43 44 3e 3d 47 3e 49 46 44 44 45 47 42 48 49 4a 4a 46 40 50 51 4b 54 4f 45 45 47 4a 4b 4e 4e 3c 42 48 48 3b 42 41 40 48 49 45 46 47 3b 49 4d 4b 49 49 4e 4e 4b 51 46 4f 45 4a 4c 4b 49 4a 46 4b 49 47 48 46 42 43 24 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1a 3d 45 43 49 4a 4a 4d 4f 4d 57 4b 55 56 54 53 54 53 56 50 5b 51 58 5e 5b 5f 57 5a 59 4c 59 55 4b 4f 52 4e 49 51 4e 4e 50 4f 4e 4c 4d 50 4c 41 4c 4e 4e 44 4b 52 44 56 52 4f 50 56 50 4d 50 4d 54 51 53 53 4c 52 56 56 52 54 50 4f 53 4a 4f 40 34 25 17 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 14 2e 35 40 46 3b 3e 44 40 47 43 44 4b 45 45 3d 45 46 47 4f 52 4c 4d 4e 52 48 4c 4b
 41 46 4c 39 42 3e 43 47 47 41 4a 4a 4a 46 42 46 48 47 4a 4b 45 4a 4f 44 4c 45 47 44 47 46 52 3a 24 33 4e 4a 44 3f 3c 42 45 48 43 3f 3b 40 3e 44 4e 48 4e 49 45 46 4b 46 50 4b 49 48 4e 52 44 45 4f 48 4a 49 41 4a 3b 45 2d 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 37 4e 4e 4a 45 4e 48 49 4e 4b 54 4c 53 59 56 4a 5a 5c 51 53 59 56 57 50 59 5d 54 54 56 4f 4e 55 4d 58 4e 4a 45 45 50 53 49 47 54 49 4a 4f 4d 4d 4f 4e 4b 4a 4a 4b 54 4a 4e 52 52 57 4e 51 4e 4b 4b 56 53 54 53 56 5b 50 49 54 4f 4d 4e 4a 3e 30 1f 15 0e 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0f 20 31 3a 42 47 41 46 3d 41 46 45 48 4a 42 4a 49 4d 4c 4b 4d 4f 48 4a 4c 49 4a 44 45 46 44 44 44 44 44 47 44 46 4d 44 4f 46 3d 48 49 41 4b 47 4f 52 4a 42 4f 45 43 4e 44 4b 47 45 49 4c 4d 44 3e 43 44 44 48 42 40 45 3e 42 43 3f 40 41 42 49 51 50 4c 54 4a 4e 50 4c 43 4b 49 4c 48 49 4b 4a 3f 41 44 3b 33 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 3a 44 4a 43 4b 4a 3e 4c 4b 4a 53 4f 59 57 50 53 4f 4f 4b 50 56 5a 54 58 5d 59 52 51 58 5c 55 49 51 54 51 4e 50 55 56 50 4f 4e 46 41 50 50 4d 47 4b 44 55 46 49 50 5b 48 50 53 51 57 51 56 53 4b 50 4b 5b 4b 55 47 57 50 53 5a 52 4e 4e 4b 32 28 1b 12 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 1a 27 35 47 49 42 47 44 38 42 42 46 46 4a 49 4a 44 4e 46 4c 3f 4b 4b 46 4e 44 47 43 40 40 3d 41 4b 3e 44 46 43 41 3e 48 4e 41 45 4a 49 49 44 4a 4e 47 49 4b 4f 43 49 46 42 51 47 44 3e 41 47 38 40 42 3a 47 46 44 45 3c 44 42 45 49 45 44 43 49 4a 43 4f 44 47 47 43 49 4f 3e 4a 4a 46 4b 41 3a 43 39 3c 29 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 2f 44 52 42 49 43 47 45 4c 48 51 4a 55 4e 50 50 51 53 51 4f 59 4b 56 57 56 55 53 48 51 4e 52 50 4c 54 49 4c 4a 49 46 4d 52 44 4a 3e 4b 50 4f 49 4b 4a 4c 48 48 4a 53 46 4e 49 4e 4b 57 4a 54 46 50 54 4c 50 51 4e 4f 4e 52 53 53 47 49 3d 30 22 0e 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 14 1a 30 3e 3f 47 42 3e 3a 43 3e 45 3f 46 3f 3d 47 49 50 49 4e 4a 46 48 41 4d 4a
 41 43 4d 3e 48 3e 43 42 41 48 44 43 3d 4b 4a 4a 44 46 48 52 41 45 3d 44 48 4e 43 3f 47 3e 45 48 47 3f 43 46 3e 3c 3d 3f 3c 43 4a 48 40 40 36 3f 43 48 46 48 43 4a 41 48 4a 44 48 4e 4b 47 4c 44 44 42 3b 46 46 3a 4f 3b 30 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 36 45 45 41 49 47 4b 46 49 44 46 4f 52 51 4d 51 53 53 4d 4c 4d 4b 4f 51 51 4b 51 52 54 53 4f 4e 4f 4f 4a 44 48 4a 46 42 4e 4d 4a 45 4b 46 44 49 50 46 4b 53 51 54 4b 4f 51 51 51 4a 47 50 52 4d 4f 54 53 48 53 4e 4f 51 54 53 55 50 43 3a 25 1f 10 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 11 18 24 3a 3c 45 40 41 45 3d 3a 44 3f 3f 41 3f 4c 48 4d 42 4d 4a 47 4c 46 4c 4c 4a 43 4b 44 44 40 43 4c 48 46 44 4c 45 48 46 4c 47 4f 45 49 49 46 47 47 47 3b 47 4b 46 47 48 46 48 45 4f 46 3e 48 43 4c 4e 41 45 43 40 3e 4a 3d 39 39 46 4b 4e 4e 4b 47 49 44 47 4a 3f 43 49 46 44 4a 40 46 45 42 42 44 30 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 32 3a 47 45 4b 3f 50 44 49 49 5a 4c 4b 50 50 49 4f 4b 4d 51 56 54 57 4b 54 57 50 54 4f 4e 4d 4f 50 49 48 4a 41 4b 47 46 4f 47 44 46 4d 40 4a 4e 4b 56 4a 49 50 4c 4c 44 4d 4f 4f 4d 51 53 4c 55 55 59 55 4c 55 4b 55 4f 55 4e 4d 4b 49 39 2b 1e 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 10 20 2f 37 35 42 36 41 48 40 46 40 47 3f 48 43 49 45 48 47 4d 4c 4a 4d 46 50 4d 42 41 46 43 48 48 4a 40 4b 4b 46 46 49 46 45 4d 43 51 4b 47 4a 48 45 44 4a 4d 53 40 3b 47 45 4a 47 43 43 40 41 41 43 4e 3e 3a 3f 40 48 45 45 3e 44 48 43 3f 3f 41 3d 42 44 4a 52 48 4a 3f 47 45 45 39 49 47 45 4c 43 31 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 2d 38 44 46 4e 42 44 43 43 47 4c 4c 4d 47 52 49 4a 50 53 51 54 50 4f 49 53 47 53 58 52 55 51 45 51 48 44 4b 4a 4d 4d 4c 49 46 4c 4e 47 52 4b 44 4a 49 51 43 47 43 4d 4b 4a 4d 4a 49 50 4a 4f 4d 4f 4d 57 50 51 55 4e 5b 55 4e 56 46 44 2e 23 17 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 19 26 30 40 48 3e 44 3b 3d 40 3e 40 44 43 3c 4b 43 51 44 47 4b 4a 47 44 42
 44 47 4a 3d 49 45 44 45 4b 46 47 47 40 47 47 49 58 48 42 4d 46 47 4d 45 50 41 41 44 45 45 4a 49 51 41 42 46 46 3d 41 47 46 3b 49 3a 39 44 3a 44 3f 3d 43 47 4b 43 45 43 4a 40 40 45 46 47 3f 45 44 49 47 43 3d 37 3e 3c 34 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 29 3d 4c 3e 4d 4c 48 42 46 4b 4a 53 4d 4e 4b 4a 57 4a 51 4e 4e 4e 4f 4e 4f 51 48 52 4c 43 48 49 4f 51 4c 3e 47 53 44 49 49 3e 4c 49 41 4e 44 4d 4a 4c 4e 43 4f 4b 4d 4b 4e 55 4c 49 4b 49 4d 4f 55 45 51 4d 4f 50 51 4f 53 5c 53 48 37 2e 17 0e 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0c 1f 33 34 3d 43 4a 3b 42 3e 4a 39 3c 45 3d 48 47 50 4e 4d 4b 49 4a 48 43 4a 4d 47 4d 49 4a 4b 49 44 46 48 42 44 4e 48 49 46 42 4a 4d 45 4f 51 48 48 44 47 44 4b 47 50 50 4e 45 40 42 3f 40 3e 45 43 3e 42 46 41 3f 3f 47 41 47 3f 45 40 50 43 43 3f 47 45 48 48 48 44 48 3e 3c 40 46 4b 43 42 3f 2d 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 2e 3d 45 40 40 41 42 48 4c 4c 45 4a 51 4b 4f 47 56 51 5c 48 48 52 4f 4b 51 50 53 4f 47 4e 4c 4a 4f 47 4f 43 4f 43 4b 4f 49 4b 46 50 49 45 49 4f 49 4e 46 45 4f 40 50 4b 49 57 4c 40 48 49 59 57 55 4e 4d 46 52 51 53 59 50 51 50 40 31 2b 18 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 1b 22 30 41 43 43 40 39 45 43 40 42 3d 47 46 4a 4b 48 50 4a 48 48 50 44 43 54 4a 4c 4e 4e 4a 4a 4e 49 44 4c 4d 4d 46 4f 46 40 44 44 3e 48 45 4a 45 43 4b 45 46 4f 50 58 58 4e 48 46 4b 3e 3d 3f 40 3d 49 3f 44 3e 3f 40 3e 44 46 45 40 4a 3d 46 42 40 43 45 45 43 45 47 45 44 42 3f 42 45 4c 46 38 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 23 3f 49 44 43 44 43 4a 41 47 49 48 50 4d 51 4a 53 50 54 4f 46 50 4d 4b 4a 4a 53 45 52 49 52 4b 4d 4c 48 4b 4a 3d 45 47 4a 48 49 41 3e 4e 4a 4b 4f 49 44 49 4c 4a 49 4a 44 40 4b 49 58 48 50 4d 4f 47 54 4a 46 49 51 60 51 51 50 37 24 17 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 12 1f 23 39 3d 45 45 44 38 46 3d 41 3e 4a 46 44 4b 47 4f 4d 4d 4a 44 4a
 52 4e 49 4b 49 53 4c 4c 45 43 4b 4e 3f 42 4a 53 43 49 48 4b 40 4a 47 46 48 43 44 48 47 4a 53 58 4f 4a 42 44 3f 3e 41 43 3e 3e 43 3f 3b 3c 3e 44 43 3c 42 42 3f 44 4e 43 42 43 47 4a 45 4c 39 44 3c 45 48 43 3d 48 3f 43 3d 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 24 3d 44 45 40 41 44 41 4e 41 53 3f 4b 4d 4a 4d 49 4c 49 48 50 4c 47 4c 4e 47 44 42 43 50 44 45 45 45 41 49 41 42 49 43 42 43 44 46 42 48 49 49 45 40 41 40 4e 4a 4a 53 4c 4d 50 46 46 42 49 4c 50 4d 4d 4f 4e 4b 56 56 4e 4e 3b 2e 23 10 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 14 20 2f 41 44 44 44 41 44 3c 40 45 47 45 47 45 44 4b 4b 48 4a 4b 52 49 48 4a 48 49 50 4c 48 4c 4f 49 3f 3d 4c 4e 4c 4c 42 48 52 45 41 4b 42 43 47 44 4a 45 48 4a 58 50 4a 3d 3d 43 42 40 44 42 3d 42 3e 3c 46 36 45 42 3d 3e 45 46 46 49 41 3b 45 3d 49 45 46 48 45 45 49 42 48 46 4b 49 44 37 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 3f 4b 41 3e 41 40 45 47 45 46 43 4b 45 4b 4c 4e 53 45 4a 4f 4e 52 4b 5b 42 45 48 4c 4d 4b 46 42 45 3e 42 47 49 4b 47 4c 3d 49 44 47 4f 4a 49 4e 4d 52 49 49 48 53 51 43 49 48 45 4e 48 4d 51 50 4b 56 4a 4a 53 4a 47 51 48 40 24 1e 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0d 15 2b 30 40 3f 45 3d 3b 44 44 3d 3f 45 49 3f 4a 47 46 49 45 44 50 53 56 46 4a 50 51 4c 4a 4a 4d 42 4a 4b 4d 4c 4b 4c 49 49 4e 41 4a 48 41 44 42 41 48 45 4e 50 4b 48 45 46 3e 3f 3e 40 44 41 3a 41 45 40 48 38 43 43 3e 3d 44 36 4a 40 47 3f 46 45 46 4b 42 3d 37 40 3c 41 44 45 4b 44 4b 41 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 3c 44 42 3f 48 46 40 43 3b 45 42 49 4c 49 49 48 4d 53 49 4b 51 4a 47 4f 47 49 45 4c 45 4d 3e 49 45 3f 42 40 3e 48 44 49 4c 44 48 45 4c 4b 40 47 49 49 4a 49 48 45 4d 4b 4a 47 44 53 4f 47 50 4d 43 4c 4a 4e 4b 56 4f 47 44 35 1b 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 05 15 25 30 37 43 43 42 43 3f 43 35 3a 3d 44 41 41 44 4a 4a 49 4a 45
 42 4e 46 4a 4a 4e 4c 4e 4b 52 4a 47 4a 4b 47 45 44 43 51 4e 44 47 46 3f 3d 40 39 42 3c 45 3e 42 40 3e 3d 40 3d 45 3f 45 3e 3b 3f 40 3a 3f 3f 41 3e 3a 3f 3d 42 41 3d 3e 42 43 4a 42 45 49 48 3d 41 37 49 3b 3d 45 49 43 3c 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 1c 32 46 3c 44 3f 46 43 3f 45 46 4c 4b 46 4e 4f 4b 48 48 44 4a 48 44 4a 49 3b 4a 45 44 3f 45 41 43 42 43 3f 3e 47 41 43 42 49 48 44 44 3d 54 45 41 47 4b 43 47 48 4d 52 4b 46 42 47 42 4b 4a 48 4b 47 48 40 47 4c 4c 4b 3d 35 30 16 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0d 11 29 30 42 3a 3e 44 44 41 49 3d 3f 45 44 43 4b 4c 41 45 47 3f 49 4e 46 49 4a 4e 51 46 4f 44 48 45 44 4a 4a 42 46 46 4f 4c 4a 44 44 40 42 3f 48 41 3f 42 47 3c 44 45 44 46 37 41 43 43 43 40 47 43 3a 41 47 44 4c 3d 44 44 45 41 3e 39 3f 4c 4a 49 4c 44 42 44 3d 3a 45 40 46 4c 47 47 3b 23 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 23 45 48 42 44 52 48 4a 4a 4b 47 4b 45 47 50 48 49 4b 49 47 4a 3e 45 42 41 48 3a 44 40 4b 47 3b 3f 3d 47 3a 3b 43 41 45 42 4b 4b 4e 4a 46 47 48 44 45 46 47 52 4b 4f 48 43 4d 44 44 4e 49 46 50 50 4a 4d 43 49 4f 4b 47 45 2d 27 0f 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 1e 2e 38 4d 45 49 46 3e 3c 41 3f 48 40 41 4c 44 4b 4d 42 46 45 4f 46 53 4d 4d 4d 4c 4e 54 41 47 45 49 4b 4d 4a 47 4b 45 3f 49 3f 40 45 41 48 40 3c 3a 3d 47 3f 41 4a 3d 44 3e 3e 3d 42 4c 40 47 3c 3d 45 3e 43 49 41 44 44 4b 44 44 40 3b 49 42 42 47 40 46 44 44 43 41 41 47 40 47 35 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 29 4a 4a 49 4f 47 4f 50 4f 48 43 3c 4b 42 4b 4a 4f 4f 51 47 4a 42 45 3d 47 40 42 45 41 44 3e 43 46 3c 43 41 44 4e 42 40 47 43 44 43 41 47 46 47 44 41 49 41 48 4d 48 46 43 4a 48 4b 51 4d 49 47 5a 50 4c 47 49 45 46 3f 36 23 16 0e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 13 1d 33 38 35 3b 3d 45 3c 40 39 3d 44 3e 42 3d 43 3e 3d 44 45
 4c 47 51 4b 50 51 48 49 45 40 49 4d 45 46 41 44 53 42 4e 47 46 3b 3e 45 3e 42 44 3c 39 3a 3a 3a 40 39 3d 3f 3d 3e 3f 3f 41 48 47 42 3f 3a 3d 3f 3c 3a 42 40 41 4a 3e 3e 3d 40 3a 4d 46 44 3a 40 42 44 43 41 48 42 3d 43 42 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 4d 54 57 54 4e 5a 56 4f 40 48 47 3d 48 45 4a 4f 47 47 40 47 47 40 45 45 3e 3a 3e 41 3e 44 38 35 40 40 3f 3b 45 46 48 3a 47 44 3e 45 46 43 45 4d 40 45 46 46 3d 4d 44 4f 4b 47 4f 51 4b 4e 43 4c 4e 48 45 4c 4d 49 3a 2f 14 13 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 12 1e 30 35 42 4c 45 44 3b 42 44 44 3d 42 49 44 4c 49 44 43 4b 46 50 4c 49 4c 4c 46 42 50 48 41 48 49 47 46 48 49 4b 45 3d 4a 44 45 44 3c 42 46 39 3c 47 3e 43 3c 3f 42 42 41 4d 4b 3e 3f 43 3c 45 44 40 46 40 45 47 40 46 4c 41 43 47 46 44 4a 46 46 49 40 46 42 40 3e 3d 45 4c 42 3a 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 45 45 44 51 50 51 57 50 4c 4a 4c 4d 40 4a 4a 48 4c 47 46 4b 41 46 44 48 40 40 41 48 44 3e 36 42 3d 3b 45 41 4b 48 47 49 3e 43 47 40 45 4b 46 47 48 43 49 4f 4a 50 47 45 56 56 57 52 52 54 63 59 51 4a 4c 4e 49 45 31 27 18 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0e 17 26 2e 3b 42 3d 3e 3b 3e 3e 3e 45 47 3f 41 41 45 46 45 49 4d 48 4e 48 51 48 4a 43 4c 4b 44 48 4b 42 4f 42 41 44 50 3b 3c 4a 43 45 4e 3c 48 40 3d 39 3f 49 3d 49 44 3e 3f 3f 42 45 41 44 41 3d 40 3d 49 41 44 4a 3e 47 4b 42 40 45 45 45 51 44 51 49 41 41 3f 42 3b 3e 3a 48 40 3e 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 3f 46 46 48 50 4e 54 50 4e 47 44 46 48 4a 47 44 42 47 3f 49 41 45 44 44 45 42 4a 4a 45 47 3c 3c 45 42 3c 3a 41 40 3f 43 41 3c 4d 4a 48 49 45 42 4c 4b 3c 53 4d 50 55 4f 55 60 5f 60 68 6b 6e 67 63 58 57 4d 47 38 27 1c 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 16 30 40 35 48 42 45 3e 3a 42 3c 3f 3a 39 3a 42 47 45
 4c 44 44 44 4f 4f 4a 43 47 47 46 47 45 49 4b 49 47 44 43 46 38 4b 40 44 3e 42 46 3e 3e 3d 47 40 3a 42 40 41 47 3f 3d 43 3f 43 41 47 40 3d 44 45 45 3b 43 45 40 43 44 44 44 41 44 48 45 4a 43 41 41 3e 40 44 47 40 47 3e 36 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 3a 45 42 44 50 43 46 51 45 47 4a 43 4c 44 42 45 47 46 37 3f 45 49 3b 48 40 3e 42 3d 3e 3f 3a 3a 3d 41 43 3e 41 48 41 4b 49 45 43 4b 4e 4b 4f 46 49 4f 4b 4f 59 5b 5f 5e 6b 69 6e 7a 7c 79 7a 78 7b 6a 5c 54 49 2d 23 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0e 24 33 41 40 44 3b 40 3e 3f 40 41 41 43 43 40 3d 44 49 4c 48 3d 41 47 47 49 47 44 48 3d 47 42 49 49 44 44 3c 49 3e 4b 3e 3b 3a 3a 36 3d 3b 3e 37 44 42 3f 44 40 43 42 40 42 40 34 46 39 45 46 43 42 44 42 3d 43 43 39 41 40 48 47 46 46 43 43 44 42 3f 3d 4e 4c 45 41 43 3f 3d 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1b 37 45 38 3e 40 45 48 45 44 4e 42 42 3b 43 44 44 3b 44 41 47 3f 45 40 42 40 45 42 43 40 45 3c 3a 47 42 44 3c 45 40 3f 42 44 47 43 41 49 48 51 4a 4c 57 54 54 5e 68 6d 71 80 7f 81 89 87 84 8f 88 7e 75 69 5b 4b 26 13 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 11 1e 28 31 3e 42 3d 40 41 3f 40 42 47 40 40 42 49 45 44 43 4e 4a 43 44 48 46 47 46 43 45 4a 42 42 46 4b 43 44 41 42 3f 42 3f 3b 42 3a 43 3c 3b 40 42 4a 40 40 44 42 3a 3d 3e 43 44 40 3d 48 3d 38 44 43 46 3e 43 44 43 3b 40 49 46 48 47 41 47 42 3d 42 45 3f 41 3d 44 3c 42 3f 29 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 2c 46 3c 3e 3a 3d 42 48 3f 46 3f 3c 46 47 4d 41 4b 49 40 40 3e 4a 49 47 43 3f 3e 40 42 43 3d 3b 47 44 3a 42 3d 44 48 46 4b 44 42 4d 46 55 50 56 53 5b 61 6d 79 82 89 8e 87 8c 8a 90 8c 8e 82 87 7f 79 6a 60 3d 28 11 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0b 14 25 23 34 42 3b 41 3d 3c 3f 4a 44 3e 49 42 41 48
 4b 44 49 4b 42 47 4b 44 4a 49 48 45 46 41 40 48 4d 46 41 48 44 45 3b 38 4a 40 41 3d 37 42 3e 41 42 44 3a 3f 39 3d 39 3f 43 35 34 38 38 3a 3c 44 39 43 41 3e 48 3b 46 4d 46 48 42 44 4b 49 45 43 42 49 46 46 47 3c 48 42 38 2a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 30 3e 46 42 48 45 3c 48 40 47 3c 42 42 45 48 44 4c 43 45 4a 42 44 43 4a 45 3e 44 3e 40 40 3a 3a 36 3c 44 49 3f 45 45 42 45 44 4c 4e 51 59 56 66 66 6d 75 83 84 90 8e 8c 91 87 8a 89 8c 84 84 7e 78 6d 5e 45 35 14 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 11 20 32 36 39 3a 3d 42 47 43 3b 4a 39 3b 4a 3a 47 46 41 42 49 3e 48 48 41 47 42 4a 3c 4a 49 49 41 46 4a 41 42 43 45 41 43 40 36 3f 39 3e 3f 42 3e 3c 3e 40 39 3a 39 3a 3e 36 44 3f 3d 46 3c 42 38 3b 37 3e 40 43 42 40 46 42 48 48 41 41 45 40 48 3d 44 3d 40 3f 3f 3f 33 2f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 2a 37 3e 3f 43 44 3f 42 45 41 47 46 50 45 42 45 3f 45 49 4d 3f 40 41 43 3e 3e 3e 49 3d 3a 3f 3a 47 42 3f 3a 44 49 46 48 51 52 53 4e 59 5d 64 78 82 8a 8f 90 91 9e 91 91 8c 89 8a 8c 85 83 82 83 77 6c 4c 42 19 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 16 29 31 39 39 44 42 3f 45 41 46 47 47 41 45 43 49 49 47 46 48 47 45 43 47 49 47 3e 4f 45 4c 47 40 4c 47 3d 45 43 41 48 3e 41 48 34 3e 43 3d 42 42 3d 37 38 30 41 3c 3c 3b 3d 38 33 44 41 3c 44 41 3a 44 34 41 45 3a 3f 47 4e 43 44 4a 48 45 46 49 48 47 45 3c 43 43 3b 34 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 33 40 37 44 42 3f 44 3f 50 4d 49 44 3c 3d 48 40 48 49 3f 43 3a 3f 42 46 48 40 41 3e 3e 40 3f 3c 3d 3b 3d 3f 4d 4b 50 4b 49 52 5b 61 72 75 7e 8a 90 8d 97 93 92 94 91 8d 8d 90 87 8c 85 7f 80 82 77 69 49 32 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 20 28 31 35 3e 3d 4f 3e 3d 43 40 3a 40 4c
 43 4a 39 41 3f 47 3c 46 46 42 47 44 48 4c 4a 41 42 46 3e 41 46 44 47 42 40 3e 3a 40 3e 3f 40 41 35 3f 3d 3c 33 3a 3c 37 3b 32 40 35 39 3e 39 39 3e 3b 3a 41 3e 41 41 3e 44 3e 46 40 3c 44 46 46 46 44 3d 46 43 3d 45 3f 3b 2b 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 29 44 3f 47 41 41 49 43 45 3c 46 42 3e 44 44 49 3f 3e 3d 42 3f 44 4c 39 3f 3f 48 40 3d 43 36 42 3f 39 3e 4c 45 4f 4a 4f 57 69 6b 74 82 8e 90 96 92 9a 93 8e 92 90 94 8d 8d 82 85 87 81 78 80 71 6c 5a 48 23 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 15 23 27 36 35 41 4c 42 3e 44 40 4c 45 40 4a 46 46 44 40 4b 3e 44 47 45 44 43 48 4a 43 3e 3e 3d 3c 45 44 45 45 35 41 41 3f 3e 3b 3a 3a 40 3e 3a 41 3f 37 3b 3f 3a 3b 3f 45 3d 3a 39 3e 3d 36 39 3b 42 40 44 44 3c 44 3e 42 45 48 3d 43 43 44 41 42 38 43 3a 40 45 43 30 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 2a 42 44 4a 49 42 3a 43 4a 44 48 41 3c 45 3d 4b 3e 44 3e 3e 47 44 42 47 37 3f 3e 39 35 42 43 41 3e 40 48 46 4a 4a 55 60 66 7b 83 89 92 93 99 98 9b 9b 90 8d 88 90 8e 8d 8a 84 7e 79 83 79 76 77 64 54 37 1f 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 12 19 18 2b 3a 3a 43 4a 43 48 43 47 4d 49 51 4d 45 42 41 49 47 47 44 48 44 48 47 51 48 44 49 3e 48 45 40 45 44 41 44 4b 36 41 3f 37 3f 3c 37 36 36 3f 36 33 37 3a 3b 3a 33 34 44 3a 3e 43 45 3b 3b 3b 40 43 42 3b 3f 3a 4d 47 48 41 3f 43 3d 43 42 41 3a 42 45 3d 39 2f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 2d 44 43 48 42 3a 3f 44 40 44 41 44 4c 40 44 46 3c 44 40 3f 49 3f 48 45 3d 42 48 45 4b 4a 47 3e 49 4a 4a 47 4f 56 69 75 7f 8b 94 94 a0 98 99 94 99 94 92 87 87 8a 8e 81 85 81 80 82 7e 78 7a 73 69 49 2e 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 15 19 25 35 3d 45 45 45 41 4a 50 49 58
 4e 50 3f 3f 3c 4b 43 4b 48 4f 42 4a 45 4f 51 44 49 49 42 4d 48 3e 41 41 42 3a 3e 3d 36 3e 3a 43 46 3a 40 3e 36 45 3d 3e 3e 3c 35 41 44 3f 32 37 3e 3b 40 3e 3b 3d 3d 33 45 36 3e 40 44 4a 44 40 39 42 40 43 42 3e 3c 39 3d 33 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2d 4b 44 4d 45 46 47 3f 44 48 3f 40 3e 40 44 47 44 4e 3f 4a 3f 3e 39 47 3a 37 40 3d 43 40 43 44 4d 4e 51 55 5e 72 74 85 97 6e a3 9c 94 9e 91 8f 8c 93 8a 8c 87 88 81 82 85 81 74 78 74 73 75 70 57 46 2a 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 13 1b 25 30 32 40 42 47 48 47 4d 4f 55 47 3e 44 3d 44 41 40 4b 4e 50 58 4e 4b 4f 49 50 4b 43 45 47 40 42 35 3c 3b 3f 40 36 38 3b 36 3b 38 39 41 3d 36 33 3a 3b 3d 37 3a 3d 36 36 40 41 3f 33 3e 38 3a 3b 32 3b 44 43 45 41 3b 3d 3f 3f 3b 40 43 43 39 39 38 37 32 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 2c 3b 3f 46 43 38 3e 3c 41 43 3f 40 41 45 46 42 43 3a 3d 41 41 3d 40 42 40 44 38 42 43 47 3e 45 51 4b 59 6e 74 83 94 92 9c 9e 91 92 91 8d 85 8d 84 88 8a 84 82 86 84 7e 83 84 77 76 74 6d 68 65 4d 42 1a 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0e 21 27 3d 41 3c 3f 48 47 53 52 4d 4d 4b 42 40 4d 43 4b 49 55 56 54 4e 54 4c 4e 4e 4d 42 40 3f 45 41 3c 38 3b 3d 35 3b 3d 42 37 39 39 3b 40 3a 39 3e 38 39 3b 2f 41 3f 36 35 3a 40 3b 3e 40 3e 3e 3a 42 38 3d 3d 3b 38 42 3f 40 3b 37 39 46 3a 3c 45 45 3e 2f 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 25 3f 3f 3c 45 37 47 3d 37 44 3e 41 41 40 42 3d 44 43 3e 46 3b 46 3b 45 38 3e 3e 44 41 4a 50 4f 5b 5f 6a 7f 90 90 9a 90 9a 95 8e 93 8d 95 8e 83 8b 84 84 8a 81 81 7e 76 76 75 76 6d 6a 6a 6e 5f 4d 32 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 11 1c 2b 31 3b 3a 44 4b 48 54 4f
 4f 51 4a 43 41 48 40 45 4a 56 55 5d 5a 52 4c 48 4a 45 40 44 3a 3f 41 3c 44 37 38 39 3b 43 43 42 3c 3e 3b 44 37 36 34 3d 38 34 39 3e 40 43 33 3c 3e 3e 38 44 41 39 3f 41 3c 39 47 3a 42 42 43 3b 3d 40 36 3d 35 45 3d 41 30 37 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 44 3f 3c 41 38 3c 41 3b 3f 41 41 39 3e 3d 3f 41 45 40 42 3e 44 3f 42 45 35 45 4d 4b 4b 4e 59 65 71 8d 91 97 97 94 98 92 99 91 92 8e 84 89 88 82 80 80 82 7d 7a 7f 71 71 71 6c 73 6f 69 5f 56 43 26 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 19 26 28 3b 37 3d 44 45 48 51 4a 4f 41 45 42 3c 4b 52 54 51 5d 4f 4a 4a 44 3d 3d 3e 4a 39 3d 40 31 39 36 38 32 38 32 35 3d 44 37 35 3e 36 33 39 36 3a 31 3e 36 37 3f 34 40 3d 3d 33 37 3b 3d 3b 3c 41 3c 3c 3e 3e 3d 3d 49 3d 3f 35 3f 3e 3b 3e 42 39 30 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1e 37 37 3f 41 3c 33 3e 39 3c 3b 3d 3c 38 42 3d 3b 44 45 43 41 42 41 3f 39 43 3e 43 4a 49 5e 6a 78 8c 8f 95 9e 9c 9a 90 8d 8f 8d 84 85 81 88 80 7f 7a 7b 78 6f 75 76 74 7c 75 6a 6f 61 64 64 55 34 1f 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0c 0f 25 27 34 40 33 45 45 4c 4e 50 4b 46 4d 41 45 3d 41 5e 58 57 53 4b 46 42 3e 3b 44 3d 43 30 39 39 3c 33 3f 43 3f 32 39 38 39 35 39 3f 2e 36 33 2f 32 39 34 3d 34 3e 35 41 36 38 41 3b 38 41 3f 3e 3a 36 40 3d 41 3c 3a 3e 3a 37 3e 3f 39 3c 44 39 3a 39 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 37 36 41 3a 42 36 3b 40 44 37 42 35 3e 44 3c 44 3c 42 3b 39 46 45 4d 3d 46 4d 45 54 64 6b 84 85 9c 9b 98 9a 9b 98 84 8d 84 87 84 88 80 7e 85 7d 81 7a 77 70 78 72 71 6d 70 66 61 5d 63 53 4d 35 15 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 19 1f 23 31 35 33 3f 45
 48 46 4b 44 44 46 3f 48 42 45 4e 4b 44 4c 43 40 3c 3c 40 43 3a 3e 3d 3e 34 3f 36 37 33 2f 3a 36 39 39 3d 39 37 3a 35 3c 40 3d 3e 37 3b 3f 31 3b 3c 3c 38 42 3a 3d 40 3b 3d 3a 32 3c 3b 3b 3f 44 41 36 3d 34 37 3c 3a 3b 32 31 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 38 37 45 34 40 3c 3a 3c 3d 38 3e 44 3f 48 3c 42 46 3e 45 43 41 44 49 3d 4b 53 50 66 73 83 8f 9a a3 9d 97 92 8b 8b 82 85 83 81 86 7c 7b 81 75 7c 81 78 6d 7c 75 71 6c 6d 6c 62 64 63 5b 50 43 1f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 09 1d 20 27 2a 33 3d 3e 3e 44 3c 45 45 3e 3c 38 42 3f 41 3d 41 46 43 37 3c 3d 38 38 3d 2d 3d 40 43 40 3d 41 36 38 39 38 37 41 3c 35 34 37 36 3d 3d 32 34 36 39 3a 3d 39 35 35 35 3d 3e 3c 3f 3a 34 3e 2d 3d 35 39 39 3a 3b 38 3d 39 33 35 40 2f 33 2c 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 2f 29 42 3c 34 32 38 3b 40 35 31 35 3e 43 41 3d 46 45 48 45 4c 42 43 48 4a 55 5f 7a 91 92 99 9a 9a 97 94 86 8a 8b 8a 85 7e 7e 7a 82 7a 76 78 79 7b 71 70 73 76 70 7b 69 6a 65 63 60 54 48 36 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 18 26 23 28 37 36 3d 42 3a 42 3e 44 38 44 3e 46 44 49 3c 3b 3c 39 39 39 43 30 37 37 2a 3b 38 3b 37 37 3a 3c 3b 41 38 3d 36 37 38 3e 36 3a 3c 34 39 3f 34 3a 3e 36 39 31 31 39 37 3b 38 38 3a 3b 3e 41 31 3c 33 3a 3b 34 33 38 3c 31 39 35 3c 2f 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 2d 3e 3d 39 32 31 32 3f 3a 39 36 3e 38 3b 3e 3d 40 40 49 48 50 4d 4b 54 51 68 7c 93 96 9b 9e 96 8e 8f 8f 91 8c 8e 7c 7c 7f 72 75 75 7e 70 70 7b 76 74 74 6b 6c 6b 60 67 63 62 5f 57 4a 3f 2c 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 02 11 21 22 24 35 39
 39 3e 3c 3b 3b 3a 40 40 3d 42 38 3c 3a 41 3d 38 41 3c 36 3a 3e 31 34 39 37 39 41 3b 3b 3d 36 33 38 39 3a 3e 37 39 36 35 3e 39 3a 3b 30 41 30 37 41 38 39 41 40 38 33 3c 32 3a 35 32 32 32 3b 38 42 39 3b 35 33 36 34 33 34 2f 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 14 38 40 3f 3a 33 3c 3c 40 38 38 3c 3b 3f 3e 47 3e 45 40 3e 3d 47 50 52 63 6e 7f 99 98 99 a3 91 96 92 87 8e 81 80 85 81 7b 7f 76 77 74 77 73 78 79 6d 6f 69 6a 72 6d 68 68 65 5c 5f 51 47 35 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 13 18 24 2d 36 2e 38 3e 3b 42 40 37 39 3c 3a 36 38 34 41 3a 34 3a 37 3b 39 30 37 34 36 34 3b 35 39 3e 42 3a 36 36 3c 38 33 34 33 3a 38 40 37 3a 35 36 3d 30 34 3a 36 33 3f 2f 37 41 34 37 36 36 38 2f 39 36 35 39 34 2f 38 33 30 36 37 31 2e 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 35 34 36 40 3e 3e 3b 39 27 38 36 3a 41 39 43 3e 3e 4b 50 4b 5e 5b 69 74 84 97 9b 9f 99 95 90 85 85 89 89 87 79 76 75 7d 78 74 73 77 6d 73 71 73 6c 6a 6e 67 68 68 64 57 64 53 5e 55 41 2f 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 12 19 25 28 30 3c 38 36 3c 3a 39 36 42 34 37 40 3a 37 35 37 3c 37 3c 3b 37 30 3b 3a 38 2f 35 39 38 38 37 34 37 34 34 3c 37 35 35 36 3b 34 38 39 37 3b 31 37 32 30 32 2f 35 36 36 35 3a 2f 37 3c 33 36 3a 2f 2f 30 35 35 30 39 34 2f 2e 2f 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 35 3a 41 39 3d 2e 31 30 3a 35 35 3d 3d 43 3e 3b 49 4f 4f 5a 61 67 7b 8f 8f 96 9e 97 88 8e 8b 8b 80 83 81 75 7d 7f 7a 75 71 72 73 72 71 6d 6a 6c 65 68 66 64 6a 67 64 69 5e 55 51 41 36 23 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0f 17 27
 27 31 36 32 35 3a 3b 35 3a 3c 41 42 36 3d 35 33 41 3a 3d 3b 37 3a 35 31 3c 3a 3f 3a 39 34 38 3f 41 3f 44 39 3f 38 38 3e 34 34 3d 35 3c 34 30 37 3d 3b 39 3b 36 34 31 37 2d 36 3a 38 2f 37 37 36 30 32 39 31 31 31 35 38 32 2a 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 30 2f 37 43 38 39 39 41 40 39 3b 3b 43 3e 45 4d 4f 53 5b 64 7e 83 88 8d 8f 9b 8e 8f 8c 8c 85 7f 7b 85 78 7e 79 72 67 74 75 70 72 6b 68 72 6b 67 66 65 60 6e 63 5d 61 61 5a 54 4d 40 2f 1f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 12 1a 1f 27 2e 35 33 3d 3e 3e 3c 3c 36 3d 3a 3c 38 3b 33 34 35 39 33 31 40 32 3d 37 36 33 32 3c 39 3a 3f 36 35 41 35 38 38 36 38 33 3d 37 39 39 3a 3e 37 3e 3c 34 3d 3a 3e 31 36 36 34 3c 33 3a 33 32 35 33 35 2d 34 2a 3b 35 2f 23 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 30 30 35 36 34 3c 3e 36 3c 3d 38 3b 45 36 46 51 58 65 64 7d 8c 91 98 99 8f 97 8c 8a 88 84 80 7d 84 79 69 7d 75 7b 6f 6a 71 74 65 74 66 6e 70 65 68 66 65 60 64 6a 5a 5e 59 47 40 31 15 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0b 11 1a 22 27 2a 36 37 33 2f 3d 36 3f 3b 37 36 39 40 38 35 2e 36 3b 3b 3a 33 33 30 2f 38 38 31 37 36 39 3a 3d 3e 39 33 3a 39 35 39 3b 39 3f 37 35 34 3d 35 35 31 2d 32 36 39 39 31 35 32 33 3a 35 3e 35 2f 2c 30 2f 27 31 32 29 2f 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 30 34 41 36 32 3b 3a 32 3d 3c 42 42 4a 4e 53 60 68 6f 7c 89 93 9b 98 89 93 84 8a 85 7b 85 7a 7d 71 75 72 72 6f 6f 73 76 72 62 6a 68 60 68 64 68 64 60 65 64 64 61 5d 50 4b 3e 38 29 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 10 1d 1e 29 2a 36 34 3d 36 3b 3c 3c 36 37 35 3c 38 39 38 38 38 3b 32 38 34 32 38 36 32 37 37 3b 3b 38 3d 44 39 3a 3a 33 3f 31 3e 3d 36 38 34 3a 40 3c 3a 35 36 36 36 3d 38 32 36 37 34 41 34 35 2e 29 33 32 32 33 36 2e 39 2b 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 36 30 33 3f 3b 38 3a 3d 3d 44 41 43 50 58 6e 74 7e 85 89 96 92 94 94 8a 8a 89 89 82 83 81 7d 78 74 75 71 73 6d 75 6f 72 6e 6e 6e 69 6e 64 60 67 65 5c 5f 64 5b 5b 5a 4e 4b 3c 29 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0f 1f 1f 20 30 38 38 38 43 38 37 39 32 41 37 34 3b 30 35 33 3d 3a 34 31 37 37 39 32 37 35 35 3d 3c 36 3b 3f 39 38 3c 38 36 3a 32 38 3f 3e 3d 3a 38 3b 3b 33 3a 33 35 3c 3d 31 33 38 39 2d 30 35 33 2d 2b 30 30 2e 35 2b 29 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 31 2e 30 40 38 3d 44 3d 44 3d 4b 55 62 71 7b 85 83 8a 8f 90 8e 89 8f 89 84 83 7a 7c 78 7d 74 76 75 79 77 77 6b 71 6d 6a 6f 66 63 6a 68 61 63 63 5c 59 65 57 66 56 5a 45 46 2b 1f 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 09 12 16 23 2a 32 30 39 34 34 3a 35 3e 3f 32 34 30 3c 37 37 32 28 35 36 3b 33 2b 37 30 34 36 38 39 37 33 3b 36 30 35 38 3b 38 40 3f 38 41 40 43 36 34 33 30 33 38 36 2c 32 37 39 2e 39 3c 2f 32 31 31 31 2c 2f 2c 2f 2d 24 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2b 33 3f 3c 3a 30 3c 42 46 4f 59 66 70 76 87 88 90 8c 8d 8f 90 8a 89 82 80 7a 7e 78 77 77 76 7b 78 78 6b 67 6a 6d 6f 71 70 6a 6d 63 67 6d 64 61 57 54 58 57 57 53 4f 4f 38 20 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 06 06 0d 1b 24 23 29 35 3c 3c 3a 3c 3d 38 36 34 36 3b 34 31 33 32 35 3d 33 34 30 2a 34 33 38 3b 33 38 39 3a 36 35 40 2e 35 37 39 37 3b 40 44 48 3e 40 35 3a 38 35 3e 33 31 39 35 35 3a 36 38 32 35 31 2a 30 27 2e 31 2b 2b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 33 37 3f 3f 3d 3f 41 53 55 64 6b 78 84 8c 90 8c 89 8e 8a 84 8c 89 84 7e 7e 7a 7d 78 7b 7a 6f 73 68 69 6e 6a 6e 6e 67 6e 64 69 60 62 62 69 61 61 66 57 64 57 55 4d 46 3b 27 16 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 13 14 1f 27 26 31 33 36 34 35 34 36 2e 3b 31 34 30 35 36 37 37 30 39 32 37 35 36 38 36 34 3b 3e 2d 39 36 30 30 39 3a 3d 39 4a 3f 47 40 39 3e 3c 33 3d 33 36 3b 36 38 39 3b 33 30 3c 2b 35 34 37 2c 32 36 2c 24 2b 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 28 35 37 42 3b 43 52 58 6c 73 82 8a 8f 91 8f 8c 90 8d 84 81 80 7f 85 7e 78 74 75 74 7f 72 6e 6b 6e 71 6e 70 69 67 6c 65 64 64 63 67 66 61 60 5a 54 4c 56 56 58 49 39 31 15 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 0f 17 22 2d 25 2f 33 32 3e 31 2e 36 35 38 35 3c 36 2f 3b 38 3a 32 33 34 2d 38 32 3d 31 37 3b 2f 2f 36 30 32 36 37 3d 3f 3c 40 3d 38 38 35 3a 34 38 36 35 31 3e 3c 38 3a 34 34 32 31 35 32 32 2b 2d 2e 2a 2f 1c 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 37 3e 3e 44 55 63 6e 7b 81 89 8c 8a 8f 89 87 89 84 87 7f 80 7f 7a 7a 6d 73 74 6c 74 6f 6a 66 66 69 69 67 6b 6a 64 65 65 5e 5d 63 60 61 4e 56 54 52 4e 4a 3e 39 2a 1a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 07 08 14 1b 28 23 2c 31 34 35 3c 35 34 36 3a 32 35 2f 34 39 3c 35 30 31 35 33 37 2c 30 35 3c 30 32 36 36 3c 32 38 36 33 3c 38 3d 3f 33 3c 37 31 34 39 3d 39 30 3c 41 45 36 36 33 33 37 30 32 2b 33 2c 39 31 27 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2c 30 3e 4b 52 5b 72 78 84 88 8f 8f 94 87 8c 82 81 87 85 76 7a 72 7b 73 73 71 6e 6f 71 6e 6c 6c 67 66 6d 65 64 6a 65 64 61 5d 60 5d 54 5a 55 55 4f 4d 4d 3f 42 33 20 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 10 1a 1c 22 2f 31 2d 3f 37 36 38 35 33 34 3a 36 40 36 38 31 33 36 31 38 3a 3a 37 33 35 35 36 2e 33 31 34 37 3a 38 34 32 38 39 32 37 3e 33 39 34 3c 3a 38 41 3e 41 38 35 37 34 2e 32 33 34 38 34 2f 26 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2e 37 3c 4b 5d 71 79 91 8e 81 87 90 85 88 88 80 84 83 79 78 7a 77 72 75 6a 6f 75 67 65 66 6d 62 67 6a 67 6b 6d 68 63 57 60 5e 5d 5d 55 5d 58 4e 52 49 43 39 2e 23 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 0f 18 1c 2c 26 2f 29 36 32 38 37 31 37 37 39 3f 2f 35 34 2f 30 35 33 32 30 31 37 34 2f 38 33 2b 28 36 30 34 37 39 34 30 2c 32 36 3f 35 32 3e 33 35 36 3d 3d 39 37 34 30 2e 32 32 27 37 31 2a 2f 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2f 3b 4a 5a 6a 7b 89 8d 8c 87 81 85 84 83 81 76 7e 7a 76 73 75 74 75 6b 68 64 70 6c 6b 68 68 61 6d 62 60 64 63 64 5c 5e 60 5e 5a 5a 54 54 50 4d 4d 41 37 2a 1d 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 02 06 07 11 1e 26 2d 2d 32 40 35 3b 39 33 35 3c 38 32 2f 2d 36 3b 36 34 30 31 33 3a 3b 2f 2d 32 32 32 3b 33 33 26 31 37 37 3c 3f 33 3b 34 37 3c 3c 35 35 3a 3c 3d 3c 39 35 32 3c 2b 2d 3b 2b 28 26 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 36 4a 58 75 7c 85 81 86 81 87 88 83 7c 7f 75 6e 70 7b 79 70 6f 68 74 6e 67 68 6f 6e 6a 6c 6a 6e 69 5e 5e 64 66 5b 59 68 56 4f 56 58 56 4d 4e 4e 47 39 2f 1d 07 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0a 11 12 1b 2d 2a 2d 3a 34 39 32 3b 3b 35 38 38 3e 3d 39 35 32 3a 35 39 30 39 36 35 3e 34 37 33 33 3a 3a 32 3c 32 35 39 36 38 3a 3b 39 42 47 4b 47 46 42 35 3d 36 37 35 36 31 3d 3e 2c 31 29 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 33 50 60 80 89 80 8f 84 85 84 7d 7d 7c 75 76 76 70 6f 6e 75 73 68 66 67 6f 6a 6b 6c 67 5f 62 60 56 68 64 61 61 5c 59 61 56 56 57 51 51 4a 4e 42 37 2f 1b 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0b 1b 18 2e 2c 2f 2f 31 36 30 39 47 40 44 3b 3b 37 3a 33 36 35 2c 21 38 2e 35 33 2e 35 37 39 30 39 30 36 36 39 41 39 3b 40 35 3f 3d 41 4d 4e 49 3a 3b 3f 3c 42 38 3a 31 3d 3c 2b 30 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 4c 7b 8a 80 84 81 81 86 87 7e 77 76 72 71 6d 71 75 6d 6a 71 67 6b 70 64 6d 6c 64 64 60 5c 67 5a 5f 5a 5a 57 55 50 52 5a 56 51 52 4a 42 3f 2d 25 17 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0a 1b 20 2b 37 3a 39 34 33 3d 46 4c 48 49 3c 3c 35 38 38 38 30 2a 2c 32 33 3e 31 2d 31 2e 3a 3b 38 36 40 3a 3e 3f 3e 36 3d 47 51 5a 50 50 52 48 43 42 3c 3a 33 3e 3d 31 30 26 20 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 29 61 75 7e 86 7a 79 80 75 75 7c 6d 6c 73 67 74 75 6b 6c 64 6a 61 6b 65 63 62 67 62 5f 67 5d 63 64 5f 5e 51 5d 5f 5b 5b 4e 4c 4c 4a 45 38 39 24 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 04 0d 16 26 26 34 35 38 40 43 4c 4c 48 4d 49 4b 3e 38 37 36 34 31 36 33 34 2c 36 35 34 39 3b 38 39 39 3f 40 41 3f 3d 34 40 42 50 4f 4a 54 4f 54 4d 4d 45 41 41 42 41 33 32 2c 2d 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2a 64 7d 82 7e 7d 7a 77 75 72 6d 73 6d 70 58 6d 68 68 6b 6d 64 71 65 57 67 60 69 60 5d 5f 5d 5d 5e 5a 5f 51 54 59 4d 5c 4f 45 4a 43 38 32 22 14 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 10 16 18 27 25 34 40 3d 45 42 4b 4c 4e 49 46 3e 3d 35 29 30 2f 33 38 31 2e 39 34 30 34 3b 40 44 40 41 40 3e 44 3f 3e 3e 49 48 42 55 4c 4f 58 4f 49 49 3c 45 3b 3d 32 3b 30 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2c 5f 73 7d 70 73 73 6d 6d 69 68 64 67 68 66 65 64 5b 62 69 62 62 5e 5f 60 5d 60 5e 60 5d 58 56 50 51 52 4e 52 50 4b 4f 4a 41 3e 38 25 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0b 11 1c 24 21 32 34 38 41 47 3c 43 56 46 41 38 37 34 32 2b 2e 33 30 2d 34 35 3b 30 3c 36 3e 3a 35 3c 3e 3d 3d 43 43 3d 48 4a 51 4b 55 4d 4f 53 51 52 4b 3b 40 32 34 2c 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 4e 67 6b 5b 68 69 5e 69 62 5b 5a 5d 5e 59 5f 6a 54 5e 61 5e 51 5a 52 4f 56 51 59 56 4d 4f 51 54 51 47 53 4e 4c 42 3e 44 2f 2e 20 14 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 18 1a 22 2b 2f 39 45 48 4b 3f 41 3d 3f 37 2d 2a 33 36 33 32 36 33 2e 36 35 3d 3c 38 35 37 3d 3f 40 3e 48 3f 4f 4d 47 51 50 55 4d 51 4f 54 54 4a 4c 43 3c 34 2f 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 47 53 5b 57 52 5b 5e 62 57 5f 51 55 57 5a 5b 56 53 55 53 50 54 54 51 52 50 54 52 4c 4c 4f 43 40 51 44 49 3c 41 3f 33 24 1b 1a 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 08 0d 16 18 19 2d 33 2f 3c 41 45 37 34 33 32 35 31 2b 2c 2b 32 35 36 34 2b 31 3a 37 30 39 37 43 42 48 52 55 4a 58 53 59 59 54 53 50 55 4f 47 4e 3e 43 3f 3a 37 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 2e 36 37 32 3a 3b 4d 46 48 4d 52 46 42 46 4a 4d 49 4e 44 4b 4a 48 45 40 40 46 4d 3e 3e 3e 3e 41 3d 34 35 2d 29 1f 16 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 10 14 23 1f 28 33 3d 2d 2e 33 25 29 27 27 2f 2c 2f 35 2c 30 26 2e 29 27 2c 31 39 42 4c 4a 52 4b 52 56 4a 56 5a 59 53 4e 4d 4e 45 41 42 37 35 2d 2b 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1b 1e 22 1f 22 2a 2a 2e 33 30 30 2b 40 39 33 39 35 35 2a 38 37 30 30 29 33 2f 2b 2e 2a 28 21 1e 18 17 12 13 0d 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 07 0d 10 17 28 26 22 30 28 35 2d 24 29 2b 28 27 2a 1f 22 1c 25 24 1f 20 2f 3c 3d 4b 4c 45 50 4a 4e 4c 51 55 4f 47 46 42 3f 3f 3c 36 35 2c 1f 21 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 11 0f 0d 0c 14 21 1a 25 1f 24 1b 1f 1e 17 22 1c 1e 1d 12 17 1f 17 1a 19 1c 15 16 13 10 0d 05 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0a 0f 14 11 1f 24 27 24 27 22 22 1f 19 14 15 0f 0d 0f 19 11 1b 1a 2d 38 3e 3d 34 2f 35 36 31 3e 36 30 39 33 2f 2f 2c 20 24 25 16 10 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 08 05 03 04 07 09 07 04 14 0d 08 08 0d 09 0e 0d 06 14 0a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 14 0e 10 0a 0a 11 0f 06 05 03 00 06 05 07 05 10 11 17 1d 16 20 1d 14 14 22 20 27 18 1e 20 14 20 10 11 10 12 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0b 0a 0c 08 06 06 0e 07 0a 09 13 03 09 0f 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
