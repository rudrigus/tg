 ff ff 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 08 06 09 03 0a 06 09 03 06 06 0b 09 0a 10 0c 18 13 15 1e 17 19 15 05 1c 1b 27 2e 2d 2f 2d 25 1e 20 18 1f 27 32 33 2e 53 62 60 5f 75 7e 7f 77 87 8e 93 aa 9d 97 8f ac d0 dc e9 e4 dd da c8 b6 a3 9a a2 ab bc e5 fa e6 e1 ce be ad a4 a7 b3 a5 63 32 20 1b 24 4e 52 64 6f 66 78 a9 e5 ff ff ff ea bc 8d 7f 7f 90 83 6d 5e 41 2c 1b 13 0b 0a 10 0d 06 10 15 11 11 0e 07 0b 0f 09 10 0c 05 0b 08 03 08 06 05 05 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 08 09 07 0e 0b 09 06 05 03 01 08 07 0e 10 0a 12 14 0b 0d 07 09 0e 06 14 0e 1e 11 19 21 1a 1e 1e 1d 1f 21 1e 31 2f 39 3f 48 54 3c 36 31 35 38 42 57 55 50 5f 73 70 86 94 b6 b8 c2 ed ff ff ff ff f2 f5 ef fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 e9 ed ee e5 a2 83 6f 49 44 70 87 7d 7a 78 7d 8b ba ff ff ff ff fb b9 a9 aa b8 b1 8c 7a 7a 60 44 36 22 17 13 18 18 31 35 31 34 28 14 12 11 10 1e 14 0b 0e 05 05 0e 0c 05 03 00 06 05 0a 05 0a 14 0e 01 09 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 04 06 05 03 01 06 05 08 00 06 07 03 0b 06 05 0d 01 06 0b 07 07 0c 0a 12 04 15 0b 12 12 0c 16 13 1a 1b 1f 20 1f 1d 1f 29 2b 29 2a 2a 24 2b 37 3d 2f 36 46 4c 61 60 53 5c 4b 52 60 73 81 6d 6e 74 93 cd f7 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef df be ad 8f 8e 86 82 7f 80 79 84 98 cf f8 ff ff fa d1 c0 c7 cb c2 9d 8c 9f 9f 80 6b 49 1d 23 24 3d 50 49 50 49 3b 35 34 26 1e 2a 18 16 13 11 0f 05 0a 0b 04 01 06 06 03 0c 0b 1e 1c 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 07 05 07 00 06 0b 0a 07 09 05 0d 0f 07 07 06 09 11 10 12 0a 11 0f 18 14 1e 15 10 1a 12 16 23 22 17 1c 1b 21 26 35 3e 3a 2d 3b 34 34 34 3a 50 50 58 67 65 81 92 94 8a 7b 76 66 6f 80 84 91 b5 e4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f0 ff ff ff fe eb d3 c5 b0 9e 98 8c 7f 83 85 8f 9a a9 c0 d1 df e2 ca c0 c2 cf c1 a3 91 ac c4 af 92 5d 3b 4b 5e 74 85 75 78 6c 65 57 44 44 38 43 34 3c 2d 24 1f 10 0e 09 04 0b 06 0c 05 0a 12 1c 1c 16 06 05 03 00 06 05 03 00 06 08 03 04 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 06 0b 05 0e 14 0f 0c 00 0c 05 0b 10 0f 1f 1d 13 14 0e 13 11 18 19 16 0f 1b 30 23 1f 21 22 20 3a 3b 39 4e 4e 4a 47 4e 43 48 49 58 73 a4 c5 dc e0 f2 f6 f4 ec cc 9d 9e cd f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e0 dc d3 e4 e3 e2 dd ce b6 b5 ab a9 9d 93 95 8f 92 a1 a8 b1 b2 b3 bb b5 bc a9 ac a7 98 95 9c aa b5 a3 8d 83 94 98 a1 a1 96 96 9a 93 8c 75 69 63 64 58 4b 3f 39 28 1b 14 0e 04 0d 08 0e 0a 03 07 0e 0d 04 08 0c 11 0f 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 09 06 08 08 0a 06 09 0c 11 16 13 12 0d 11 1a 12 14 19 14 12 15 1f 16 1c 22 2e 2a 2c 27 26 32 38 42 51 50 59 68 72 68 70 67 69 7a 9e ae dc ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec db d4 d3 d9 d0 e2 d0 c6 c4 bb b7 b0 a9 a5 a1 a5 a8 9f aa b0 b3 ac ac a9 9b a7 9f 91 8c 9a 94 a4 a8 ab 75 b3 b1 ae b8 b1 bb c0 c4 b9 b1 9d 9c 8f 7d 69 4b 41 38 29 26 18 1b 10 11 12 0f 0f 07 13 03 0e 06 09 13 0e 09 08 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 0a 03 06 05 07 07 06 07 06 0c 0c 05 0d 0f 15 13 12 10 11 1e 23 1b 18 20 19 20 28 2a 35 30 2c 29 2d 30 37 40 4c 5e 69 6e 83 8a 80 7d 7c 89 8b 97 ac b7 cb dc f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 e7 d6 e3 e3 e1 df db d3 d0 c7 cd c9 b7 be b4 b0 a8 a7 ae a7 ac af b2 a7 a4 9d 98 9b 97 98 95 a8 ae bd bf b4 ad bc ba bb cc da da d4 cd cc bb a6 93 74 55 54 4e 32 2e 2a 23 22 17 15 14 09 07 03 0c 06 05 11 0b 06 06 03 00 06 05 03 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 0c 07 09 06 05 09 05 06 05 0a 08 0f 09 0d 0f 0a 0f 07 10 11 13 17 1e 1b 25 15 24 20 24 28 27 27 30 35 37 4a 45 49 46 45 64 69 68 69 79 7e 7b 85 89 8b 9c a5 a7 b4 bd c4 cf e7 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed f4 f2 ed ee e8 e2 dd d6 d7 d5 d0 cb c4 c2 b8 b8 b6 b0 ad a9 ab aa ae ab a9 a5 a6 9e 99 a0 ad b1 bd c4 be c4 c9 c5 cc da de e7 e0 e0 cd b8 99 7a 6f 69 53 4f 40 3b 38 31 34 38 26 1d 1f 05 10 07 07 0a 11 16 08 04 01 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 02 06 05 08 01 06 05 09 04 06 05 09 07 0a 14 11 0e 09 05 05 14 11 14 1d 26 30 21 26 20 27 2d 2a 34 36 38 48 4f 54 59 60 60 6e 77 71 7b 7d 7d 7e 89 8b 8b a0 a8 ad b8 b8 ba c9 d4 e4 e6 f2 ff ff ff ff ff ff ff fd fb f9 eb f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fc f2 f4 ef e0 e9 e0 d8 d0 cc ca c9 c0 bc b4 b8 b3 c2 b5 ae b4 a9 a8 a9 a8 ac b4 b8 be c4 c9 c7 c8 c8 ca df de e4 e5 db d4 b8 92 8b 71 5d 52 4b 3e 3f 35 3a 45 40 3c 37 2a 19 12 0c 06 08 05 16 14 04 00 06 05 03 04 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 05 03 00 06 06 09 09 07 05 06 05 0e 10 0f 13 0a 07 14 1d 13 18 17 19 19 16 1f 1e 25 21 29 38 34 34 3d 4b 4b 51 68 6e 7d 78 80 81 81 86 88 90 89 97 97 9a 98 a4 a3 b6 c1 c4 c9 ca ce d5 df ef f4 ff ff ff ff fe f5 e5 dd e1 e5 e9 e8 f1 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f8 ec e4 e4 e3 d8 d3 ce c2 c4 bb be c3 c1 c5 b9 b7 ba b9 b5 b2 c4 bf c8 cd d7 da cf d8 da e0 eb ef e6 d9 d5 ac 9d 85 79 68 59 5e 4d 40 42 3d 47 46 41 4a 3d 2f 2f 28 23 11 11 0f 07 03 00 0b 0a 03 08 07 09 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0c 0e 0d 06 0d 13 05 10 18 19 15 15 18 16 1f 25 16 1e 26 2e 36 39 40 4e 52 59 63 75 7b 7e 8d 85 95 92 99 9e 9b 9d 9c 9b 9b a6 ac b2 b3 ba c6 bf d1 d9 dc da e8 ee f3 ff ff fe f8 f4 f3 eb e9 e1 df f2 f0 f2 e8 f0 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ef f3 f3 ef e4 de d9 ce cb c7 cf d1 d1 c9 c0 c2 c6 c1 c2 ca cb d9 db da d7 dd e2 f1 fa fb fe e1 e5 c8 b6 a0 8d 73 72 6a 5e 5a 54 47 4f 53 49 45 41 3f 49 4b 49 28 12 15 09 05 0d 0e 0d 0e 06 07 0e 05 06 06 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 04 07 07 05 0a 0c 06 0e 0a 14 19 0d 20 18 0e 1d 1e 1e 28 2a 25 35 41 4b 52 5c 69 6e 7f 8b 95 a3 a5 a8 a8 ab a9 ac bb bf bc ae b6 b8 b7 c3 c2 cb d5 d0 d6 dd e1 e7 ef ef fe fe ff fd ff ff f6 f3 f7 f2 f0 f4 f8 fe ff f7 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fd f1 e4 e2 de dd dc d7 db e2 dc db d0 c3 cd d4 df e0 de e3 d7 dc e7 f6 ff ff ff ff f5 e1 d4 b9 a6 96 86 72 6f 64 5e 55 4e 4c 4e 49 43 38 49 47 51 51 51 38 2b 13 0f 08 0c 0c 0b 13 03 06 05 04 07 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 04 06 05 03 00 06 05 0a 0b 09 05 07 06 0d 0a 0f 11 0e 13 0a 15 17 18 1c 1f 21 28 2d 33 3e 40 4a 56 5e 74 77 7b 8b 89 95 a1 b7 c6 c8 ce ce cd d1 d7 e6 e4 df de da e0 e0 e1 e6 ef ed ec f1 ee ee f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ed ef f0 f3 e3 ee f3 ee ed e6 de e7 e5 f6 f5 f5 f4 f7 fd fe ff ff ff ff ff fa e8 d8 ba a5 95 89 80 75 63 61 5e 64 56 4e 4c 4b 45 46 48 3e 50 50 52 49 3c 32 22 23 16 0d 10 0d 0e 05 06 06 09 06 03 00 09 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 07 07 0f 07 05 07 00 06 05 0c 05 07 0b 03 09 0a 12 0c 10 0d 13 17 1c 20 24 1f 28 37 35 43 50 5d 59 61 75 73 84 8c 97 a5 af bd c9 e0 e3 dd db da e0 ef f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f3 ff ff ff fd f5 ff ff ff ff ff fd ff ff ff ff ff ff ff ff fe e4 d4 c1 af a0 93 84 76 77 65 62 6f 5b 57 58 4c 4c 45 49 4b 43 52 52 4e 50 51 44 3b 2e 26 16 0f 10 0f 0a 0e 06 08 08 02 06 0b 03 03 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 05 06 05 09 00 09 08 04 01 07 08 08 08 06 08 11 14 0f 17 19 22 27 37 38 40 48 54 58 68 70 71 78 82 84 91 9e a9 c0 ce e2 e8 e0 df d3 d1 e0 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e7 df be b3 9c 91 87 7e 7d 79 71 6d 67 56 55 53 43 49 4a 4a 4b 56 59 55 58 55 4e 54 43 38 2f 2a 14 09 03 07 06 05 03 05 06 06 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 05 06 05 0c 0b 06 0d 07 0f 11 0d 10 22 20 2a 2d 31 31 38 4a 51 5a 68 6b 74 76 81 91 96 a0 a9 b8 cb e6 e0 e6 e5 e2 e1 e0 e7 ee f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 eb d8 ce b9 aa 97 94 90 8b 7f 7a 76 6d 5c 63 58 52 55 51 48 57 5f 5d 63 60 5a 4c 48 46 44 3e 38 30 24 10 13 07 07 0b 0a 0d 05 03 06 06 05 09 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 02 06 05 04 04 06 06 0a 04 08 06 0d 11 14 11 16 13 15 24 29 2b 2b 38 3d 3c 4a 52 52 63 65 75 72 80 8f 93 a4 b2 b6 c6 d2 d9 e4 e4 e8 e1 ee f7 f8 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f8 f9 fe ff fb fc f2 ea d4 c7 c2 b2 a5 99 9e 93 80 7c 6c 5e 6f 68 5e 5c 5a 55 61 62 61 64 69 5e 52 54 54 47 46 3f 3c 3e 3f 34 25 1b 14 0f 0b 06 05 03 04 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 03 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 03 06 05 03 00 06 05 03 0a 06 06 07 0a 09 05 04 02 12 0a 13 0d 0b 14 18 13 20 32 36 40 3d 49 4f 4d 60 5f 66 76 74 7e 83 8a 99 a3 af c1 d4 da dc de ef ef eb f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f5 ee e2 eb de de e4 e1 da d5 c3 b6 b3 b5 b3 a7 91 7f 76 75 6d 75 6f 6e 6a 60 67 65 66 6a 67 6b 64 60 5a 58 4b 4a 40 49 40 3f 39 33 30 21 14 12 0f 0c 03 06 06 05 0f 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 05 06 05 03 03 06 05 05 00 06 07 03 06 0c 10 15 19 14 27 27 32 35 3d 3e 43 46 52 5c 65 69 71 74 79 81 94 95 9f 9f ac b6 be d8 e3 ef f0 f6 f1 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fa e5 ef e4 e3 d9 dd cd cf cb c8 c0 bc b6 c2 b0 95 83 76 75 76 79 75 6f 6d 6e 68 65 71 72 6d 6c 64 5a 53 54 53 4e 4e 4f 4e 4d 3a 40 3d 35 20 21 13 11 08 04 0a 05 03 07 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 02 06 05 09 00 06 05 07 07 0a 10 0e 0b 0e 0a 11 10 10 1c 1a 1d 26 31 31 3e 3e 49 54 59 5b 69 66 73 76 80 81 8b 93 a1 ac b3 b8 bd c0 cd db ea f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 fc f3 ee ec e3 de d3 d1 ca c9 bc b6 be cc cc b9 9b 86 7e 86 79 81 89 81 81 78 78 73 74 71 71 65 6f 62 5a 5f 5d 50 56 51 53 56 4c 4c 42 43 3b 32 2c 1b 17 13 11 05 07 01 06 0a 04 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 05 06 05 08 00 06 05 0c 08 06 13 0d 14 13 16 24 30 2c 37 40 3b 4e 4f 60 64 6e 73 7d 7d 85 8c 96 9c a5 a9 bc c8 d9 d2 da d3 dc e7 ec f6 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f4 ed f1 e7 e0 d0 c4 ca be c0 c7 d1 c9 b5 9f 91 89 86 89 84 8b 87 82 82 81 7d 75 73 73 75 68 5f 66 62 5e 60 51 57 51 56 54 4a 4a 4f 4d 4d 32 2a 1e 1b 1d 14 0e 14 06 0e 03 00 08 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 04 06 05 07 00 06 06 03 08 06 11 09 0a 0e 10 12 14 1e 2d 35 3b 34 44 48 54 5c 64 6a 77 83 86 8a 97 95 97 9a aa b4 c0 d1 e0 ea f3 f1 e7 f0 fa fc fc f8 f9 ff ff ff ff ff ff fa ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fc f6 f2 ed e6 de cf cd c5 bf c9 d7 c9 ac a3 9c 87 90 8f 8c 90 95 90 8b 82 89 79 79 71 75 74 6d 68 66 64 64 67 67 60 5f 5c 59 4e 4f 52 4c 46 35 21 25 21 15 0f 11 06 0f 03 0b 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 05 03 00 08 05 03 08 06 05 06 10 0f 0f 14 0f 16 11 1e 24 32 40 3f 3b 3e 45 51 57 63 6a 73 81 92 a4 af b0 b1 bb ba c4 c8 cb e0 f2 ff ff ff ff fd f9 fd ff f8 f0 f4 f9 ff ff ff fe ef f1 f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 fc f4 f0 e8 e1 ce c8 ca d0 ce db d8 c5 b9 aa 9a 9a 92 96 96 8f 8e 80 8c 87 82 83 85 78 71 73 66 75 69 67 67 72 67 5f 61 5d 61 53 5a 55 57 45 3b 2e 22 23 1b 15 12 05 03 01 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 07 05 03 0a 06 12 0c 0f 0a 12 14 18 20 24 2b 37 38 3f 3a 42 44 53 54 5b 6d 67 7f 8f 96 bc c8 d5 e7 e7 e5 e4 e2 e4 f8 ff ff ff ff ff ff ff ff ff fa e5 de dd de e7 e5 e6 eb e4 f2 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fd e7 ec de db d4 cd d5 d3 ea e6 d6 cd c0 b8 a0 9d 9b 99 9a 96 96 8b 8e 87 80 8b 85 7f 75 72 72 70 76 73 79 68 6f 65 60 5e 59 64 58 57 4d 3e 30 31 21 1f 17 14 0a 03 04 06 06 07 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 0b 08 0b 0a 0a 11 05 0b 11 14 14 17 24 36 27 36 3b 38 44 48 4b 4a 56 62 68 66 7c 84 94 ac c3 d6 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 e9 d5 d3 d6 d9 e2 e1 da e7 f0 f4 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fa ea d3 d9 d4 da f5 ff ff e9 d7 d3 c3 b6 b0 a4 99 9c 94 99 92 8e 85 80 89 87 82 78 7a 7a 75 83 73 74 78 72 6b 66 68 61 59 59 59 50 4a 37 2f 24 21 13 09 06 05 00 08 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 06 06 0c 0c 0f 12 08 08 19 1a 24 2e 30 38 38 3c 3e 47 45 4a 4f 53 62 71 69 7a 84 88 98 a9 c0 e7 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e2 d8 d6 e1 e4 e2 e8 ea f0 f1 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d4 ee e4 e4 e5 f3 ff ff ff ff f2 f1 eb d7 bc b2 ad 9c 9e 96 95 9b 96 88 8c 89 85 84 74 7a 82 8a 89 86 85 7e 75 71 74 63 5f 60 5b 55 57 4b 40 38 2e 25 0c 0c 03 0c 07 05 08 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 0a 14 0c 13 0c 0a 18 17 1f 29 2e 36 3b 3d 40 47 4c 51 56 53 5a 5e 6c 68 6f 85 8a 96 9e aa bf d5 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb de e2 e0 e3 ec e8 ee ef fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f7 f4 ff ff ff ff ff ff ff ff ff e7 c8 c3 ad a2 a1 98 9d 96 98 8f 8f 8e 8c 8a 8b 8a 86 87 8b 84 87 7b 7a 73 68 69 62 59 55 5d 5c 5c 58 49 4b 27 12 17 03 09 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 07 0a 0c 0c 11 12 24 25 2b 32 27 3a 41 3d 41 50 57 58 5a 4e 57 60 64 70 7b 81 8c 95 a4 a2 ab c4 cf e0 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e4 e6 e4 ec eb f0 ef f5 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 da d1 be b4 a5 97 97 a2 97 95 92 92 94 90 80 87 84 8b 8e 8e 87 7e 78 75 6d 6d 67 63 68 64 72 68 6a 68 4c 34 13 0e 0b 04 06 07 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 0b 06 05 07 07 0e 08 0c 0d 11 1a 20 2c 2f 3a 3c 3b 36 3f 4c 4e 49 53 62 6b 6b 66 68 6d 76 84 89 8f 9f a2 a1 ad b6 bb c9 d9 e3 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e9 ef f3 fe fa f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 d0 d0 c1 ae b5 a7 a2 a5 97 9a 97 90 94 95 88 8e 8d 8c 85 89 82 76 7f 78 77 6f 6f 70 75 76 7d 77 73 5b 44 30 1b 07 0b 0a 07 06 06 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 06 07 05 03 0d 0c 05 09 16 15 21 31 3a 45 44 48 46 48 4a 48 4f 5f 53 66 7b 77 83 7e 80 87 8f 96 94 a2 b0 b1 b4 b9 c8 cf d7 d8 f3 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f7 f7 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 eb d3 c1 b7 af b0 9d a1 9e 96 93 98 93 95 94 8c 8e 90 8b 83 82 83 85 7c 81 76 73 69 75 7f 84 82 7c 63 4b 3c 22 10 04 06 06 05 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 03 03 06 05 06 00 06 08 04 09 09 0f 10 21 31 32 40 46 45 46 41 50 49 51 5b 5f 61 6a 77 84 88 97 96 91 8f 9f a7 a6 ad b3 bb ba c0 c0 c4 cb d9 e4 eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f1 fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 eb d6 ca ba b3 ac a3 98 9e 9e 99 9d 9c 96 97 8d 96 90 8c 98 95 8b 88 7c 79 77 77 7a 71 7a 8d 8c 84 69 59 41 22 0f 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 06 06 05 03 00 06 05 03 02 06 05 03 06 06 05 0e 13 09 11 21 3b 42 3c 44 4b 41 3c 4b 52 54 57 59 66 66 68 72 89 9a ab af aa b1 b6 aa b5 b2 bd bc b8 c4 c8 c9 c7 d1 df eb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 df c5 bd bc ae a9 9f a1 aa a2 9b a1 9c a1 97 9d 9b 98 a0 99 85 88 79 84 84 82 85 7c 79 7d 8c 84 79 59 43 2c 17 05 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 07 03 02 06 05 03 00 06 08 09 12 15 1b 33 4d 40 3f 4b 45 4d 4a 55 59 66 68 6a 73 7b 75 81 8d a2 b5 cb c6 c8 c7 cc c8 c4 c4 cf cb c3 c5 c7 cb da d7 e7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 d6 c9 bf b3 a7 a7 aa 9f aa ad a8 ab a6 a1 a4 a5 a1 ab 97 90 87 84 87 81 8a 81 80 74 75 79 84 8e 82 5d 47 2d 0f 05 06 05 09 09 06 05 03 00 06 05 03 03 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 05 06 05 03 0f 06 0f 14 10 16 28 32 41 42 4c 4e 4c 50 5c 63 6d 6b 70 71 7a 85 86 8a 96 b1 c3 d3 d9 d6 d9 d9 d4 da da d7 cb c8 c7 ca cb d3 d6 e1 ef fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ed d7 c6 bc b7 ae b3 b6 b2 b8 b1 b0 a7 a8 a7 9d a6 a6 a2 99 8e 89 8f 85 86 88 7a 7d 79 75 7b 85 90 90 6d 44 22 17 0a 06 0a 0a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 04 00 06 05 0b 0f 06 06 10 1e 33 2a 3c 49 44 4e 59 56 59 66 6a 76 6f 7b 78 8c 84 93 a1 9f b2 c7 d5 db d8 e4 e7 e2 eb e3 d9 cd c5 c3 cd d2 d8 da dd ec ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec d6 cf cd c8 c2 be b9 ba b6 b1 a9 a4 a4 9f 95 b0 b2 ab 8d 88 88 96 8e 8b 81 7e 73 6a 7a 87 90 a4 97 6d 42 26 15 10 06 0a 08 08 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 04 06 05 03 07 09 05 04 05 06 13 1e 29 41 45 43 41 4b 50 5f 60 65 73 73 74 80 8f 91 98 92 9e a6 ae c2 d9 de e5 e3 df df ea e7 e4 e2 d3 c8 ca d2 d2 dc e4 e1 ec f2 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e7 df dc d2 c1 c1 b4 b8 b1 ae af ab a4 ab a2 b5 af a5 9b 93 8b 8d 88 80 7d 76 7d 82 84 8b 95 9a a0 77 4f 2e 17 10 06 09 0a 01 06 06 05 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 01 06 07 10 0d 12 15 1e 35 40 3f 42 49 48 58 61 5e 68 76 78 7c 89 97 98 95 9e 9f b2 b9 c4 d5 e0 dd da c8 cb d4 dd d8 db ca cd cf d2 d3 e4 e5 ea ef f2 f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 e9 d8 c5 c1 c3 bc b8 b4 ae ad ac 9d a9 a2 b4 ad a3 a5 a2 8c 8b 81 7e 7e 81 81 88 8c 95 a5 af 9c 71 51 28 20 11 0b 07 07 03 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 0b 0d 06 0e 06 10 13 17 25 3a 43 41 42 50 4d 5b 62 66 70 71 89 89 94 a0 a5 a5 a3 a9 ac b9 c1 d5 d3 d1 ca be bc c9 ce d0 d1 ce d5 d1 d9 d9 e3 e3 f0 f6 f1 fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e7 da cd c4 c4 b2 b5 b6 af ac a2 a0 9c 9b 9f aa ab 9d 9e 8e 8a 81 86 87 7d 7c 8c 98 9b a4 aa a1 7b 49 25 15 16 0b 0f 09 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 04 0a 09 0f 10 12 22 44 4a 49 44 4f 54 4d 56 6a 78 7a 83 8b 97 a2 a9 af b3 af a9 ab b9 c4 cf d0 c5 b6 b5 b0 af bf ca c9 cb d0 d3 dc e7 ec ef f0 f8 f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec dd d3 ce c4 c0 ba b3 ad a5 9a 97 98 9c 9f 9c a5 a7 9f 98 8f 8e 8b 87 85 7e 8b 93 ad ac a3 a0 a4 77 4f 29 19 18 0a 15 08 04 06 05 0d 00 06 05 04 00 06 05 03 04 06 05 03 00 06 05 04 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 05 05 0c 10 10 11 24 33 45 48 4d 47 4b 4f 58 60 68 7a 7e 88 92 a0 a7 b8 ad b8 c2 b5 a4 b1 b5 b0 c0 ae b1 bc b3 b5 b9 bb ca ce d0 ce e0 e4 ed f4 f7 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 df d3 c9 bb b8 b7 ad a3 9b 95 93 a2 9a 9b 9b 99 9b 97 a1 9e 9e 8b 83 88 87 8c 9f b0 b2 b8 b9 aa 87 56 39 1c 11 13 0b 0a 05 06 05 05 03 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 03 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0d 0d 0a 11 0e 13 13 28 4f 52 49 53 4c 4e 58 5f 6b 6a 74 7c 91 a3 a4 b1 c1 ca cd bd a9 a4 a1 ab af aa b5 b1 b2 b8 c1 bf c2 c6 d3 d2 d9 e3 db ea f4 fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f1 df cc c3 b7 b0 a2 a3 9e 9b 91 92 9c 9f a0 94 91 9b a1 a2 a3 9f 8a 8b 8b 8b 83 97 ac bd c7 be a9 8e 60 39 29 12 06 09 08 07 07 05 04 00 06 05 03 00 06 05 03 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 0c 15 13 1c 37 41 5f 63 59 55 59 64 60 62 62 6f 73 83 8f aa b4 ce ca d9 d2 ca b6 ab a3 aa b1 b4 b0 b4 c3 bc c0 c7 be ce da da d4 db e7 e9 f5 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec de d1 c3 b6 af a4 9f 96 99 96 9a 9a 9a 92 9d 95 a2 a5 b3 9b 9a 95 93 93 8f 8e 9e b9 d2 d0 c0 9f 86 63 3a 21 1c 14 09 0e 08 08 05 04 02 06 05 07 02 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 05 0b 10 0c 12 11 19 30 43 5e 69 76 69 5e 5e 61 60 68 62 6a 73 7b 90 a4 c4 d7 e2 da dc cd be aa a5 a8 a8 b0 b5 b9 c5 c5 bf cd d1 d5 d9 d9 df e3 e7 f0 ee fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e8 dd c7 be b4 ae a5 a3 9d 9e a1 9f a7 9f 9e 99 99 98 ab a7 a5 97 97 8a 98 90 97 a4 c8 e0 d9 b2 92 78 65 35 27 15 11 08 0a 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 07 06 05 13 13 16 1f 3b 51 6b 7e 8c 80 6b 60 52 64 62 6a 73 6f 7a 87 a7 c3 e6 eb e9 e6 d0 bb ad a6 ab aa b1 af b9 c6 bf c8 ce d4 db df e1 e4 f2 ea fb f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f0 e1 d1 d0 b9 b6 af a8 ac aa a2 a4 9f a0 99 9e 98 9c 9f a7 a8 9e 97 8f 93 92 8c 98 b5 d7 d4 c6 a8 88 7d 66 42 20 15 09 07 0a 07 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 06 03 05 06 0f 0d 0f 1f 27 45 6a 74 89 97 95 89 6f 67 62 6b 71 6f 72 7b 85 ab d3 ee f7 ee dd c8 be b2 af b5 b9 bc b8 b8 c9 cb cb d7 d3 df e3 e7 ed ed f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e9 d6 cd c2 c2 b8 b6 ac a2 a4 a0 97 a0 95 9b 96 9c a1 a4 a8 a6 97 92 90 8e 8d 98 9d c6 d6 c8 b5 a2 91 77 76 55 31 1b 0e 08 0d 0b 12 05 03 02 06 08 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0d 0c 16 18 18 27 38 5a 6f 8d 9b a3 a7 9b 7c 75 70 74 6f 6e 74 79 8b a9 da fd ff f4 e6 c8 bc ad b0 bc bd bf c2 c2 cb d1 d6 d9 de e2 e1 e5 f1 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e5 dd d5 c7 c1 bd b6 ab b0 a3 a2 97 90 92 a0 95 9c a1 a2 a2 9d 89 95 8c 8d 94 9c ad b0 ba b7 ad a2 90 83 7c 62 46 21 0b 0d 0c 08 14 05 03 00 0c 05 03 00 06 05 03 00 06 0a 03 00 06 05 03 00 06 05 03 01 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0c 0d 13 1b 26 47 60 77 99 a5 ac b2 ae 96 7f 84 80 76 76 76 7e 82 a2 d9 ff ff f9 df cc b6 b4 b9 c6 c0 c1 c7 c7 ce cd da d6 d7 e8 ec ef f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb f0 e5 dc ce cc ba ae b5 ab aa 9f 9f 9d 9e 94 96 a2 9c 95 98 8d 8e 90 86 86 89 93 a2 b4 a9 a8 ac ab 98 8c 7e 76 70 4c 26 19 0d 0e 03 06 08 03 05 06 05 04 00 08 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 09 05 0b 13 19 1f 2e 4a 69 8c 9d b5 bb bc be a6 91 93 8f 80 84 81 8d 95 a7 c8 f7 ff ff ec d4 bc be c6 c9 ca bd ce ce d4 d3 d6 dd e4 ec ec f2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 e9 e4 d9 ca c4 bc af b2 b1 aa a1 a0 a0 a4 98 9c 95 91 99 8f 92 88 8e 8a 82 8b 92 a7 b0 a8 a7 a9 9e 9f 94 8a 83 83 5b 36 15 0d 06 06 06 05 03 00 07 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0a 12 12 1c 26 30 4f 6d 96 a6 c6 cb c8 c9 b3 ac 9c 8d 94 8e 91 99 a5 b0 cf e5 ff fd e9 d4 c0 c1 cc cd d6 d3 dc ce e5 e8 e1 ec f0 e7 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fe f5 ed e4 d1 cd cb be b3 b4 b1 a5 ac a1 a3 9b 9d 9c 99 95 93 8f 85 8a 86 80 84 88 8f a4 a8 ab a8 a7 a3 9c 93 8f 85 84 6f 3c 21 07 08 0d 06 09 03 0a 06 07 03 01 06 07 03 05 06 05 03 00 06 05 03 00 06 05 05 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 03 03 06 05 06 0e 10 11 1f 20 37 45 73 9d bb c7 c4 ca c8 c4 bd aa 94 8c 95 9e a5 b5 c3 d2 ea f6 fe e6 cd ca bf c9 cb da da e2 e0 e4 e1 e9 f0 ed fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f1 f0 ee e0 d5 ce c7 c1 b3 af ae b0 ab a6 aa 9f 9a 94 94 95 90 8c 8a 81 89 81 88 86 90 97 a0 9e a8 ab a6 a6 a9 a7 a1 90 6e 3b 1c 18 10 0e 0d 09 05 06 06 05 03 01 06 05 04 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0b 07 03 07 11 0f 23 28 35 4f 70 9b c3 c7 c0 c5 bc c6 c3 be 9b 8e 90 9a b0 b2 c5 dd e5 f8 fd f1 d1 be c0 bf d1 df ea e7 e8 f4 f0 f4 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff eb e6 e6 df db cc cd c5 ae b5 aa b5 af a0 a2 a2 97 91 95 91 91 8f 86 83 85 7e 78 81 83 8d 9d a3 a0 ab b6 b7 cd b5 a0 8b 6c 4f 2d 1d 0f 07 07 07 04 0e 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 07 05 05 11 0a 1c 23 2f 36 58 77 9e c7 cd ca bf bd c1 ca c9 a7 9d 96 9f a7 b5 b8 da e6 f9 ff ff ec c7 bf be d1 df e3 f0 f7 f6 f8 fc fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fc f0 f1 ee ed dd cf c4 c5 bc ba b6 ab ab a1 a6 a5 a2 a6 92 96 91 91 88 8b 87 7e 84 84 88 83 8f 90 a2 ae b3 c5 c6 b4 96 89 78 52 30 22 1a 0e 0b 05 08 0b 06 08 03 07 06 05 03 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 06 06 09 0b 13 18 24 2b 3e 52 78 9f cb d9 d5 bd ab c1 cb d8 bb a8 a1 9f a7 b2 c2 d9 eb f8 ff ff ff d6 c0 be c6 da e5 eb f1 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f7 f3 e9 e3 d4 cf cb c1 b9 b2 b2 aa aa a5 a2 a0 99 9a 8a 98 8b 90 87 8e 89 82 7d 86 7e 7d 88 89 8f 90 a5 b8 b8 a7 90 89 75 59 37 2d 21 11 0e 05 03 0b 06 05 05 00 06 05 03 02 06 07 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 16 0b 0e 18 1c 30 47 6a 87 af cf e1 c6 a9 a2 ac c4 d9 cf b2 9d a0 a7 b2 be d4 e4 fa ff ff ff eb c8 bc c6 ce e2 eb f3 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 f1 e9 e8 de ce c6 bf bd b6 b1 aa a0 a7 a1 96 95 91 94 96 90 93 86 84 8f 82 8b 84 8a 7e 7f 7f 81 88 90 94 9a 8c 82 83 6d 58 45 29 20 14 16 05 0c 05 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 05 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 06 0d 06 11 09 15 0a 1c 24 2f 4b 69 96 b9 e1 e8 c6 a7 9e a3 ba c2 d0 c1 b4 a9 ab b0 c5 cc e0 ed ff ff ff eb d2 c2 c9 d1 d8 ed f5 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f5 f2 ea e2 cf c9 c6 b3 b4 aa ab 9b a0 a1 94 93 92 93 8f 8a 8e 7d 86 89 89 85 8a 84 7c 86 82 87 84 85 84 89 83 86 88 86 6d 46 31 20 11 06 06 03 0a 06 05 03 01 06 09 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 07 00 06 11 0a 18 16 22 2b 3b 58 75 a0 c5 ef e6 b7 96 9e 97 ac b9 bf c0 bc b1 ad b5 c1 cd d5 e5 e6 f0 f2 e9 cc c7 c7 db e4 ea f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa f5 e9 df d4 c4 b5 b4 a8 a5 a7 a0 9d 8f 91 92 99 95 8e 8a 85 91 8b 87 89 86 88 86 8a 83 89 85 85 84 82 7f 7b 83 84 6a 4a 3b 2a 1d 12 06 03 06 06 05 04 01 0b 05 03 01 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 06 11 0d 0e 12 16 25 32 59 8d a9 db f8 ec b3 9a 89 8c a1 ab b6 b3 b9 b4 b6 bd bb c5 d2 d6 d9 e4 df cd d4 cf cf dd e0 f1 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f7 e9 dd d4 cb bd af af ae 9f a2 9e 90 8a 8b 92 88 7f 8c 89 87 84 86 82 86 8a 8b 87 84 7d 80 85 7e 7d 7b 77 8d 81 77 55 3c 29 18 11 05 07 03 06 08 07 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 05 05 06 10 11 07 1b 23 28 3e 66 96 c4 e6 ff e0 ac 97 8c 87 9a a4 a5 b1 b7 c5 c8 c0 c2 c0 c8 cb ce cd d5 cb c8 ce d9 e2 e7 f0 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f8 f2 ed ec e4 d5 ca c7 b3 ac ac aa a9 a3 99 8d 88 8d 8a 82 8d 8d 8b 8f 8a 88 87 7f 8b 8d 82 82 87 77 7b 7f 7b 7f 89 91 96 7b 5a 39 28 17 12 14 03 01 06 05 03 04 06 05 03 02 06 07 03 02 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0d 06 0b 11 16 15 22 2e 39 6f a0 d2 ee ff da ad 95 92 94 9b 99 a1 ad b8 cb cb bf b8 bd c0 c2 c5 cb cd cf d2 d4 e0 e4 ec f0 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fa fa fc f5 ea ec ee df e2 d9 ce ce ba bc b1 b3 aa a1 9e 97 98 97 8c 8b 91 85 88 90 87 93 86 89 91 88 8a 81 85 89 7e 80 7c 78 7b 80 8d 9f 98 7f 52 3d 2c 16 10 0a 0c 05 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 0e 0a 10 14 1a 2e 45 69 a8 da f6 f9 d0 a9 99 97 95 96 95 96 a5 af bd bc b5 b4 ba bd ba c1 c7 cb d5 da e0 e0 e9 f0 f4 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff fd fe fa f4 f7 ec ea e6 e3 d9 da c9 cf bf c0 b2 ac a9 a5 a2 97 95 97 91 91 8e 8b 87 88 8a 92 88 8e 86 8a 80 8c 86 89 83 84 81 7b 74 76 83 85 8d a1 93 71 56 3e 27 1e 11 06 05 06 07 05 04 00 06 05 03 00 06 05 03 07 06 07 03 00 06 05 03 00 06 05
 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0f 0c 12 1a 21 2c 45 76 a9 d9 f6 f7 c5 ac a1 9d 9a 92 9e 96 a2 b7 b1 bb b7 ad b6 ae bb c7 c2 d7 d5 cf de e8 ef f6 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 fd f9 f6 f8 fe f9 ef f0 ed e4 d7 d3 d2 d0 b8 bc b5 ae a3 a0 9b 8c 8e 8e 8e 89 8b 93 87 8f 86 8a 80 87 88 84 84 7f 83 81 83 85 76 72 82 79 8a 8e 98 a2 8f 7e 5b 3c 2c 1b 0f 05 03 05 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 10 14 11 13 11 23 30 3a 6f a5 d6 e9 e1 c2 b0 a5 a5 a8 a9 a6 a9 a8 ad b0 ab b4 b1 be b3 c4 bf cb d5 d1 db e1 ee eb f2 f6 fb fe fa ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff f7 f7 ff f1 f3 fb f4 f7 ff fb fa f6 e3 e1 e0 d3 d1 c6 c6 b7 ac a6 a1 95 8f 96 8d 81 8a 89 88 8f 88 81 87 8d 8e 90 88 8b 85 84 84 84 7d 7e 7a 76 76 84 8c 9c 9a a5 92 6a 53 42 24 18 0f 05 06 02 06 05 03 00 06 05 03 00 06 05 07 00 07 05 03 06 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 03 00 06 05 03 03 06 0b 03 10 19 17 24 40 6f ac cb e1 d5 a9 a3 a7 9f a5 ab b1 ab a9 ae b2 ae b5 b4 bd b6 b8 c5 c1 ce cf db e9 e7 f5 f8 f4 f6 f4 fe fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f8 f4 ee f8 f7 f0 f0 f2 fe f2 ff ff f8 f5 f0 ee e5 df df d2 ca be b1 b3 a3 95 90 8e 89 94 86 84 87 80 8a 89 89 8b 8e 8b 88 8d 8e 8c 87 8c 7b 7d 7d 7a 7c 7e 91 98 9b 9f a4 8b 70 51 34 23 16 08 08 06 0a 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 06 09 0b 12 11 10 15 31 42 6a 9e c6 d7 c3 a5 a9 a5 a2 a3 a0 aa ab aa b7 aa b6 b5 b1 ba c0 ba be c4 d3 d9 dc e9 ef ff ff fa ea db f2 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ed e6 f2 e9 f9 ee f4 ef f5 fa f5 ff ff ff f5 f5 e6 eb dc d6 cc c8 c3 b5 ab a9 9d 97 8d 87 8c 7f 89 7b 7a 88 8a 8d 85 94 8c 99 93 90 8b 91 84 7c 7f 79 73 7b 8a 8f 9d 91 a7 9e 8f 74 51 45 26 0f 0a 05 07 03 06 05 03 00 09 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0a 0b 10 12 22 33 41 66 9d bb cd b9 a3 9f 9e a2 a5 a2 ad a9 a4 af ad af b9 b4 b6 bd bf c1 ca d1 de eb f3 f5 f4 ed e8 ef ed ed ed f9 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f2 ea e3 e5 eb f0 ee f1 e6 f3 ec ee ff fd ff ff f5 f6 e5 dc d1 ce c7 b2 b6 a8 a5 9d 91 95 95 91 8d 85 88 7c 89 87 92 9b 8b 93 98 95 95 8d 8c 84 82 7f 88 7a 86 91 93 93 a3 a5 a8 82 66 57 3a 27 1d 0b 07 0a 09 09 05 03 00 06 05 06 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 08 06 05 11 09 14 1c 2b 3b 56 8d aa b3 b1 a9 a4 9e a1 9a a4 a0 a6 a3 ad af b3 b5 bb ad b5 b9 c7 d1 d2 d6 e8 ef e9 e1 db d9 db e4 e3 ef f4 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 ef e3 e0 e0 ec e6 f4 f3 e8 f3 ec e7 f2 f7 ff ff f6 ee df d8 d1 ca be ba bb b1 a4 9f 98 94 8d 8c 8c 87 8f 89 8d 89 91 8e 99 98 94 93 8f 88 8b 80 86 7a 7e 80 8a 9a 9c 95 9c a7 a5 7c 65 56 30 27 12 0f 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 07 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 08 07 08 06 10 10 1b 27 37 57 79 9e aa a0 9c 9d a3 a9 a0 a2 a8 a6 a6 a1 ac af b1 b4 ba b0 b8 c5 ca d7 db d4 de d4 da d6 da db e0 e2 e4 f2 ec fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ef ea ed f4 fa f4 fc ec ed ef eb e9 ea f1 f7 f3 ec eb dc d3 d0 c7 be bc bd ae af a8 a0 9b 9b 96 91 8f 8d 85 8e 8e 8f 99 97 94 a0 9d 93 8f 8c 80 86 87 8c 92 96 96 93 93 93 a4 9d 84 68 4a 3d 20 1e 0a 05 06 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 08 07 11 0b 0e 13 16 2a 40 55 79 95 a1 9b 9b 9c 9c 9f a3 9e 9e 9a a7 af aa a7 b2 af b3 b5 b8 b9 c9 cd cd c9 d0 cf d3 cf d2 d0 d3 da e1 eb ee f2 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ed e7 e7 f7 ff fe ff ff ff f9 ea e8 df e1 e2 ee e2 ea e9 d6 cc cd c1 c3 b9 b0 ae aa ae a2 a5 9b 95 92 91 8b 91 90 92 99 9e a4 9c a7 a1 9f 95 93 8a 8c 92 91 91 9c 99 90 8c 9d a1 a1 7e 6e 44 3a 2d 0e 0c 05 03 0a 06 05 06 00 06 05 03 01 06 07 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 06 0a 0f 0b 18 24 35 55 77 91 9f 9b 96 a0 9e 9c 9f 9b 9f 9c a4 a6 aa a7 a4 aa ac b4 b1 b7 c3 c0 c7 c7 be c2 d1 c7 cf d5 d7 da da da e0 f2 ec fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e7 d5 d2 d9 e4 f6 ff ff ff ff f8 eb e0 d5 de d8 df e0 e0 e1 da d1 d0 bf c8 ba b6 ba b5 aa a9 a5 a0 98 9a 98 9c 9a 9a 9b 98 9f a2 aa aa a4 a4 98 97 98 91 9a 9d 9b 95 81 81 8c 9a a2 99 72 5f 3e 3b 1d 14 0b 05 0c 08 06 05 03 00 06 05 03 00 06 05 0c 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0f 08 13 0d 1e 2f 3a 51 73 81 91 96 95 94 9c 9e 9b a0 a3 a5 a7 a2 a3 a9 aa ad a8 ae b0 b2 b4 b4 b7 c2 c1 ce cc d0 cc d5 d3 d1 dc df d9 e0 e7 f1 f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ee e2 de d1 d5 d7 e4 f0 f3 f8 f3 f9 ee e3 df d7 d2 d2 d5 dd dd de d4 d0 c6 c6 bf bb bb be b7 af a7 b0 a0 a3 97 92 97 94 9f 9a a0 a0 aa ad ac a0 a2 a2 a3 a7 a4 a6 a3 9b 92 8b 7e 89 95 9d 8b 78 5d 45 33 1d 0a 0d 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 06 0e 04 10 09 17 2c 38 56 68 89 87 89 96 98 9d 9b 95 97 9c a2 a4 a5 a0 a2 a3 ad a7 a6 a9 ab b3 b5 b9 b4 be bf ca cd cc d1 d1 d2 d6 dc d9 dc e0 ee eb fd fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 ed db d4 d4 d6 da eb e6 f2 f6 e9 f4 e1 d8 dc d6 d2 ce d2 d1 d7 dc cf d3 c5 bd bf bd b6 bc ac b2 aa b0 a4 a7 a1 a4 a0 a1 a1 a6 9f a2 aa a4 b3 ad b1 a9 9e af ac b0 a4 97 8b 7e 79 86 8a 92 91 73 55 47 35 1e 11 06 05 03 06 06 05 03 00 06 05 03 04 06 05 03 00 07 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 00 06 08 0f 03 11 20 2c 33 4d 69 77 7f 86 94 91 9e 9e 98 9e 99 9c 9a 9e a3 9b 9c a3 a7 a4 a2 a5 a1 aa b6 b3 b7 c4 c3 c6 c1 c7 cb c5 c9 d6 da df dd e6 f0 f8 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ee e7 e0 d4 d1 cf df e9 ef f0 ed ea ec f0 d6 dc d7 cf d0 d0 cb ca cf c9 d0 cd c5 c0 bc c1 b4 ba b3 ac a6 a2 a4 a7 9f 9f a2 99 a5 9c 9e a9 aa b0 b5 a7 b9 b9 b1 b2 aa a6 9a 8f 89 7b 7e 71 8f 93 84 70 5b 3d 2a 1f 12 0d 05 06 08 08 0b 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 07 08 0f 0b 19 28 39 47 66 75 86 89 8c 94 90 97 93 94 9b 99 9b 9c 9c 9c a2 9d 99 a4 a6 9e a6 ad a6 b7 ae c0 be bd c2 bf c7 ca c7 c8 d4 d6 d9 e3 e5 f1 f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e7 e0 df d0 d7 d2 e0 e6 f0 f4 f3 f1 e1 e7 d9 d7 d7 ca d1 cd c5 c9 c6 c0 c8 c3 c2 bd b9 bc ae b0 b3 b0 aa a9 ab aa a1 9e 9e 9c a0 a7 a0 a9 ad ae b0 b9 b6 b2 ae af a5 99 8f 84 71 75 79 76 7e 8b 82 6b 4f 34 24 16 15 06 05 03 08 06 05 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 06 06 08 08 10 0f 17 2c 2f 48 66 75 80 86 8c 92 91 97 99 8f 92 94 99 96 9e 98 95 a0 9f 9d a3 a8 ab ad b2 b6 b6 be b5 be c2 c7 c4 c7 c1 cc ca d5 dd d8 e5 ef ea f4 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ea e3 de e0 dc da e4 f1 f3 eb ec ea e3 de e2 db d7 d0 d0 c4 c4 ce c9 c1 c5 be ba b8 b5 b7 af b2 b1 af ab b1 a5 ab a4 a6 aa a3 a9 9e a0 a1 ae b1 b5 ba b9 b4 b2 ac a4 91 85 7b 6f 6d 74 77 7e 85 7d 61 4b 3a 33 16 19 10 05 04 0b 09 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 00 06 08 08 0d 0a 1d 26 34 49 5d 72 82 7f 94 8b 8d 9a 95 90 94 96 90 9d 99 8f 96 97 9c 99 9f a3 a3 ae ac b2 b6 b1 b7 c0 c4 c2 ca bf c2 c4 ca d4 d6 da df e5 ee ef ee f6 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f6 ea df de d8 de e2 e3 ec ef f0 f0 eb e6 e4 e8 df da d7 d3 d1 d1 c6 c9 bd bb bd b7 b5 b4 b2 b5 ae b0 b7 aa a5 a9 ab ad a3 a6 a8 a4 a5 a9 a7 a9 ac af b4 b5 b4 b8 b6 a2 9c 8e 81 7b 78 66 6f 76 7f 82 79 60 4d 34 22 1f 13 0d 05 0a 08 06 07 03 00 06 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 07 03 0a 07 1b 1f 32 42 5e 78 7a 84 81 90 8f 8a 8c 90 97 8d 93 93 91 92 90 9a 99 a1 9e 9b a6 ad ab b9 b3 b3 c0 c1 b9 bd c0 c1 c2 c5 c9 d5 cf da d7 da e7 e9 f1 f7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ec e7 df de df e1 df e3 e4 ed ec e9 e2 eb e6 e1 d9 d9 d3 ca ce ca c1 cd c1 b5 b8 b5 b0 ad ac b3 a8 ab a9 a3 a7 a2 a5 ae ab a7 a5 9a 9f a6 a1 aa a8 b0 b9 ae b7 a8 aa a2 95 86 6f 75 72 6b 64 77 7b 7e 6d 57 48 38 30 25 18 12 09 03 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 08 05 08 0f 08 17 24 2e 4e 5f 73 7b 80 82 8d 90 8d 93 95 97 92 94 96 94 99 92 9a 9b 95 9f 9d a0 a8 a5 b2 b2 b5 b8 bf b6 ba c3 b9 c5 cc c8 cf cf d9 d9 db e0 e9 ec f0 ef fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f6 eb e8 de e6 ec e2 e4 e6 e3 e6 ec e5 ec df d7 e4 e3 d9 df d3 d1 c8 cb cc be c1 b8 ae b1 af aa a8 ac 9d a3 ab a1 a6 a6 9f a7 a0 a6 a4 9e a0 a1 a2 a6 aa ac b4 b0 aa ae 9d 97 83 74 7b 6b 6c 68 71 78 76 83 70 5a 4f 3e 2b 2b 18 10 05 03 05 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 01 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0e 0c 08 11 17 26 2f 4a 59 70 74 79 83 85 8b 91 90 97 9b 9c 9b a0 9d 99 90 99 9b 9a 99 a1 a5 ab b5 b4 b8 ad b1 ac ad b3 b7 be bf c2 c7 d2 cf d4 d6 da dd e1 e7 ed ef f3 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e3 ef e1 da e1 e5 e2 ec e9 ef ea e8 e4 e3 e2 dd e2 d7 d6 d4 d1 cc cd c4 bf be b6 b5 af a5 aa a1 a8 aa a7 b2 a3 9e a2 a7 9e ab a3 a2 9f a4 9f a5 a3 aa ae b4 aa a9 a3 8d 85 80 70 73 74 6a 68 6b 70 75 80 74 5d 51 3b 2d 1c 1a 15 05 03 08 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 1a 0e 19 2a 2e 42 57 6d 74 6f 79 7e 82 8e 88 94 96 96 9d 9e 9a 96 99 94 9a a0 9f a6 ae a7 ac b0 b1 b1 ad a9 b0 b1 b2 b3 b0 bf b6 cc cb ca d1 d7 d8 df e0 e1 eb ea e7 f0 f6 f8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f8 f5 f3 ef ec e4 e4 e7 e5 eb ec ea e5 e3 de df e8 dc e0 d3 d1 d0 ce ca cc bf bc ba b4 b4 ae a3 a5 a3 9e a2 9a 9b 9c 9c a3 90 9b 98 a1 9e 99 9d 9b 96 9f a9 ae ac a9 9c 96 88 7f 7b 75 6d 63 63 67 64 70 79 81 71 57 45 3d 24 22 16 0d 07 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 05 13 11 20 24 3b 41 59 69 73 76 7e 7d 7b 81 8a 8c 92 92 8f 95 98 98 9b 97 a1 9e a1 9b a6 a0 a6 a0 a4 a7 a9 aa aa ab b0 b1 b8 ca c4 c9 c4 ca c8 d3 d3 d1 d7 db dd de eb e8 ed f4 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 ee fa f0 ee e5 e4 e7 e5 f1 ef e7 eb e0 dd d9 d6 de d1 cd ca cb c4 bf b8 be b5 b1 b4 aa b0 a1 a6 a2 9b 9c 99 98 9c 9d 9d a3 8f 98 96 93 97 93 9a a5 a4 a4 a6 a7 9b 89 86 76 72 71 6b 5f 6a 65 71 70 7f 7f 75 56 4e 3c 2e 25 20 0a 05 05 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0e 0a 03 12 16 22 2a 2e 49 55 6a 73 77 76 73 7d 83 80 87 8f 88 91 91 97 95 8d 92 96 94 9f a2 9f a2 a3 a1 a0 ac a9 a6 a9 b0 b1 ac bb bc ba bd c3 cb cb cf d1 d7 df d8 d9 e2 e3 e6 e9 f1 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc fe f6 f4 e9 ef e7 ee f3 ec f0 e8 e4 e9 df d5 e1 df d2 cb d0 c6 c4 b9 b3 b1 b3 b0 a8 a6 a3 a2 a0 99 9e a1 9e 92 9f 94 95 99 9d 9d 99 9f 91 94 99 a3 9f a4 9e 91 90 89 7a 73 6e 74 6e 6b 69 6e 6d 74 84 88 7d 62 4e 40 33 31 15 0a 05 03 07 06 05 07 03 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 06 08 10 25 2f 36 40 57 68 76 6c 73 7b 7c 7e 7d 89 83 88 83 8b 90 91 89 92 90 90 99 9b 96 9e 9e 96 96 a5 a1 a5 a7 aa b0 b5 b2 be be c8 bf c3 ca cc ce ca d2 d2 dd df e7 e2 e9 ed fb ff fa fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ff fb fd ed ef f9 ef f6 e5 e8 e7 e4 df e1 da dc da cf ce c6 c9 c4 b7 b5 b5 ae ab a2 9e 9e 9b 9b 96 92 95 91 8e 8e 98 99 8f 95 96 94 97 8b 95 93 9a 96 9d 9b 8b 89 79 77 75 74 6c 6e 68 68 68 6a 77 85 82 7e 62 53 42 33 25 11 1a 05 03 07 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 04 11 10 1c 2d 2b 48 5b 65 72 68 6d 76 70 7b 82 85 8b 8c 8b 8f 8b 8a 90 90 8f 92 92 99 9c 98 9e a1 9e a1 a1 a3 a3 a9 ba ac b4 bd b6 c0 bd c2 c7 cc cc d5 d6 d8 d2 dd d9 e5 e4 f1 f6 f3 ef f1 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f5 f6 f4 f8 f5 f9 f3 ea ec e4 da dc dd dd d9 cd d0 bd bf bf b2 af a7 ad a4 a1 9f 9f 99 91 94 89 91 93 96 94 97 93 8c 9f 8d 9a 8a 91 96 97 a2 95 93 91 8a 83 78 70 71 64 6d 6d 66 66 6e 75 71 7f 84 74 61 55 40 35 26 1c 0b 05 08 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 06 06 04 08 19 1f 29 3b 45 55 6b 6e 6b 72 74 72 7b 7d 81 86 8a 83 8e 8e 8e 8f 8e 8d 92 94 92 94 98 9b 9e 95 9b 9c a1 a2 a5 b5 af ae b8 ba bc bc c8 cd c5 ca c9 d2 de d1 d5 d6 de de ea e9 eb e7 ec f5 fc f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 f7 ff fc f1 f3 f2 f0 e5 e2 e3 d3 d5 d5 ce d9 c9 c1 c5 c0 b4 ae b1 a8 a1 a0 9a 92 9a 97 95 95 8e 96 8d 8e 90 87 8b 91 90 98 9d 8c 9c 8e 93 99 9d 98 8d 7d 80 7b 79 76 6b 6d 6e 6d 6a 70 75 81 84 85 7c 60 60 47 37 2e 18 16 0a 03 0a 06 05 03 02 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 10 12 2a 37 41 63 6f 6f 6d 68 6c 70 77 7c 80 86 8a 8b 8f 8d 88 8c 8e 94 91 94 98 92 92 98 96 9e 9f 9d a0 a6 a6 af aa b1 b4 bc bd b8 c2 c5 c2 ca ca c5 d1 ce d4 d6 df dd d9 db d9 da ea f0 f3 f0 f2 f4 fb fb ff f7 ff ff f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 fc fa fa f4 f7 f3 ee e6 e1 db d8 d5 d1 cc ce cb bf b2 b7 ae ab aa a1 98 9f 8d 96 8d 95 9c 8f 8b 88 8a 8f 89 85 8c 8f 95 94 96 8e 92 91 92 90 95 84 86 7b 77 73 77 70 6b 72 6c 6b 6e 6f 79 88 8d 82 67 5c 4d 3a 21 1a 10 05 03 00 06 09 03 01 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 07 0b 1f 28 35 42 59 67 6b 73 6c 6b 72 72 79 7d 7f 81 82 8d 8d 85 8a 8c 8a 8e 93 93 91 9a 98 91 9a 9c 9f 9e 9b 9c a5 b1 a6 b0 b9 b8 b7 c2 c1 bd c2 c9 c0 c6 c4 d3 d5 d0 d6 d5 d3 d5 d9 e2 e6 ea e6 ea ec f3 e4 f0 f0 f5 f0 f5 fc f3 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa fc ff ff fa f6 f6 ef ee ef e3 e1 da d6 ce d0 cd c2 c0 c1 b2 af ad a7 9b 96 9b 92 95 8d 8d 90 92 8b 91 8f 88 86 86 84 88 87 8d 8b 8e 8f 89 8c 8c 90 88 89 83 78 6e 70 70 69 6d 69 5e 64 6a 79 7a 78 89 7c 6d 60 41 37 2c 10 14 07 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0d 0a 0c 1d 20 36 4d 54 6b 6e 6d 6d 66 6d 6c 77 7c 80 7f 84 7e 8f 8b 8d 90 90 8e 92 95 93 95 9c a1 99 9b 9d a3 9f 9e 9f a9 ab b7 bf bc ba bc bd c1 bc b8 c4 bf c7 cf cf c9 cb cb d0 da db d1 dc dd e4 e6 e4 eb e9 e6 e9 ea e4 f0 f4 f4 f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff f6 f7 f6 f5 f4 ed ec df de d8 ca cb c5 bf c2 c0 b5 b9 a6 a3 a4 a3 9b 95 95 8c 8e 8d 8b 95 8e 8e 84 8d 88 91 91 85 89 87 8f 89 8f 8e 93 92 92 77 84 75 72 76 6e 6b 6c 6a 68 69 62 66 6f 72 80 89 86 72 63 47 38 2e 21 11 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0b 0c 10 1c 26 30 43 5b 6c 7c 6e 6d 6a 6f 70 6f 73 7f 7c 87 89 88 88 8d 8b 90 8d 96 99 93 9d 95 9c 9d 94 9e a2 9a a1 ab a8 ad af b9 bb be bd b7 bb b6 b6 b9 c1 c7 c7 c3 c4 c4 c6 c7 ca d0 d1 d7 da da e0 dc dd e4 e1 dd e5 e1 e7 eb f2 f9 fa fd f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed e3 d6 cf d6 db d4 c7 ca e0 ff ff ff ff fe f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f8 ff ff ff ff fd f6 f6 f0 ec e1 d2 d4 c3 ca cd c6 bb bb b5 b3 a6 ad 9b 9c 93 93 87 90 91 87 93 8f 8b 90 8a 84 8b 86 86 85 8d 86 87 89 8f 8d 92 90 91 86 83 73 74 70 6f 6e 65 6a 6b 69 6e 6a 68 74 7b 85 88 72 62 51 49 2e 1a 11 05 07 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 01 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 0b 18 28 34 52 59 69 68 6c 65 61 6e 71 73 77 70 76 7a 87 84 86 92 86 88 8b 8a 97 91 90 98 96 97 a0 9c 9f 9b 93 9f 9f a6 ab b3 ae ad ab ae b1 af b2 b0 a6 b0 b2 bc b3 be c8 c0 c5 c9 c7 ce cf d1 d6 d9 dd d6 e1 df e3 e4 e9 e8 f8 ec f1 f3 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e2 cf b5 a6 aa a4 9a 97 92 9a 95 9b 99 a0 b3 b2 c2 bf ce dd eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc fb ea ed e3 e6 da ce c7 c6 c3 c1 bc b6 b9 a7 a2 9a a3 9d 90 8a 80 88 8e 8e 91 8d 8d 92 83 88 80 88 88 85 8a 82 8c 87 7f 8b 84 88 89 84 7e 78 71 6d 6b 66 60 6b 64 6b 60 6c 67 73 74 85 80 73 6f 51 46 2b 1d 11 07 03 00 06 05 05 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 05 07 0a 14 17 29 37 43 54 60 70 6a 70 65 6f 73 74 6e 73 7b 81 81 8e 81 85 82 8d 8a 94 8d 95 94 99 97 95 97 94 a1 9f 97 a1 9c a6 a8 a8 b4 af a3 aa a9 a9 ac af ae b3 ae b3 b5 b7 be bc c5 c6 ba c9 c9 ca cf d4 d9 d6 d4 e0 e2 e4 e7 e8 f1 e7 f1 f6 fd f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb d2 b3 a8 9b 95 86 77 5c 7b 78 71 73 75 6f 75 79 7e 7e 80 8c 94 97 a5 b6 c0 e0 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff f2 f1 f0 ed e9 dd db d0 cc c6 c5 cb be b6 b5 a4 a5 a4 a2 97 97 92 8a 8b 8d 8e 8a 88 87 89 8a 87 87 86 87 7f 7e 80 7f 87 87 8d 84 81 7c 79 79 74 6e 6a 6a 69 67 65 6c 6c 65 6e 69 69 71 84 84 77 66 53 45 32 23 18 05 05 00 06 05 03 01 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 02 0e 17 22 37 48 5d 63 72 61 63 6e 66 69 6e 6b 7b 76 7c 7f 82 8b 82 80 89 90 8d 98 91 93 9c 93 94 95 97 9e 96 9d a0 95 a1 a9 a5 af aa a7 a4 aa a2 a7 a7 a4 b2 a7 ad b5 bd b8 bd b9 c2 ba c3 c2 cb cf ce d7 d0 d3 da d7 d9 e5 ec e2 eb ee f5 fb fd fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa dc b8 92 7d 6e 76 72 67 60 3d 5c 5f 65 5c 61 61 5c 5f 5d 6c 6a 70 77 7c 89 8d 9e c0 d9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 f7 fc f5 f0 e6 e6 e2 dd d8 cd cd c8 c7 c4 b3 b6 b3 9f a3 a2 9c 99 94 89 8f 8f 8d 90 8e 90 8d 88 89 84 80 87 7e 7b 79 7e 8b 7e 7c 7f 83 83 7c 73 74 70 67 64 6d 6a 65 67 63 63 64 64 64 6d 76 82 82 7c 6b 5a 3e 39 16 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0d 1d 27 38 4b 5b 68 64 68 60 69 60 6a 71 69 72 74 78 85 81 89 82 84 83 85 92 93 90 94 92 93 94 8e 91 8f 94 97 92 98 93 a1 9c a5 a4 a8 9e 9d 9f a5 a5 ac ae a8 ae b5 b0 b7 b8 b3 bb ba bc b8 c5 c9 cf cf cf d4 d3 d2 d5 df df e7 e8 e8 f6 f6 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 c8 a9 83 67 64 62 5b 55 57 54 50 54 4c 4a 48 4e 52 54 59 54 57 5c 67 5f 6e 74 76 88 98 b1 db ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe f4 f8 f9 f2 fa fc f2 ec e9 e0 da d9 d2 d1 c9 c7 c3 b7 b9 ac ab aa a3 96 99 8e 8e 8d 8c 83 83 82 94 88 8a 8e 81 7e 7e 7c 81 7e 7f 7d 7e 71 76 7a 73 7d 74 71 7a 67 69 6c 64 64 66 62 64 6a 61 71 65 6c 71 82 8e 73 6a 5e 45 2c 1f 19 05 07 01 06 05 06 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 0e 13 24 37 48 55 67 70 67 64 5f 62 62 68 72 6e 74 75 83 80 83 85 86 83 85 85 8c 8c 8d 94 8b 93 93 95 99 97 99 98 94 99 9c 9f 9f 99 99 9e 9d a5 a2 a5 a1 a0 a6 a5 a9 af b0 ae b2 b4 c0 c4 bc c0 c9 c1 d7 cd d1 d4 d7 d8 d6 de dc e1 f0 ec f8 f8 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff da a6 7d 6c 5c 5a 57 51 50 50 4e 4b 4e 4a 4e 46 45 4a 50 4f 47 54 50 59 5c 5e 5e 66 70 88 9d be e7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fb f8 f3 ef ea f4 ec f2 ec e5 e2 d9 d6 d4 d1 bd bf c1 b9 af b3 a5 9d 9f a5 91 99 97 89 88 82 89 93 86 85 7e 7e 7e 7e 80 7f 7c 70 75 7c 7d 7b 74 82 71 78 71 76 6f 6a 6c 6c 74 6a 6c 5d 5f 63 6a 68 66 67 68 7d 83 78 70 57 4b 37 24 19 05 06 04 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 04 06 05 03 0b 0c 1e 26 32 49 60 65 6f 6c 66 5a 67 69 6c 6d 6f 79 73 78 84 83 84 81 85 89 8e 90 89 90 91 8c 90 8e 92 90 94 9b 97 9f 90 97 9c 9a 99 9b 9f a4 95 a2 99 a1 a1 a4 a7 a4 ae a4 af b0 b4 c0 b7 bd c9 cd c1 ca cd cb cb d2 dd d5 e0 e1 e0 e5 f2 f0 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 bd 89 6f 60 56 4e 4a 48 3c 47 49 41 42 46 41 45 45 44 47 41 39 4b 4f 43 54 55 55 60 62 72 83 97 ce ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f7 f2 f5 ec f4 f0 f0 ec ec e4 df dc d6 ce ca c5 bf c2 bd bc b1 b2 a4 9c a2 93 94 8d 82 87 86 92 8e 8e 8b 83 84 80 7d 75 7b 7d 6c 80 73 75 77 79 70 76 71 78 6d 71 69 6d 63 5f 61 66 64 63 63 5f 6a 60 63 66 6f 7d 7c 6b 63 50 3e 24 0d 0e 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0a 06 14 24 31 45 59 63 6b 6d 5a 5a 65 60 66 66 67 6d 73 75 77 7c 7b 74 79 85 8a 94 8c 8a 89 8b 8c 8a 8b 8d 89 96 93 8c 95 92 95 97 99 9e 96 95 99 98 9b a5 9c a3 a2 a0 a0 a2 b0 aa b3 b2 b9 b6 c0 c6 c1 c6 c1 ca ca d5 d0 cd d7 e0 e0 e6 e8 f3 ea ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d9 9a 75 6c 5d 50 45 3b 44 42 3c 40 3c 38 3e 40 38 3d 40 41 3a 42 40 3c 44 3d 4b 4e 53 5e 69 6e 8a c8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f9 fa f8 f4 f6 f2 f3 ef f1 e5 e8 ed e9 e0 d5 d6 d1 c5 bf c5 b7 ba b7 ae a6 ab 9c 9c 9b 91 8f 8b 8c 87 89 86 90 84 86 83 7b 79 77 7c 77 6c 74 70 78 76 69 75 68 75 73 6c 78 66 64 64 64 67 62 62 69 67 66 60 5d 67 64 65 68 75 77 6e 61 4b 3c 24 1f 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 07 0e 16 2a 37 4e 5a 6a 6f 71 66 5f 68 63 66 69 6a 70 6d 73 79 77 87 7b 7e 84 84 89 85 8f 8e 8a 8e 90 92 8f 8a 92 90 8f 94 94 8f 95 94 93 90 9c 9c 94 96 9a 9d 9e 9c 9b a2 9f a9 aa ad b3 b5 b6 bc c5 c4 c1 c0 c7 cc c7 ca d0 da dd df e5 ea ea ef f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe be 8f 76 62 53 3f 3b 36 3a 3c 41 3a 36 36 36 3a 33 3e 3d 3d 43 37 33 37 40 39 3d 4d 4d 56 5f 6c 7b ac f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe f8 f6 f7 f5 f7 f2 f6 f1 e8 ec e6 e4 e6 e2 e0 e2 d4 d1 d5 c8 c7 c2 c0 be bd a9 a7 ac 9c 95 98 90 92 8b 85 88 7b 87 81 85 83 7c 82 7b 73 72 74 72 71 6d 6a 6d 6f 70 71 71 75 71 70 67 67 60 60 62 62 67 61 66 5f 5c 63 64 64 5e 6c 65 6a 70 5c 56 3d 2b 1b 15 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 03 0c 10 20 28 3c 40 52 72 72 68 64 63 5d 6b 63 65 69 6f 6b 71 76 77 7c 83 82 87 89 89 82 8d 8b 89 81 8e 8e 8c 8d 8c 91 8c 8b 92 94 90 95 93 93 9b 92 96 9e 96 9d 9c 9a 9e a5 ab ab ac a9 b4 b5 b9 b6 b6 bd bf bc c8 c4 bf cf ca d5 d9 d2 dd e3 e2 ed ef f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ac 7e 6d 5a 48 3b 37 31 3a 3c 30 2f 36 34 35 3a 34 38 31 47 42 3b 34 33 34 2c 35 3e 46 52 55 6d 7a 95 e3 ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 fb f3 ec f2 f6 ec ef e9 e7 e1 e5 e7 e0 dc e0 e0 e3 d5 d3 c8 c7 c4 be c1 b9 bd ab a5 a1 95 9f 8e 8b 87 89 8a 84 81 8a 82 83 7f 7e 79 7d 6f 74 76 77 70 70 68 70 67 70 75 71 67 67 6e 74 67 64 62 64 69 66 63 64 6c 61 69 5b 5b 5d 60 70 6c 70 5d 58 48 32 22 14 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 19 14 28 38 48 56 6b 70 65 63 5c 64 66 65 61 66 67 68 6f 6f 6d 7c 80 82 85 8d 8b 80 87 87 88 8c 8c 8d 80 7f 8b 84 8a 8f 90 8a 92 8c 99 8a 92 92 99 94 90 95 91 95 9f 9f a1 a6 a5 a3 b5 b0 b7 b1 bb b4 b9 be c7 bf c6 c6 cd db d7 dd d6 e5 e5 e6 e8 f1 f8 fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 a3 74 6b 48 3f 32 2b 38 30 35 35 30 2f 2f 2e 2c 34 34 37 41 35 36 35 32 31 37 35 3b 3c 39 51 64 6b 98 d7 ff ff ff ff ff ff ff ff ff ff fc fb f2 f4 f8 f0 ec ec ea ee e8 ed e5 e4 e3 df de e1 e2 dc d3 d0 d6 ca ca c7 bd bb bf b1 ae aa a6 a5 95 97 97 8d 87 87 87 80 88 81 7d 83 7c 7f 7a 74 72 6f 6f 65 69 6b 69 70 68 69 65 6e 64 67 6e 65 62 64 61 62 61 61 61 66 62 5d 62 63 5d 59 5d 62 68 6c 65 58 43 30 23 0b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 0d 1c 24 44 54 60 6b 6a 66 5c 58 57 58 65 5e 62 69 68 6f 75 6f 78 73 7c 80 82 85 84 83 81 80 80 85 84 87 8a 7e 89 89 8b 8b 8f 8b 8e 8f 89 92 9d 95 97 96 98 95 91 9c 9d a2 a5 a0 ad a5 b2 a7 b2 bb bc c3 c2 b7 bf c1 c6 c6 c5 d4 db d6 d9 db df e9 e7 f9 fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd a3 76 69 45 38 2e 2b 30 2e 26 32 2c 2e 2f 2a 33 2f 2d 33 3d 44 39 2e 2e 31 31 35 30 32 3a 3d 58 74 9d e3 ff ff ff ff fd fb fa fd f7 f8 fe fb e3 ea ee e7 ec e4 e7 e1 e4 db de de de dc dc dd e0 da d9 d1 d1 d1 c8 c2 be bf be b7 b3 ab a1 96 92 95 8a 84 80 7a 84 86 82 82 80 7f 77 74 6e 77 6c 6f 75 6f 64 60 60 6b 6d 71 69 68 64 67 66 64 62 5a 66 64 65 5d 66 63 60 63 5e 60 53 5b 5c 5a 60 65 69 52 4d 2d 25 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 05 0d 14 1e 27 37 4f 60 6b 70 72 65 57 53 5e 60 62 6a 64 72 66 6f 71 74 7f 80 85 81 84 88 85 86 7c 7e 7a 84 87 8b 8a 91 8f 8f 89 8b 91 90 8a 94 86 8f 98 91 93 91 93 98 98 9c 9a a1 a9 a5 ac ac ad b0 bb b9 bc b5 b8 bb c7 c2 c4 c8 d1 d1 d9 e5 e5 df e5 e6 f6 f0 fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff a9 7c 60 3d 2f 2d 24 2c 30 2e 31 25 20 2a 27 2e 32 2c 39 42 42 38 2c 29 2f 28 33 37 37 3b 40 54 74 a8 e7 fb ff ff fc f6 fc f8 f7 f9 e7 ea ea f1 e0 ea e3 e5 e4 de e2 e3 db d7 e3 d7 de e1 da d9 d5 d8 cc cb c3 c4 bd c1 bd b9 b2 ae ad a8 a2 9b 8a 85 7b 80 80 78 84 7f 80 72 78 79 78 76 72 6a 72 6b 64 64 67 6c 71 64 6b 6b 68 75 64 6a 65 5f 68 67 60 6a 61 5f 65 68 66 67 57 56 5e 5f 58 58 60 61 52 4d 38 24 1b 07 05 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 13 17 1a 30 3e 45 64 62 71 70 5d 56 5d 5f 5c 66 61 62 6b 6d 66 6d 74 6d 7c 82 86 86 87 83 87 83 8a 80 87 80 7b 87 8a 8a 8c 86 8b 90 8f 8f 8b 87 8c 8b 92 90 94 99 95 93 9f 99 a0 a9 a6 ab a5 ac a9 b1 ab ba b5 b6 bf b4 bd c6 cc cf d2 d0 d3 db d8 e6 ea f2 f1 f6 f8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c0 89 5d 3d 2c 27 22 28 2d 25 24 26 2a 2a 2e 2c 28 2d 35 44 3d 3f 2e 2d 2f 35 32 27 2e 36 46 43 78 ba e9 f1 ff f6 f9 f2 f2 ed e8 eb eb e7 e7 e3 e2 e2 df e0 d6 d9 da d4 d3 ca d9 d1 da db d4 dc de d4 d1 c5 c8 c4 c0 b8 b6 b5 b2 af a2 a2 9c 93 8a 84 79 70 75 79 81 73 76 71 73 6c 6c 70 6b 66 69 66 66 68 66 64 67 68 60 69 64 6d 5e 5c 68 59 5f 67 63 61 61 60 63 5a 5a 5c 5a 5c 55 5a 51 52 5e 5e 55 50 37 2b 0f 06 02 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 0f 10 22 34 42 4e 54 60 70 65 58 5e 5a 60 5c 58 66 66 6a 6d 6a 74 64 71 7c 7f 84 84 84 83 80 7d 82 81 86 84 89 8b 8d 83 8f 8b 8c 8c 86 8b 87 88 87 82 91 93 8f 89 95 92 94 9a 9d a4 a2 a5 a8 a6 ab ab b5 b6 b8 ae bb bb bc c7 ca c5 cc cd dc d8 de dd e3 ef e9 f5 f4 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d9 89 60 33 2d 20 25 24 29 2b 26 23 27 1f 24 29 20 29 35 3d 4f 3c 2c 27 30 32 30 31 36 3b 3d 4e 74 c7 ec f2 f7 ed ee e8 ee e1 e1 de e6 df e1 d9 db e0 de df d4 d2 d3 d5 d3 d0 d2 ce ce d5 d1 d2 cd ca c9 c4 be b7 c2 bc b1 b2 a1 aa 9e 9d 93 91 8b 82 72 6c 7d 76 75 6e 72 73 71 73 63 70 6b 64 66 61 64 5f 63 64 5e 5d 6b 66 63 67 60 67 60 64 60 67 61 66 60 62 5e 58 5c 53 52 53 50 54 5a 57 57 59 58 4d 44 29 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 13 18 27 2e 3a 54 5e 66 6c 5f 55 53 54 67 5f 5d 64 5c 66 65 73 73 70 73 72 72 7d 7e 84 86 80 8c 84 82 83 8c 82 87 8c 84 8c 83 89 88 84 83 88 89 8b 92 8a 89 90 93 94 96 92 97 9e 98 95 a0 a7 a1 a7 ae a1 b1 ab b5 b4 bb b5 bb c4 c5 c9 d0 d1 d2 da dc e5 e9 e6 f0 f4 f0 ff f9 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 8e 57 3d 2b 26 23 24 29 24 20 23 28 21 22 26 2c 2e 32 3e 43 39 35 2a 31 35 31 33 31 39 35 42 67 c4 e2 f3 f1 ea ec e7 e3 e1 dd db df d9 dd d1 d2 d0 d6 d2 d0 d6 c4 cd ce c7 cd c7 cb c7 cc d3 d3 ce c5 bc bd bf b9 b4 b1 b1 ae af 97 9d 97 89 85 79 7c 76 76 78 76 6b 71 6d 6d 70 68 6d 62 5d 60 6a 69 62 61 5c 65 62 64 64 64 66 5f 5f 68 5f 5e 5f 5d 64 5f 5a 55 58 4c 5f 54 5a 54 5b 52 4f 58 5e 54 53 3e 27 15 04 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0b 05 15 1d 2b 37 37 4f 65 5b 67 62 59 55 53 5a 63 5e 62 65 5e 65 69 68 68 6c 73 74 83 79 7b 87 83 7e 85 85 87 90 8e 8d 8c 8a 83 85 8f 8c 8e 8b 84 8a 8e 8d 84 9c 90 86 90 97 95 9a 9e 95 9a 9f a5 a3 a5 a9 a8 af a6 a7 af b4 b8 bd c1 c4 c7 c3 d2 d3 d8 d9 da e6 f0 e8 f1 f3 f2 ed f6 fa f8 fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb d7 89 58 33 2d 24 25 20 28 1b 25 24 1f 22 24 23 1f 20 26 3c 4a 36 2c 2f 29 34 36 33 2f 2c 3a 42 69 bb da e6 e8 e4 e5 d8 dd da de d7 dd d4 ca cb cc c3 cd ca cf ca cc c3 be cc c6 cd cd c9 cd ce c4 c2 b6 ba b2 b2 b6 b1 b4 ab a3 a3 97 9a 8c 7a 74 7b 77 75 72 6a 70 72 63 69 70 6c 6a 62 62 60 63 61 64 66 5c 65 63 62 65 66 64 62 62 64 5f 60 66 67 59 5d 61 59 62 5d 50 5e 5e 54 57 4c 59 4d 56 58 5b 57 42 2a 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 15 1e 25 2f 49 56 5f 6d 66 59 55 4f 50 54 5f 5d 66 5b 64 63 5c 6d 6e 6e 73 6b 80 79 80 80 87 88 85 8b 89 82 8a 87 89 84 84 86 80 86 8b 7f 87 8d 84 82 86 88 8b 87 8e 8f 92 93 93 92 a0 97 a2 a3 a3 a9 a7 ac a6 a9 ad ad b2 b9 b9 c1 c1 c4 ce c4 d2 d7 d7 de e0 de e9 e8 ee ec f1 f4 f5 f4 f8 f2 f5 fd ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e8 9b 54 30 22 21 17 1e 1a 1c 1f 1e 1b 1b 22 22 21 27 28 3c 57 31 35 26 24 30 2e 35 35 38 34 42 62 b6 dc e5 e5 de d9 d3 d9 d8 d0 cf d5 cb cd c8 c6 ce c5 bf c4 c7 c4 bf c3 c2 c4 c6 cd cb cd c8 c9 c1 ba bb b0 af b3 ae a6 a3 a0 a5 8f 93 89 7b 73 74 72 70 71 69 69 6a 68 6b 6d 5f 5d 62 65 62 5f 62 5b 5a 5e 5f 5e 57 5f 61 5e 61 54 5e 64 61 5e 5a 59 65 55 5e 61 56 57 55 57 4c 56 4e 4a 53 4e 56 55 4c 48 27 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 11 19 1c 29 3d 40 50 5c 60 64 56 51 55 5e 5b 5d 57 67 62 6d 60 65 6b 62 6c 6b 70 75 78 7e 83 84 7e 82 8b 84 8b 8f 8a 84 8c 81 8b 84 86 86 82 84 8d 8f 85 8d 86 83 8d 8f 8f 90 91 94 91 98 a1 94 a0 a6 a5 a4 a3 a7 a9 ae b4 b6 b6 b9 ba c5 c4 c4 c6 cc ce ce d7 dd d9 e1 e7 e4 df ea ed e6 ea ed e7 f0 f6 f4 f6 ef fb fa fd f9 fe fa ff fb fa ff f1 e0 a8 59 33 27 22 22 1b 1f 1b 18 1d 19 19 1c 23 20 26 25 3e 5a 3b 2e 21 30 35 2e 31 33 43 3f 42 60 a9 d4 dc df de d5 d4 d8 d5 d1 ca cd be c5 bd c8 c0 c3 c0 be bd c2 bb be bb c0 c7 cb c9 c5 c7 c1 c5 b6 b9 b0 a8 ab a8 a4 a6 9d 9f 8e 86 8b 80 72 6d 6d 70 68 76 70 61 63 64 6f 62 64 62 5b 5d 64 64 5c 5f 64 65 5e 5d 5b 5f 65 5c 68 5d 64 61 5a 5f 55 63 60 63 59 56 56 5e 4f 59 52 59 51 49 54 57 53 51 40 25 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 06 05 16 1a 20 2e 36 3f 4f 63 69 62 52 52 49 51 65 5f 62 61 5c 64 65 62 68 5c 62 6f 6a 73 73 71 7e 7d 7f 86 81 82 8f 83 8b 87 7f 82 86 86 83 88 85 86 8a 80 81 86 91 8a 87 8e 8e 8a 8e 93 90 9b 94 a3 9b 9c 9f 9b a4 a0 ab a8 a8 b5 b3 b6 bf b8 bc c5 c4 ce cb cd d5 d0 cf dc d5 e0 e1 dc dd d9 dd e5 e0 e5 ed e7 e8 ed ee f2 f0 f0 f1 f9 f5 f0 f2 f6 e4 d9 a2 65 3b 22 22 1c 19 1d 1e 1e 14 18 1d 24 1a 1e 1d 28 3c 53 43 25 2a 24 2f 35 34 41 38 40 44 63 b8 d4 da db d5 d2 ce d5 ca c9 c5 cc c0 c2 ba bb c5 bd bd b8 b8 bf b3 bc be bd bb c7 c1 bc c4 bb bd b4 af ae ad ad ae a4 a1 97 99 8c 87 81 71 70 71 70 68 6b 6a 66 68 67 68 66 60 5e 65 65 61 5a 57 5f 5c 61 5c 5f 5b 69 5b 64 5f 5c 61 60 5e 59 5a 5a 5d 5f 53 5a 57 54 5b 4b 50 4f 4c 52 50 4f 56 5b 52 3e 1f 10 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 0a 1f 23 29 3b 49 60 63 63 60 54 53 52 52 54 5e 59 60 60 59 69 63 5c 63 61 6d 70 74 74 71 7b 79 76 79 86 8e 7e 89 85 85 78 80 8a 86 85 89 8a 81 84 86 87 7d 8a 86 83 86 89 8e 8f 8b 92 91 98 98 99 9f 93 9f a1 a5 a6 a7 a1 a0 aa ae b5 b6 b4 c3 bc bc cd c8 c8 cd c7 c8 d6 ca d7 da d8 d8 d7 d9 d8 db da dd de e2 e5 e8 ea e8 e7 e1 e7 e8 e7 e1 d6 d0 a2 65 34 20 13 15 1a 13 1d 1e 18 13 16 19 16 15 1c 27 31 3f 38 26 29 27 2b 31 35 38 3d 47 48 5f a5 ce d5 d4 d2 cd c6 c5 c6 c9 c3 bd c0 bb b1 b6 b3 b5 b7 b0 b2 b3 b3 b4 b5 bf b9 be b9 b8 b5 bd ac ab ad a7 a1 99 9c 97 92 98 87 89 81 7e 6f 6e 70 64 64 65 5e 64 61 60 63 61 5e 5f 64 58 56 5f 5a 5f 64 5b 61 63 5d 63 59 5f 5d 62 5b 5c 54 57 58 5b 5d 61 5c 52 53 56 53 57 55 53 4f 50 4a 50 58 59 4d 38 25 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 05 0b 0c 0e 20 22 2b 3d 45 53 5f 64 61 55 55 55 50 55 55 4c 59 59 5e 63 60 61 64 64 68 68 70 73 71 77 71 71 78 7f 83 7d 80 79 86 85 85 90 7d 80 84 83 7d 8c 7d 87 84 87 94 7e 84 94 90 90 8a 8e 95 94 97 93 90 9a 94 9c 9e a4 ae a6 ad aa a7 b0 b0 b7 bb bb bf c3 ba cc c8 c9 cb cf cb c6 c7 ce d3 cf cd d0 ca cc d6 d9 d4 e5 d8 de db da de e8 e0 dc d5 db ce b0 6b 3c 1e 18 15 18 1f 19 16 14 11 20 1f 1a 19 1b 25 3d 46 36 38 28 31 33 3a 41 37 44 44 4e 62 a9 c9 d9 ce cc ca c6 c7 cb b7 be bd bb b2 b4 a9 ae b3 b1 b6 b0 b1 b7 a9 ad b9 be b4 bb b6 b3 af ab ab ae a7 a5 9f 9f 98 8b 90 85 7f 83 76 70 67 69 70 67 60 61 62 61 61 68 59 67 5e 57 5a 52 59 59 62 5c 5f 5a 5a 57 56 5e 59 5f 5a 5d 69 5c 5d 5a 51 60 58 5e 58 58 5b 53 56 50 4a 50 4e 4b 4e 56 59 4c 31 18 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0a 09 0d 0c 17 25 3a 40 46 58 60 69 61 5c 50 51 50 55 52 59 5c 5e 55 61 5b 67 6a 61 69 6a 6c 71 6a 68 70 77 6f 80 80 88 7e 7e 83 80 7e 86 82 84 86 82 82 7d 85 7d 82 87 84 8a 88 89 8d 8c 89 92 95 99 91 90 96 8d 98 96 99 a0 a2 a5 a0 a7 a8 ad b2 b5 b8 b2 b8 bf c1 c3 bd c7 c6 bf c5 c6 c2 c8 b6 ca c0 d1 cb ca cb d3 d0 d0 cf d5 d7 d6 db da de d7 d3 cc c7 a5 61 30 20 14 14 1b 16 19 14 1a 18 19 19 1d 12 27 22 36 4a 3e 2d 2d 29 30 37 39 43 48 48 56 67 b0 d2 d1 d5 d0 c8 be c4 c2 b6 b4 b8 a8 b5 a8 ab ae a7 b0 b3 a6 b0 a7 b2 b0 b9 b9 b7 bc b6 b1 b0 ab ac a3 9f a4 9b 9f 94 89 89 86 7c 77 77 65 5f 6b 63 61 65 5f 61 64 61 5e 6a 65 60 60 5b 5d 55 5d 60 5a 61 5d 54 5f 68 57 5d 5a 61 52 58 55 5e 60 5b 5a 5b 64 61 53 54 52 51 55 4e 50 43 48 51 50 54 49 3b 15 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 06 0a 12 12 2b 2d 40 53 59 64 73 61 55 47 4b 50 4a 45 55 58 5e 63 5f 5d 5b 67 61 59 6a 68 67 71 6d 6a 6c 6f 70 74 77 7a 7e 84 82 77 7d 83 81 7d 7e 82 7b 83 7d 85 7e 84 89 88 86 89 8e 8c 91 8d 8b 90 8e 96 8e 89 92 91 93 9b 97 a0 a4 aa a9 a4 ac ae b4 b1 b1 b4 be b0 bb bd b4 bf ba be c1 b9 b8 be bd bd c1 c2 c4 c4 c9 c5 ca c7 c7 c6 c9 cd cc ca c4 c3 a5 6c 37 1c 11 0c 15 0a 17 12 13 0c 0f 14 1a 16 26 24 2b 48 42 2e 30 2c 31 3d 45 43 4d 55 5e 67 b6 c8 d6 ca be be b4 bc b7 b3 b1 ac ad a1 a4 a1 a5 ad a3 a0 a2 9f a6 ab aa b6 b3 af af ae a8 a3 a6 a4 9f 93 9b 9a 91 8f 8d 7e 7f 74 68 70 65 6a 67 64 62 5e 5e 62 58 68 5e 5c 60 58 5e 57 51 59 56 5f 56 5b 5e 63 5b 5f 59 55 59 59 5a 58 56 5d 56 54 56 59 5c 5c 50 54 4e 51 49 4d 4b 45 47 4d 51 4c 3b 2e 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0e 08 0e 1b 22 34 3b 46 55 65 6f 64 54 4d 4f 4a 58 50 52 59 54 59 66 5c 60 5e 5c 5b 65 64 74 6e 67 6a 6b 6f 6d 76 6e 74 71 78 76 84 82 7d 7c 81 80 80 84 78 82 78 7d 87 7f 82 88 83 84 8e 8c 8b 94 8c 99 90 8d 8c 92 93 92 9c 97 9f a7 a9 a5 a8 a9 af b3 ae b1 b6 b4 b4 b2 b4 b5 b1 b0 b0 b5 bc b8 b4 b3 bb b4 b9 b7 ba c6 c0 bc c4 bb b5 b9 c2 bf bd c9 b5 a6 6d 2f 18 13 19 11 10 18 19 16 14 10 13 0e 16 18 28 32 4a 47 38 30 35 3e 45 48 5f 67 6c 72 7f b6 d4 ce bf b9 bf b4 c2 b2 ae aa a2 a2 a7 9f 97 9f 98 a2 a3 9f a5 a5 a3 a6 b4 b6 ab b1 af a2 a5 a4 97 9f 9a 9a 8b 8c 84 83 78 79 70 6d 6a 65 5f 60 62 5f 5f 56 61 63 61 5d 64 5e 63 59 54 52 59 55 4f 59 5a 58 5a 53 5f 59 5a 59 59 56 5c 57 59 58 59 5d 55 5e 5a 55 51 50 4a 4c 46 47 43 46 4d 4c 4a 38 20 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 0f 15 1b 27 3f 3f 4e 5e 6f 68 70 5c 54 50 53 4b 4c 47 51 52 56 62 5a 60 64 62 5a 5c 67 69 67 64 66 62 68 77 6c 6b 78 77 7e 7a 7f 83 83 79 7b 80 79 80 7e 79 7c 7c 7f 85 80 86 83 8a 8b 92 8c 8e 8e 85 90 8e 8d 90 8f 91 97 98 91 99 9f 9d 9a a8 ad a9 a6 ad ae b3 b3 ad b4 b1 b7 a9 ad b3 af b6 af af b4 b2 b6 be b1 ba b7 bb b8 b4 b6 c3 ba b0 b9 b4 ad 98 73 2a 1b 14 10 17 11 11 18 0c 0d 0b 14 1b 17 1f 21 36 4e 49 43 33 2f 3b 41 50 7a 8e ad af ae cb d8 d3 c9 bd b4 b2 b4 ad a5 a7 a9 a8 a6 a0 98 9a a2 9a 9b 97 9a a1 a5 b2 ad b3 af a7 aa 99 a0 9b 9c 9b 94 96 8e 84 82 7e 7e 76 6c 6c 6c 65 64 64 67 5b 5a 66 5c 61 5b 5f 5b 62 62 5b 5a 5b 5a 62 56 54 5c 5e 57 58 5c 55 59 5d 58 57 5a 5b 5e 5b 5c 5f 5e 5f 5f 55 53 4e 49 49 49 49 4c 3f 46 4a 3b 2c 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 04 06 0e 18 15 31 2d 3d 51 58 6b 74 73 6b 54 52 51 47 4f 4a 59 54 5a 61 5f 60 64 5f 5a 63 61 64 69 68 62 62 64 68 70 6c 70 72 76 72 77 7e 7a 74 85 7b 74 7b 82 76 7e 83 84 79 78 80 82 82 87 8d 86 84 8d 8c 8d 8c 92 8d 8c 8d 94 95 97 9b 98 9d a2 a2 a8 a9 a5 a8 ab a8 a2 a1 aa ad a5 ad aa b1 ab a7 9c a7 af a9 ad b3 a9 b1 b2 a5 b1 b7 ba aa ae af aa b7 a6 92 69 30 1d 0f 08 18 0f 10 0c 08 11 0e 15 1a 14 29 27 32 43 44 3a 34 3a 37 58 79 b3 e7 ff ff ff ff f5 d4 c3 b7 b6 b2 b3 aa a4 a2 9f 9b 9b 9a 9e 9d 99 a2 9d 96 98 97 9f ab ad b0 ad a7 9e a4 9d 9c 97 8d 94 85 87 80 79 7d 73 6b 60 62 68 62 63 63 52 57 5b 5b 63 54 56 5a 5d 52 64 53 58 50 52 5a 56 55 54 5a 5b 57 59 4d 56 54 5d 5a 5d 5e 5b 5f 5b 57 55 58 57 51 50 48 49 48 4a 48 4c 3b 3c 3d 33 25 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 09 12 22 26 35 49 53 5e 6c 65 70 6a 5e 4d 50 51 4d 51 50 51 56 5d 5d 5d 58 5e 64 67 61 65 61 63 63 6a 65 69 6a 6a 6d 70 6e 73 74 6e 79 76 73 79 76 75 77 76 79 7b 7a 7b 78 81 85 85 8c 8a 80 85 92 87 8e 8d 81 92 84 90 88 92 94 94 94 9f 9e 9e a4 97 9f a9 9e 9d a9 a6 b1 a5 a9 a4 98 a7 a1 a5 a8 aa ac ad a5 a4 a5 a4 a7 ae a3 b0 ae ad ab a9 a8 a7 9f 93 62 2b 15 0b 0b 11 10 11 15 17 06 10 0c 0d 20 20 1a 29 3d 38 35 31 3b 45 6d af f5 ff ff ff ff ff ff ed c6 ab a5 a8 ad 9e 98 95 96 9e 97 9a 8f 99 9c 93 8f 99 a4 9a a0 99 ac a6 a6 a2 9d a3 90 90 8f 8e 8e 87 87 7d 79 6f 75 67 66 65 60 5f 56 5a 5c 5b 61 53 5f 59 5f 5a 61 5b 54 5a 55 53 56 59 53 58 55 51 58 4f 5b 57 58 5a 59 64 57 65 51 55 5c 53 4e 57 4f 41 4e 52 43 49 4b 48 43 38 42 38 29 18 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0d 10 1f 24 2f 4a 4b 66 71 71 6f 68 62 4c 53 45 4a 4e 4a 54 51 51 58 59 60 58 60 66 61 62 63 62 64 62 65 66 65 64 66 6d 69 67 6f 74 71 74 76 79 74 7b 7c 82 76 7b 7a 7d 7e 7d 82 7a 7e 84 91 8f 8d 87 8a 87 94 89 8e 93 8c 8e 96 92 99 94 9b a1 a0 a1 a2 a1 9e a1 9f a8 a3 a8 a5 9b 9c a3 9a 9c 9c a2 a7 9e a1 a4 a5 a4 a4 a4 a0 a2 a5 9f 9f a2 9c 9b 98 8e 59 2d 17 09 0d 0c 13 0d 13 0e 0e 06 12 18 14 1f 21 29 3a 44 3a 33 35 4d 82 e3 ff ff ff ff ff ff ff fd ca ad a0 a0 a4 9c 98 94 92 90 99 8e 94 93 92 94 90 92 94 96 9b 9e b1 a4 9f 9f 94 96 96 91 86 84 83 7b 7f 78 7a 71 71 6d 63 64 5e 5a 5e 5e 53 5d 53 63 5b 57 5e 58 5b 53 57 5d 5b 5a 51 58 57 5b 5f 5a 5a 4c 5a 56 59 54 5b 58 5d 59 59 58 58 55 55 51 52 50 52 56 4a 4c 45 4b 40 3b 34 25 22 1c 09 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 10 15 19 2e 38 45 50 5c 6a 70 7a 73 64 4a 50 4a 53 44 4f 4d 51 57 58 56 56 59 5e 65 66 68 62 63 67 64 60 64 61 63 6b 64 68 69 63 69 6d 6e 6d 75 72 71 7a 6f 76 7c 82 7e 78 7b 7c 83 80 87 83 8a 87 86 8a 8d 91 89 82 8b 8b 8b 86 91 96 9a 9a 95 9d 9c a4 92 a2 9e 9a 9a 9e 9d a0 9e 9f a1 9b 9d 94 97 97 98 9e 9a 96 a0 99 9d a4 9c 97 9a 9c 9f 95 94 93 7d 55 23 1c 14 05 0e 09 0a 0f 0b 0e 09 0a 11 16 13 1c 23 46 3d 38 36 38 54 a5 ff ff ff ff ff ff ff ff ff c9 ac a0 96 98 91 90 8d 8f 91 8f 8f 89 8b 91 91 8e 92 99 9a 9d 98 aa 9d a4 9f 8b 93 8b 8a 88 84 7d 79 7b 74 70 6f 60 68 62 64 5c 5b 5a 59 59 5f 56 56 4f 53 5b 59 58 55 56 5a 53 4f 4f 51 59 53 51 56 53 55 51 5e 59 5c 5b 5d 64 57 5e 5a 52 51 51 4d 4c 4f 4d 4c 49 48 45 42 44 3c 31 26 1c 12 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0d 17 1d 31 31 40 50 5c 67 68 7c 72 65 55 4a 50 48 4c 53 41 48 4c 4d 4c 56 5d 5e 57 63 5e 5a 6e 5e 62 5a 5d 62 62 67 62 64 6b 65 63 67 66 74 70 71 68 71 70 6d 75 72 75 7d 7c 71 82 82 7e 87 88 91 87 8a 8c 88 8b 92 87 86 90 8f 8d 8f 92 90 97 9b 98 9d 99 93 9a 97 9b a0 93 9e 97 9c 92 8e 97 99 91 98 9b 92 98 9a 9e 9e 95 9a 95 92 96 91 92 92 87 8d 7f 55 23 12 09 06 0a 07 0b 10 0b 09 0d 07 0a 0f 12 1c 22 32 38 36 36 38 6c b7 ff ff ff ff ff ff ff ff ff d0 ad 9d 9a 8a 88 8d 8b 8f 8f 8a 8e 95 8a 90 89 94 89 96 8c 9e 96 9f 96 9d 9d 8f 95 8a 85 88 76 7c 7e 72 77 67 6f 69 62 60 66 5c 5a 58 5b 5c 5a 5a 51 56 53 59 57 62 54 4b 4f 51 52 55 4e 4d 56 56 57 56 51 57 57 56 60 61 59 57 51 52 51 52 4d 55 4a 47 4a 49 49 4c 46 44 36 3f 2e 31 1d 10 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 21 2c 34 41 4b 5c 6c 6d 7c 76 6c 5b 57 44 44 49 45 49 4e 4e 4c 54 4a 59 51 54 56 5c 66 67 63 62 60 55 66 5f 59 65 64 61 61 67 6e 63 71 6a 69 6e 70 76 74 6d 70 74 73 75 81 7b 7f 7a 81 85 84 86 84 8a 83 8e 8c 86 91 8f 8c 90 93 93 99 8d 8f 8d 96 93 9a 9e 98 9b a2 8e 92 94 87 92 92 93 8c 8e 8b 90 94 98 8e 98 8d 9d 90 94 90 90 94 8f 90 8b 85 74 4a 1c 0e 07 11 09 10 0b 0e 04 04 15 0d 11 10 13 17 20 37 3d 39 38 3b 63 b4 ff ff ff ff ff ff ff ff ff cd a5 97 94 90 8c 81 88 84 86 8a 85 85 83 86 8b 8b 8b 99 8f 9c 98 9a 9e 9b 93 8d 84 87 80 7e 71 76 79 70 6d 71 63 6b 6d 5f 5e 60 5b 5d 5f 57 56 5d 56 57 5b 58 53 52 53 59 51 56 4b 4f 50 56 59 56 5a 54 53 56 5c 5c 5c 64 53 5f 54 4f 56 4b 53 50 48 4f 4e 53 4e 50 4d 41 3d 37 31 25 16 11 09 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 1c 1a 2d 49 4d 5e 6c 69 78 76 77 62 55 48 4f 4c 4e 4f 4f 52 58 55 49 4f 4f 4d 5e 61 61 60 5a 5e 5f 5a 61 64 57 5b 5c 64 61 67 61 62 64 68 6e 6a 68 6e 73 71 76 71 71 78 74 79 7a 79 83 81 84 83 82 8d 81 8a 8a 86 8d 8c 84 90 91 90 94 95 94 8c 93 94 92 93 8f 97 97 9e 95 91 92 8c 8a 8c 97 91 92 93 97 92 8b 99 88 89 91 96 92 8c 86 87 81 7e 80 74 4a 1e 14 0a 08 0c 0d 12 17 08 0b 06 0a 07 0d 18 13 22 29 38 3a 2c 45 58 9b f8 ff ff ff ff ff ff ff fa c3 9d 94 8c 8b 8b 84 84 7c 85 81 88 89 8a 89 80 85 86 8c 90 88 8e 95 96 94 8d 83 84 7a 77 75 80 75 76 73 6c 62 65 59 62 5c 57 63 4d 5b 58 55 59 56 55 55 52 50 56 54 54 56 58 4f 4d 50 57 54 50 54 58 4f 52 5e 57 55 59 5f 58 51 4d 51 54 46 50 4e 48 4e 4c 4f 4a 48 4b 3c 3e 32 21 22 12 16 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 0e 1a 1d 32 34 41 54 63 62 70 7b 78 61 4e 4d 43 41 4f 47 48 45 51 4d 46 51 4b 4f 55 54 5c 54 57 58 50 5b 5b 60 61 5b 5c 63 5f 61 60 66 60 60 63 62 67 6b 6e 6a 71 6b 78 71 6e 72 78 73 75 7e 7e 81 7d 86 88 90 8b 82 89 89 8c 8d 8e 8e 87 83 96 93 8c 89 90 9a 85 9d 8e 8a 90 88 91 89 88 8b 8a 86 8f 8b 8b 91 88 8c 88 87 87 7e 86 87 83 7d 7c 74 76 69 49 22 0e 06 05 03 08 0a 0f 0c 06 06 05 0b 0d 0a 0e 13 2e 31 2e 2b 34 48 7d d0 ff ff ff ff ff ff ff dc a9 8f 86 85 8b 83 83 81 80 7f 80 7b 86 81 83 84 89 7e 87 8c 8d 86 88 90 8d 85 80 7d 7f 81 7a 72 6b 6f 6c 64 67 61 60 5a 52 57 59 54 56 59 57 52 54 57 51 4d 55 55 4f 52 4c 4d 56 46 44 51 53 58 50 4a 54 4f 56 55 5b 54 5a 4e 5a 42 4d 4a 48 4d 51 49 4f 47 4d 4b 45 3e 34 39 35 1a 14 0a 0a 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 18 24 2f 31 43 50 5f 65 78 76 79 6d 5d 4a 4b 44 4e 45 4e 48 4c 51 50 45 4e 4f 53 55 51 4f 4d 55 58 5b 63 5e 5d 59 5b 5e 5f 61 61 5c 64 56 65 6a 60 71 6c 70 6a 6a 74 70 70 7a 75 6f 76 79 78 79 7a 7f 86 85 86 8d 86 89 86 82 87 8b 8c 91 8f 8c 8d 8c 88 92 90 8f 8e 89 94 94 90 8e 8d 85 92 91 83 8b 8f 84 85 85 86 7d 86 83 88 7d 79 7b 78 72 76 6b 4a 1b 14 06 0a 0e 06 07 0e 0b 01 0a 06 06 08 10 0b 14 2c 2f 2a 2e 29 42 63 95 df ff ff ff ff ff e8 c1 a3 90 88 89 86 81 76 73 78 78 7f 7e 7a 7b 7c 7c 79 7b 82 87 8b 8b 92 84 88 7b 83 7a 76 71 77 74 6e 6a 5f 62 6b 60 5b 60 5a 5c 5a 4e 51 52 56 58 56 4d 54 54 52 52 55 51 4e 4d 4d 54 4e 58 52 53 52 59 5c 57 53 5a 5a 54 51 59 52 46 4a 4a 4f 50 4a 50 50 44 45 46 3d 3c 34 37 29 23 19 0e 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0b 10 20 2e 26 38 4c 54 5e 70 71 79 6a 5e 53 49 4b 4a 47 45 4c 42 49 47 44 4b 47 4a 4c 50 4f 51 50 5b 5e 61 64 61 5b 5c 5d 54 5a 5a 5e 60 65 5c 5c 64 66 63 63 6e 6a 6d 73 77 71 6c 73 75 7a 7a 7b 7d 82 81 7e 82 84 81 7c 80 89 85 8d 88 8c 88 8a 8a 8d 90 90 8d 8e 8d 8a 8d 86 87 8e 8a 8b 86 86 8b 8b 8a 82 83 84 80 7c 84 80 7c 76 77 76 6d 6a 6c 65 45 15 0f 06 06 05 0e 0b 0c 03 09 06 05 05 04 06 18 0f 26 39 21 21 2d 2b 4d 66 99 c0 e5 e2 ce be b4 a5 a0 8c 87 7c 7b 7d 7f 79 79 76 7a 70 71 7d 7b 74 7e 7a 82 7f 85 85 88 7e 81 78 7d 7c 76 6e 73 74 6f 6c 65 61 5c 5e 59 5c 57 5c 51 5d 56 51 55 53 53 54 4b 53 55 56 51 4e 4d 4d 4e 4c 55 57 4a 4a 53 56 64 55 5d 55 54 4e 59 56 58 51 45 49 44 4a 4d 49 53 4a 4c 47 43 43 30 2d 2a 1c 10 08 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0f 11 29 26 37 47 4d 5e 65 7b 6f 74 65 4d 3f 3c 44 49 49 4c 47 4f 41 49 40 47 44 47 50 4b 50 50 53 5e 62 5e 5f 67 67 60 5e 65 5c 5b 58 5a 58 5f 5a 62 66 68 68 6b 66 67 70 6b 74 77 72 6e 78 74 79 7e 80 84 7f 7f 77 7b 81 83 7e 81 80 7e 85 87 8a 7d 87 89 85 84 89 84 88 81 87 8c 88 88 88 7f 88 82 83 7c 7a 83 7f 86 7a 80 7d 72 72 7b 71 66 6c 66 50 17 08 06 05 0d 0b 06 09 03 00 06 05 04 09 0d 09 17 1c 28 20 18 22 29 2d 45 54 6f 84 7d 7f 7d 9a 9a 91 8e 87 80 7c 7c 75 74 76 78 76 77 6b 72 71 79 81 80 81 87 7e 85 88 77 84 78 7d 78 71 73 76 6d 6b 69 67 5a 5c 56 56 57 54 5a 54 55 52 56 54 51 52 4c 4e 53 4f 4a 52 50 4d 56 50 4c 4e 4c 4c 50 53 4d 52 52 52 4b 53 56 4e 4c 48 46 4a 50 41 49 48 53 40 4e 4e 41 43 37 31 2d 1f 10 06 08 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 16 22 2a 2f 3c 43 53 64 73 7d 77 64 54 43 44 43 45 49 45 4e 43 45 45 4a 53 46 4b 4d 48 51 4e 4f 62 62 64 67 64 64 63 61 5a 5f 61 5f 63 5d 62 5f 65 6d 62 6d 67 69 71 72 66 70 73 6e 7d 75 6f 73 76 78 7d 84 75 83 7a 7b 81 84 86 8a 86 85 7a 7f 81 81 82 84 85 85 80 82 86 89 8d 89 88 88 85 82 7c 76 7e 79 71 7e 7a 76 78 73 72 69 74 79 6a 64 66 41 16 05 0a 05 03 03 09 07 03 05 06 05 05 04 0f 0f 13 23 21 22 14 16 1c 25 36 33 45 49 4e 50 55 7a 90 86 85 7e 73 7b 77 73 76 79 74 7c 70 75 7b 71 7c 70 76 79 7f 85 80 84 7b 78 75 75 6f 6d 66 67 62 60 6d 67 64 64 5b 61 59 5c 5e 4e 4e 50 4f 4b 56 4f 54 4f 52 50 4e 4c 50 4c 52 47 49 4d 4f 49 54 51 53 54 50 55 56 58 5c 52 4a 4a 4a 45 4e 49 52 51 4e 43 44 42 44 47 38 34 2a 24 0d 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 14 14 26 25 38 3d 4d 5c 62 6d 77 64 4f 44 44 4a 4b 4b 51 4c 49 40 4e 42 4e 3f 45 4e 51 44 48 50 50 60 67 6b 6b 61 5d 5e 59 5f 5a 60 60 5c 5f 5c 62 5d 6d 67 5e 6a 6a 6e 68 73 72 73 72 78 73 79 75 75 6e 73 7e 7f 7f 78 7d 81 7b 7c 84 7e 84 86 7d 80 89 7f 85 80 81 81 87 89 84 84 7d 84 85 85 7e 7b 7f 81 87 79 77 7b 75 73 72 69 69 6b 62 58 5c 41 14 09 06 0d 06 08 06 06 03 0b 06 0b 04 05 06 0e 0e 19 25 15 12 0a 14 22 28 2c 2f 31 33 29 42 70 83 8b 7e 81 71 7a 7b 76 6b 72 75 6d 6d 6e 76 75 6c 74 7a 80 7c 86 7e 81 75 76 73 75 6b 6b 73 6a 66 69 66 5b 61 5e 5b 5b 5b 5a 53 62 5b 50 55 55 4f 51 59 49 4f 55 54 56 55 57 51 49 48 4e 52 4c 50 52 53 4b 52 54 58 52 4d 55 50 57 4f 55 4f 52 53 4e 47 46 43 45 43 42 38 2e 1c 20 19 0b 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 16 1c 2a 26 3a 3a 45 60 6d 72 67 58 43 40 45 47 48 4a 43 4a 3a 36 3e 40 46 49 3d 49 45 46 46 4d 5a 62 67 6d 71 5a 55 59 5d 57 60 57 5b 5e 61 5f 66 65 66 5f 6e 66 60 70 6e 6e 6e 70 72 74 68 75 71 76 6c 71 74 72 78 7e 79 7b 7a 77 81 77 7d 7a 7b 89 74 7a 80 84 83 83 86 88 7e 83 80 7d 81 7d 78 7a 6f 77 75 72 75 77 6e 6c 69 6b 65 62 59 5c 3d 14 09 06 05 0d 00 06 05 03 00 06 05 03 03 0b 06 12 1c 16 0d 0a 0a 0e 15 1c 20 1a 21 1a 27 30 60 7c 79 80 75 69 6e 72 6d 72 70 64 71 70 6a 6d 67 75 75 76 7f 81 79 79 79 6d 78 6d 71 6e 68 6a 6b 66 6a 5f 5e 5c 5d 55 59 51 5b 5a 54 53 50 57 5a 52 52 4b 4f 43 50 4b 4a 4e 4d 4c 59 4a 4c 55 48 51 52 54 52 56 50 5c 53 4f 56 4d 4a 50 4b 4a 4e 54 49 4a 3f 45 45 3d 3f 33 22 27 15 13 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 14 14 20 23 27 38 35 4f 62 69 60 4d 44 47 3b 4a 44 46 3f 43 45 44 43 3f 48 4d 47 3f 44 53 4a 4c 58 55 63 65 66 65 62 66 61 5f 58 58 5c 51 5a 57 5d 64 62 65 69 66 6e 5f 6e 70 64 6f 6d 6b 73 67 72 6d 74 71 75 6f 76 78 75 73 78 75 7b 73 73 7a 7c 7a 7f 86 7d 79 7a 7a 80 85 7e 81 80 7c 75 75 71 77 7b 7a 75 70 72 69 74 70 6e 69 57 5d 5a 56 44 12 0a 07 05 06 00 06 05 03 05 06 05 03 00 0a 0b 0a 14 17 16 04 09 11 15 15 11 14 15 1b 18 2f 5b 7a 78 73 7a 69 74 72 6c 70 6c 6d 6e 66 6a 6e 6f 73 70 71 78 76 7d 6e 75 76 75 6a 73 66 6b 66 64 5d 66 5e 62 5f 60 5c 5e 5c 51 55 4f 4b 4d 51 4a 53 51 4d 4a 52 53 51 56 50 4d 56 54 51 54 53 52 56 55 51 4a 52 48 4c 59 4d 4f 4f 47 58 51 4b 47 47 47 42 43 3b 3c 42 3a 37 1f 1c 18 0c 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0d 12 15 20 28 31 31 43 4e 54 60 4f 45 43 45 40 49 45 49 41 48 47 47 44 41 41 4e 4b 42 49 3e 47 52 57 5f 63 66 5c 60 61 5f 5f 63 5f 5a 58 55 61 60 5d 6d 6a 67 64 69 65 63 66 6f 6a 72 69 6b 74 71 77 67 6b 6d 78 6d 75 75 70 7a 70 7e 79 79 75 7d 77 80 79 7f 7f 79 80 83 77 86 83 76 76 75 74 75 6e 70 79 78 70 72 71 6c 6a 65 62 62 5d 5f 55 3b 15 0a 07 05 04 01 06 08 04 08 06 09 03 00 0b 0b 06 0f 0f 0e 07 05 06 08 18 0e 15 1c 1b 20 1d 53 77 71 70 72 65 6f 74 75 65 6f 71 6d 6a 6f 77 70 73 7a 76 77 7d 76 73 77 70 67 76 72 69 6b 6e 6b 61 63 63 60 5c 5b 57 5a 58 5a 59 60 56 4e 59 50 54 53 4e 4b 47 52 54 55 59 52 53 5a 53 58 5b 5a 58 55 59 56 55 51 5b 5b 4c 4f 45 57 57 54 52 54 42 4b 49 45 4b 39 3f 36 29 21 15 11 0c 02 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 0e 11 21 20 26 35 37 38 43 44 4a 44 41 47 3e 3e 46 42 3a 48 41 46 42 44 47 44 43 44 44 43 46 44 4c 53 5a 65 56 5b 5a 5e 63 63 5a 57 5d 54 5a 5e 5d 60 58 67 69 63 65 66 5e 6b 65 6e 63 6d 6b 67 6a 61 6b 70 64 69 6c 74 6b 6e 69 6a 75 76 69 77 72 79 7a 78 7b 7a 78 6c 80 75 7a 7e 76 72 72 74 72 70 64 64 67 65 68 6b 6b 5f 5e 55 57 5a 4f 40 17 06 06 05 08 00 06 05 03 03 06 05 03 05 06 09 07 14 12 0d 04 0e 0a 0e 0b 0e 0f 0e 0c 1a 16 56 69 7b 78 6e 6b 6f 6b 64 6b 65 69 6b 69 64 6b 63 6f 75 79 7b 77 70 6a 73 67 6f 6c 6d 6d 69 66 66 65 5d 61 5f 63 60 58 55 58 50 58 53 50 50 52 51 4e 4d 4b 4b 51 4a 5a 57 55 51 51 53 55 4f 4f 55 5b 54 5a 4f 50 48 4a 51 51 50 4f 51 4d 4d 51 41 46 48 4a 46 47 3b 39 35 31 1b 15 0c 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 0d 15 1e 24 27 2f 35 3f 42 41 46 3d 47 44 41 43 38 45 3d 42 46 42 49 48 47 44 50 43 47 49 49 45 55 52 5f 61 66 6b 5d 56 5e 51 5b 5a 5c 58 5b 61 64 5e 5b 5e 5f 64 65 67 61 68 68 68 5f 63 62 68 60 66 67 68 67 69 66 6e 70 6e 77 71 6f 6b 76 74 78 79 69 72 74 6f 79 73 6f 70 79 74 73 6c 6e 68 72 6e 67 64 67 6c 62 5f 5f 63 54 54 4d 54 3c 10 06 06 05 03 02 06 05 03 05 06 05 03 00 06 05 09 08 0f 0d 03 02 0a 05 10 0b 15 14 0d 0a 1d 43 70 73 6c 6b 63 62 66 6b 64 63 65 64 6b 65 6b 6e 70 74 78 76 77 6d 6e 6d 66 66 73 69 69 6b 69 6a 64 62 6b 61 5d 59 5b 5a 56 53 5a 4f 4e 4f 57 4f 52 4e 51 58 57 5c 59 55 52 52 5a 49 4a 50 5a 4d 49 49 53 4d 4a 52 4b 4a 4f 4b 4a 54 4c 4f 47 45 4c 3c 44 40 41 3b 37 32 21 1f 0c 09 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 17 24 29 2e 33 33 39 3d 37 44 3e 44 3b 47 3f 49 39 42 3d 3d 44 40 40 48 44 41 42 46 48 4a 56 54 57 60 58 65 68 57 5d 60 5e 55 53 52 51 59 52 62 5b 5e 66 5f 68 5e 60 65 6d 68 63 63 60 66 64 63 6e 66 6f 6d 60 69 6e 69 6d 71 69 6e 73 6f 73 68 6b 6f 73 6c 73 75 75 74 73 6a 71 74 76 69 6f 71 67 6d 6b 69 64 67 55 5e 5e 54 50 5c 4c 36 14 01 06 05 0a 00 06 05 05 00 09 05 03 00 06 05 04 0b 06 06 03 04 0b 05 03 0f 07 0b 0d 0a 19 49 6d 69 72 65 5e 66 6a 69 6b 6e 5f 61 66 6e 71 72 79 7a 72 79 6c 6d 67 71 6e 6a 62 6c 68 64 6f 63 61 60 5c 58 59 5e 5b 51 54 51 56 4e 4f 56 4b 5b 57 59 56 58 53 59 55 57 62 5e 57 4b 46 49 50 4c 4d 56 54 57 4a 4f 4e 4c 52 59 4e 50 47 4c 43 4a 47 4a 47 42 3e 37 3c 30 25 11 15 0d 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0f 18 23 27 34 33 35 3b 3b 3e 3f 44 3a 46 40 46 42 38 39 44 3c 45 45 49 4a 45 46 48 4a 4a 4d 47 4d 53 59 5c 5b 5a 57 5e 56 53 5a 5a 57 57 5e 52 5b 56 5e 64 5b 5d 69 60 61 5e 65 63 5e 67 67 60 5e 5d 67 63 62 6d 6f 6d 66 6a 5c 6a 70 69 71 64 6c 6b 73 66 67 6b 71 74 6d 75 6c 6c 6d 60 6d 68 60 5e 5f 6d 62 5d 5f 63 59 59 4e 52 4e 3a 0f 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 01 10 0b 03 00 0a 05 03 09 06 08 0d 0c 14 44 61 6e 71 6a 5c 6c 6d 59 6e 64 6f 67 66 69 67 6d 6d 69 6e 66 67 65 65 69 61 68 63 6f 69 67 63 5d 5e 60 5c 5e 58 57 55 54 55 54 51 4f 4b 49 52 55 53 58 55 5d 62 5a 56 50 59 5b 51 54 47 4f 51 54 4b 52 4f 44 46 4a 4e 45 49 50 47 48 42 49 44 46 46 45 41 3f 38 40 31 2e 1c 13 0e 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 09 1b 1c 22 2b 33 2f 3a 36 41 37 39 42 45 43 4a 46 40 43 43 43 42 41 46 47 49 42 4f 47 43 4a 41 4b 54 59 5f 5d 4d 52 57 52 4b 54 54 53 4e 52 56 5d 50 56 57 55 5f 5e 5e 5d 5b 5f 5a 69 57 62 5d 61 61 64 65 65 6e 6c 66 6b 60 6c 6b 6c 65 6e 63 6d 6d 61 63 68 6b 6b 6e 64 5e 68 65 68 66 64 66 5f 61 57 62 65 64 5c 55 53 50 4e 51 49 37 0e 03 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 09 07 09 0e 01 0f 3d 63 66 6c 64 61 6a 61 65 5e 68 61 65 65 6c 6d 69 72 7a 71 73 6a 70 65 66 62 61 67 64 5d 62 67 65 61 60 5b 57 4e 5b 52 5b 51 4f 53 54 4f 4c 53 55 53 50 56 5e 60 59 50 56 52 54 4a 4b 4b 52 49 45 4b 4b 46 4b 49 51 54 51 52 49 49 46 49 4d 4c 45 46 47 3e 41 3d 32 32 21 14 09 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 10 21 1e 23 33 36 37 36 3e 43 3a 36 3d 45 44 41 3f 3b 3f 44 43 42 4a 46 45 40 3c 4b 46 48 49 44 48 52 59 57 54 59 56 52 54 54 58 51 5a 52 55 52 54 58 59 53 54 60 59 60 5a 59 60 5c 64 5e 5f 60 58 58 67 60 65 65 5d 5e 6b 67 69 6c 5a 67 6b 6b 6c 67 6d 5f 67 67 5f 68 6e 65 63 6c 61 62 5c 68 64 5b 5f 59 5a 57 5e 58 5b 55 4f 52 3e 11 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 08 0a 00 07 07 09 02 0a 34 63 64 72 6c 6a 65 64 67 5e 6a 66 69 6a 64 6a 70 6f 74 69 64 6c 64 62 6a 61 64 5e 6c 5c 6b 68 63 63 60 5c 5b 4f 55 52 58 52 54 54 4c 4d 55 58 55 52 5c 5f 68 60 57 50 53 52 4b 4c 4f 46 52 4a 4c 4d 50 46 4a 4e 4d 4d 46 4f 4f 45 4d 48 4b 49 49 4a 41 42 43 31 3b 23 23 17 0b 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0c 17 28 29 27 2c 36 39 44 40 3b 44 3e 45 4e 40 42 44 3e 3f 45 48 47 44 3c 46 43 4a 50 4e 47 4d 4a 4b 4e 4f 53 53 56 58 55 53 52 56 56 4f 53 53 5a 5b 58 56 50 5e 58 55 5c 56 5a 51 57 57 5c 59 63 57 5d 5d 5e 62 60 58 61 60 5d 5a 60 6a 60 65 6b 69 5c 67 66 64 66 65 6b 63 67 6f 65 5e 66 64 64 5e 61 5a 5d 5b 61 5b 50 57 52 56 40 14 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 06 06 04 0d 14 32 5e 6a 6c 67 5c 63 68 68 66 67 62 65 69 64 70 6c 71 72 6f 6c 65 60 66 68 5b 61 6d 60 64 5d 5b 63 58 57 5f 54 5e 5e 5c 5b 59 58 59 57 50 4a 5c 5a 55 5d 57 60 5a 55 4d 5a 51 4a 51 4a 49 4b 49 48 4c 4f 48 4c 4d 54 4b 4a 4c 4f 49 47 53 48 43 43 49 4a 42 43 31 2e 26 1d 1a 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 18 23 29 32 3d 3d 3a 38 41 37 40 3d 42 3a 46 3c 45 4c 46 45 44 3e 3b 42 3e 4a 49 48 38 3e 49 4d 4a 4b 56 54 55 50 4d 50 55 4d 4d 50 50 54 4a 57 52 61 56 51 50 60 52 59 57 56 5c 60 60 52 5b 4f 58 5b 59 56 5a 5b 5e 61 62 63 5a 64 5f 65 61 5d 65 67 5e 5c 67 6a 5e 63 67 6c 67 60 5f 5f 62 5a 5f 59 5b 59 53 58 57 5a 4f 52 3e 16 00 07 05 04 00 06 05 03 00 06 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 05 09 07 32 53 6e 64 62 60 64 6b 67 69 68 65 68 70 66 72 6e 63 6f 6b 67 67 64 63 65 68 5f 64 5d 5f 5c 62 62 5d 5f 5e 53 56 59 54 56 51 54 52 52 54 55 53 59 56 53 56 54 54 4c 49 4f 4a 4c 49 44 46 4c 4a 4c 4d 4f 44 46 49 50 4c 4a 43 4a 4c 4c 4b 44 3e 44 46 3d 3c 3b 2e 30 27 14 0c 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1d 21 1d 3a 39 3d 3f 3a 3a 3b 43 41 3f 42 3f 41 3e 41 43 40 41 43 45 3f 41 45 45 4a 46 4c 4d 3f 4a 4a 4f 5c 52 4f 4f 4f 55 52 50 56 57 4d 56 47 5f 55 52 57 52 4f 58 4f 4c 5a 54 55 54 5d 57 54 5a 56 55 58 5a 5c 5a 55 54 5b 61 63 61 5e 5d 5c 60 61 58 62 58 61 5f 61 5b 5d 5b 56 62 61 5d 5f 60 5f 59 57 5b 5a 51 51 54 51 3f 16 05 06 05 03 00 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 0a 12 30 62 65 71 66 64 6b 65 64 6d 69 6a 6d 73 6c 6f 65 70 66 62 66 69 65 65 64 64 66 63 66 6a 5f 5e 59 58 54 52 51 59 54 55 58 5b 59 5b 51 5a 5e 58 59 58 54 4e 54 4e 45 4e 49 44 3e 42 48 42 47 47 49 4c 4e 54 49 4a 4c 46 43 47 5a 46 48 45 4f 48 42 46 41 42 35 2c 24 1f 0e 13 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 13 20 25 2b 3d 3b 44 3a 3e 3a 3d 47 43 42 43 35 3e 41 4e 40 4b 48 44 40 3d 49 45 44 46 48 46 4b 45 3e 4e 51 45 4b 4b 4d 52 47 4c 55 51 57 59 52 4f 55 4b 52 52 4d 5b 52 50 58 48 58 53 50 54 50 5b 60 58 5c 58 5d 5b 55 5d 5c 5c 5b 5a 59 5b 5c 54 5c 59 5c 5e 5f 57 5e 60 58 5f 59 66 63 66 59 5f 5a 58 60 5f 5a 4e 55 55 54 46 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 06 0c 2a 58 72 65 6b 56 5e 64 61 63 66 6e 6d 6e 70 6d 67 64 6b 6b 64 65 61 64 67 62 5d 58 5b 5f 5c 61 5c 55 58 5f 57 5b 50 55 54 59 52 55 54 4a 5b 55 61 55 58 59 4c 51 45 4b 4a 43 41 3f 3f 45 4a 46 47 4d 51 4c 50 4c 4d 41 44 4d 4f 52 50 4b 4e 41 41 3d 39 37 3e 2c 21 1b 0f 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0f 17 24 2a 2f 37 3e 3c 3a 42 40 42 47 47 47 44 41 40 3f 3a 45 42 42 41 3a 39 4a 3e 41 46 43 41 43 48 4b 46 4d 48 49 46 4a 4c 52 4d 50 47 56 54 4d 4f 51 4a 51 4d 52 47 4d 54 5c 58 54 57 51 4e 4a 57 54 55 5c 51 4f 57 51 4f 52 56 52 56 56 54 60 60 5b 59 57 5a 5c 5c 58 5f 56 5a 5b 61 64 60 62 59 5d 5b 5e 5e 54 57 50 5c 45 14 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 06 03 0d 09 21 52 62 6c 6e 65 60 69 5f 67 67 68 69 6b 6c 66 62 69 61 64 5e 5c 64 5d 64 61 59 57 63 56 60 59 53 58 53 56 54 51 55 57 55 54 49 48 55 4f 53 50 58 54 4c 58 50 43 4b 43 44 41 43 40 3b 47 48 4c 4d 4e 44 43 4e 46 49 4a 4a 48 4a 3e 4b 46 4e 49 44 48 3e 3e 3e 2a 25 17 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 06 12 11 14 30 2e 34 3f 39 3a 40 45 45 43 39 42 40 3e 43 40 43 3d 4b 3f 42 47 44 3e 41 4b 4a 46 4e 3e 4d 4b 4a 49 4a 46 47 4d 4c 50 56 51 5a 4f 4f 51 59 4f 49 4f 51 51 4d 50 54 53 50 4d 4f 4c 52 51 56 56 58 59 4f 54 50 54 57 55 5c 50 53 52 50 56 58 57 51 54 58 5b 51 63 5a 57 62 5a 5c 57 67 5b 65 5e 58 59 5b 62 58 5f 56 48 1d 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 03 00 06 05 06 00 0f 21 52 5e 66 68 59 64 65 64 57 5d 64 6b 6d 69 69 5b 61 66 61 60 57 65 5e 5f 5f 5e 57 5c 5d 5a 5b 52 55 58 5c 56 48 5d 56 53 55 4f 4a 5b 55 51 55 56 4a 49 50 45 44 4a 3e 45 48 44 43 43 4a 46 4a 47 46 4c 43 40 4e 51 49 4a 4a 50 4b 48 48 45 47 44 4a 3b 41 2e 2c 1b 16 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0b 1d 20 39 38 36 42 41 3e 3c 42 40 41 41 3a 3e 3b 39 48 43 45 44 37 3b 42 40 4c 47 4a 49 43 4c 4e 4e 50 4b 46 4a 50 4d 49 53 55 59 52 50 59 5c 56 5e 53 52 50 53 55 4e 4a 4d 50 51 48 4d 4f 52 55 4e 51 4e 4b 58 4a 55 4b 51 54 52 53 54 53 53 57 52 5c 58 58 57 59 5b 53 56 5d 5b 65 64 55 65 62 61 66 62 65 60 59 5d 5c 4f 17 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 20 4d 64 66 68 5a 5f 61 60 62 60 5d 67 6e 64 65 63 60 5f 5a 5e 60 65 52 68 55 61 5a 61 5c 5e 5d 5d 59 4f 55 59 51 50 4f 4f 4e 51 4f 53 57 58 5d 4c 51 4a 43 4a 47 4b 38 40 4f 44 46 3f 4a 4c 49 43 49 47 4d 49 44 4a 4b 42 4c 53 40 49 4c 45 48 3d 45 42 40 2f 25 16 12 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 08 12 21 2c 2d 37 3e 3c 39 3b 43 3f 3d 39 42 44 3d 36 39 41 42 44 3f 3d 43 47 41 44 48 3c 42 41 41 47 48 4e 48 47 42 3f 41 4f 53 47 55 4f 51 5c 55 57 59 54 5b 55 46 56 50 4e 47 4a 4d 47 47 48 4a 47 52 50 52 53 49 53 4f 49 53 4f 4f 58 58 52 54 52 56 50 5d 54 53 5a 5e 5b 62 5c 63 5f 69 5f 67 6b 6a 5f 5a 65 65 64 60 4b 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 4b 59 64 69 59 5f 5f 61 57 61 62 67 62 61 63 5b 62 64 61 66 58 5f 58 60 5e 5b 5a 54 56 55 56 55 4b 54 4f 50 53 50 4d 51 5d 4f 53 57 50 52 4c 44 3f 43 4d 4f 47 41 3e 3f 43 43 3e 45 42 46 44 44 49 44 4f 4a 43 45 4a 4e 4c 40 4a 44 3d 4a 4a 45 4b 43 3d 2a 1f 15 0c 05 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0c 15 21 25 39 3a 3b 37 3e 3e 45 46 3b 41 39 45 3c 3a 3d 4a 41 43 41 40 45 44 40 41 45 44 42 47 46 4b 47 4e 48 41 44 46 4d 49 42 4d 3d 4a 4d 50 5c 58 59 55 57 51 49 4f 51 4c 48 4b 4a 49 44 48 4e 54 58 56 4e 4d 4a 4a 54 50 4d 50 4e 53 55 52 49 56 58 4d 57 56 58 51 55 5d 61 65 67 70 6b 73 65 6e 64 6b 68 66 67 6b 6e 55 1e 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 15 46 57 5e 57 54 60 61 58 56 52 5f 5d 59 62 58 5c 5b 60 62 62 5d 5b 57 66 56 5b 54 5c 51 53 50 60 58 52 58 47 52 52 53 57 56 56 50 54 53 4d 4b 49 3f 44 40 48 44 46 49 44 44 3e 43 49 41 47 42 45 4b 3e 4a 42 48 46 52 45 46 46 4a 41 4c 4e 4a 4b 40 42 30 25 1b 0e 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 0a 1b 26 38 3b 44 41 3e 3e 43 3f 39 40 48 42 40 44 3b 3a 41 41 42 3f 45 3e 43 46 45 40 45 45 4c 4a 4e 45 49 44 4d 44 3b 47 41 46 4a 4a 48 51 4c 45 54 53 55 52 55 50 53 47 51 4e 53 46 47 4b 45 53 4a 4d 4b 4d 48 4f 4e 49 4b 49 4f 4e 52 50 55 52 52 52 56 4f 5b 52 5a 5e 5d 62 67 66 64 6b 6e 6d 67 6c 65 71 66 75 68 57 25 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0d 43 60 57 55 54 56 58 51 56 55 5b 5b 5c 5e 61 60 62 5f 5c 61 5e 59 5b 5a 5a 5c 59 51 59 59 55 54 58 4d 4a 55 51 55 55 4e 52 51 4e 4d 4e 4f 4d 45 3e 42 47 48 49 4e 42 45 4f 4e 4a 3e 3e 44 46 46 48 45 49 46 4b 5b 49 43 44 4a 49 4d 40 4d 48 43 4c 36 34 1c 17 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 14 1e 30 38 38 48 40 39 44 40 3e 3f 3b 45 3b 3b 3d 46 40 40 3d 3e 42 42 40 42 3f 44 3c 40 40 4d 44 45 48 41 46 48 40 4c 44 47 4b 48 43 38 4d 47 47 49 4b 51 51 47 4e 4d 4a 4e 44 46 3f 4a 54 50 52 4f 45 45 56 4f 50 47 4b 50 55 53 4e 4a 51 4f 54 52 51 56 53 4e 56 58 57 58 5e 5b 5f 60 67 6b 68 5d 63 60 60 5e 66 56 15 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 15 3a 55 56 54 51 56 57 4d 57 50 52 5a 55 57 5c 54 52 5f 5e 5d 4d 61 50 5c 51 53 4f 4d 48 50 56 4f 51 52 52 4e 4a 57 49 45 59 4b 48 50 46 46 44 46 4b 3f 44 41 47 4a 4a 45 43 4a 46 46 40 43 41 45 48 4b 46 46 48 3e 4a 43 43 4c 46 42 47 46 4f 45 3d 36 29 21 10 08 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 1c 36 38 38 43 33 41 3c 3f 3d 3a 3d 39 40 47 36 3d 3c 3d 43 39 41 3f 39 40 45 42 47 48 48 44 4b 45 3e 46 3f 41 44 40 4a 41 43 45 41 43 45 47 4c 4c 4e 40 50 45 49 50 4b 48 46 40 4c 45 4b 4b 3f 4f 4e 4a 49 4d 44 43 46 49 4c 54 43 4b 49 4d 49 4b 4e 4c 4d 4e 57 52 4c 55 55 56 5b 56 57 59 55 5e 52 4f 59 59 47 1e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 36 4e 4c 50 54 54 51 4f 4a 58 50 53 4f 53 53 53 54 59 5d 56 59 58 52 50 52 4f 49 4f 46 56 4c 4c 4d 4a 4c 4b 4f 45 49 4b 4d 50 42 43 40 46 43 3d 4d 3d 48 4d 40 47 40 48 43 45 40 40 43 4a 42 43 44 4a 45 48 42 42 41 43 45 48 45 46 3a 41 3b 39 37 27 27 14 0b 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 10 1b 30 35 38 3e 3c 3e 3a 42 41 3c 3f 46 41 35 40 40 39 40 42 42 49 40 43 44 45 3d 43 43 44 3f 47 47 4d 4b 49 47 47 45 46 42 46 49 40 40 43 49 4b 45 47 44 49 52 46 55 4e 4e 4a 41 45 47 4e 4c 42 47 4a 49 50 47 47 4e 4a 47 50 4d 45 46 4b 4e 4b 50 4c 4d 4b 56 50 50 52 58 55 55 4f 51 48 57 54 52 53 4b 4f 4a 45 1c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 35 44 4f 51 50 50 4f 43 53 4b 57 56 4e 56 59 52 58 5a 52 5b 56 50 55 50 4f 4e 4b 4d 48 48 48 4a 49 4d 4d 4f 4d 44 52 44 47 4d 45 44 41 48 45 4a 44 49 48 3e 46 49 40 4b 44 41 48 45 4a 45 44 4a 45 48 44 44 44 49 3c 47 49 40 49 43 3d 42 42 3f 34 24 26 15 06 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0f 1a 23 2d 37 40 3e 42 40 3e 39 3a 42 3b 34 3c 3b 3f 42 3f 3b 3b 40 3e 44 41 46 40 46 46 44 46 49 3a 45 45 47 42 45 45 41 3d 3d 3e 49 42 46 43 41 44 44 45 43 46 48 4b 4f 55 4c 40 3c 48 4a 41 46 49 45 49 46 50 48 4c 4c 48 4a 47 4b 4f 4b 4d 48 48 4c 4a 52 50 50 4e 55 56 52 4c 56 4e 51 4d 4c 44 48 43 46 40 40 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 31 44 51 57 4d 51 52 4f 50 4f 4c 4d 4d 58 4d 50 59 59 55 52 4d 57 4c 53 4d 46 4b 45 44 48 48 43 46 47 47 4e 50 51 48 45 48 46 40 40 44 42 48 4a 42 4a 3a 42 40 47 41 4c 3e 43 45 43 43 44 4a 4c 48 44 45 49 45 42 47 4b 44 44 46 49 41 3c 3a 32 34 27 17 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 1c 2a 2f 38 3f 45 44 41 44 39 39 44 37 35 41 3d 40 39 3c 36 36 45 44 3a 48 40 44 40 45 44 41 3b 42 45 46 37 45 40 54 40 3f 49 50 44 40 3c 43 3d 45 47 3d 42 42 49 4b 53 3a 48 44 4d 4d 41 41 42 4f 43 42 44 49 51 4c 47 4c 4a 4f 44 50 4f 49 49 50 44 51 4c 51 55 52 51 53 50 4a 50 4c 4a 4c 44 45 41 3e 47 3a 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 29 45 50 4e 3f 52 4a 46 4f 50 4d 4e 45 4a 50 52 56 50 55 5a 52 4b 46 4f 48 4f 52 4c 4e 4b 4e 46 55 46 4d 52 4e 4f 49 46 43 42 47 46 37 39 3e 3a 45 3a 48 45 41 48 4c 47 40 3e 3b 45 40 46 49 44 48 43 45 47 3d 40 40 3d 46 46 44 49 38 3c 35 30 2c 1e 1a 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0d 08 14 21 32 39 45 47 47 44 40 3d 46 44 3f 3b 3f 3a 41 41 3b 41 3f 3f 3f 41 46 38 38 3a 44 40 46 43 44 42 46 42 51 43 41 4d 48 3f 45 47 49 45 47 3c 4c 44 4a 42 3b 47 46 46 4c 4a 4b 4e 4f 4b 46 3d 47 3d 47 4c 46 4b 44 4b 4a 44 4d 48 4c 4b 4d 4e 52 48 59 52 4d 51 4c 56 4e 52 46 4d 48 49 46 4e 46 4e 44 3b 3a 1c 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 32 50 45 48 46 4e 4e 48 4a 4a 4b 52 48 49 4c 50 52 4d 47 54 4e 57 4a 4c 4e 4b 4a 51 4d 4a 4d 4a 4a 4b 4a 4e 48 46 45 48 3f 3e 44 46 40 42 48 40 40 36 47 42 3c 3e 3f 49 4b 44 49 46 44 45 48 42 43 4c 49 4a 41 42 41 45 3c 40 43 40 3d 3d 2d 2c 28 16 0d 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 10 1f 27 2d 41 4c 48 42 44 3e 3d 3c 43 44 39 42 43 3a 3b 37 42 40 47 3c 40 3d 3a 44 3c 3f 49 45 43 42 3a 3c 49 43 4a 44 49 44 47 49 43 49 45 40 41 3d 44 44 44 46 3f 40 4f 4f 4c 52 4a 4d 4a 47 48 4b 3f 42 45 4e 4b 4b 4e 40 4a 48 46 50 4b 4d 4e 42 51 54 56 45 4f 53 4c 4f 4a 47 48 42 4d 4b 45 40 3f 42 3c 1a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2a 3e 41 4b 47 4e 4b 46 45 4f 44 4d 4b 4f 4c 4d 55 4f 4c 53 52 4f 48 4f 50 54 51 4e 4c 4e 4d 48 47 4d 4d 4c 48 44 3f 41 3d 41 3f 43 3e 3d 49 46 43 41 47 40 3f 43 40 40 4a 41 42 41 45 46 3e 48 48 42 46 41 46 41 44 42 40 4a 43 45 34 2f 31 2a 1b 17 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 0a 06 16 25 2b 3f 3d 3b 44 40 3c 45 39 42 33 36 3f 39 49 3f 3e 36 39 3a 3b 40 39 3d 3a 42 38 48 3b 44 3c 39 3d 3e 3e 42 48 40 43 41 3a 4d 42 44 45 49 3e 45 41 45 44 42 39 4e 3f 45 4a 4d 46 45 4e 49 51 40 43 4b 48 4a 46 41 42 45 49 45 50 47 4e 4a 47 50 4b 49 4c 4c 52 50 4b 44 47 4e 4d 4e 4a 45 41 3e 47 2f 1b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 21 44 3b 51 3f 46 42 41 48 45 48 4b 4b 43 4a 45 48 48 45 54 4c 50 4e 4a 55 4b 4e 4e 4c 4f 4f 48 4c 47 4a 52 47 40 44 48 39 3d 44 45 41 41 45 3f 41 3f 49 44 3f 40 3e 46 41 45 4d 48 41 44 50 45 4a 47 44 45 38 3f 3e 3b 41 3c 33 40 2b 2c 30 25 1a 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 07 0a 12 20 23 31 3e 39 44 3e 3d 44 3f 49 36 3e 3d 3c 44 43 38 36 44 39 37 3b 38 47 41 47 36 3d 3e 41 44 41 3a 44 48 43 4b 44 45 47 48 47 47 41 41 44 47 42 40 4c 49 41 42 3f 46 49 4f 44 4b 4d 45 4d 42 46 4b 4e 51 47 48 42 4a 47 44 48 4e 4c 4e 4c 4b 55 52 4a 4b 50 4d 4b 4a 54 58 55 48 4a 49 45 45 41 40 3c 20 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 24 42 43 44 41 46 4a 47 46 45 4d 4a 4e 49 43 4d 43 46 46 49 47 4b 4b 54 4d 4e 4b 4a 54 52 49 51 4f 45 49 48 43 3a 41 43 4c 47 44 43 42 40 4b 4f 46 43 3b 44 43 40 3f 47 44 41 48 3e 3f 49 48 40 43 4b 3c 48 43 47 40 41 3f 42 37 3c 32 2d 2d 1f 17 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0c 1b 26 29 34 38 3a 41 43 40 33 36 3d 3f 3e 3e 35 3d 3a 42 39 48 3b 43 41 41 41 38 3e 40 3c 40 44 3e 3a 42 3d 3d 3f 45 45 3e 45 46 46 41 4b 3e 40 46 47 45 45 44 44 43 40 3d 49 47 50 4a 45 45 48 4a 52 4d 4f 4b 4f 4c 49 48 46 46 4c 44 4c 53 4b 4d 4d 4b 48 4a 4f 56 4f 53 54 4b 4e 44 41 3f 3f 38 36 3e 18 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 19 3c 3f 44 43 43 4b 3d 43 45 3e 4f 47 42 3f 4b 45 45 43 45 4a 4c 47 48 4c 50 4b 49 54 53 4f 54 4a 4a 45 4b 41 43 39 46 44 3c 3e 45 43 3a 40 42 3d 3d 4b 47 46 3f 40 45 40 41 4a 44 3b 3a 49 46 48 3f 44 47 36 41 3a 3a 3e 44 3c 3e 2a 2b 1a 14 17 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 19 29 2d 30 3a 41 42 38 43 3f 40 36 42 3f 36 38 41 43 3c 3b 43 47 3a 3d 3b 36 3c 39 3d 3f 39 3a 45 3a 46 44 40 3e 44 44 41 45 47 47 45 41 3a 48 4a 45 50 4a 40 40 44 45 47 4f 4e 3e 46 4a 4c 42 48 4a 49 51 52 4b 4b 49 3a 49 4c 47 49 48 4c 4b 49 4e 43 4c 46 4e 50 51 4b 4a 43 45 42 3e 3e 3c 38 38 15 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 20 39 3e 3a 3f 41 41 42 42 3e 48 3d 47 48 41 40 40 3e 44 3e 49 41 48 52 50 55 4c 51 52 45 52 4c 3f 41 3f 3b 38 3d 3c 3c 3d 3d 3f 3e 42 45 45 3a 44 46 47 3d 45 4a 3c 4d 4a 45 46 4d 47 45 45 40 46 40 42 41 38 3e 3f 40 3a 37 34 31 30 20 22 0f 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 13 20 2f 2d 36 40 3c 41 3e 3f 42 3a 39 2f 35 35 37 3f 43 3e 3e 41 47 3c 43 42 3b 41 46 33 3d 39 3f 44 44 3b 46 44 48 42 3f 43 43 46 45 47 3f 43 47 40 49 42 42 40 43 41 4e 38 23 32 4f 4c 48 44 41 4b 4e 54 4f 47 40 44 42 45 4e 46 4d 45 40 43 47 43 4d 48 49 4f 54 56 41 41 49 3e 41 3d 37 3e 31 3a 21 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1e 34 43 46 40 3a 44 3d 3e 41 3d 45 3c 41 47 44 37 46 49 3f 42 49 49 4c 47 50 54 4a 49 4c 43 40 45 3a 45 3d 38 31 35 40 45 3b 3a 47 3f 41 48 46 48 46 48 44 43 42 42 4b 41 46 47 47 4b 42 43 40 3d 3a 45 3e 3e 3b 3e 44 3a 31 36 2e 25 21 19 0c 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0e 19 28 35 38 44 3a 3c 41 40 40 42 37 3c 3b 3e 3b 3b 3c 3d 39 3d 41 3e 41 3c 3c 3d 3b 3f 3d 3f 3f 42 3e 41 45 3e 4a 41 39 43 45 3b 48 42 47 4a 43 3d 4c 41 40 4a 3f 47 42 41 46 48 4c 44 41 46 48 49 50 4b 4c 4e 46 48 45 40 41 41 3f 4a 4d 4c 4a 4f 47 4e 52 50 46 4a 44 44 40 3e 3e 3d 34 36 3a 31 25 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 38 3b 40 38 40 43 34 40 3f 3b 44 3f 47 44 3b 3d 39 3c 39 40 49 4d 48 50 54 4f 46 45 4b 4e 44 37 3e 42 3e 3d 3d 45 48 40 41 43 3d 38 48 48 44 3f 44 3c 4f 3e 3f 47 50 3e 46 48 47 4a 43 4a 44 3b 3c 37 46 33 3d 2e 3f 38 37 3d 2f 24 1e 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0a 12 27 31 36 46 45 37 3e 3e 41 3e 41 3c 3b 35 3c 36 3b 2f 3b 3c 39 3f 38 3b 3c 38 3a 38 3d 46 39 3e 40 3d 3a 38 41 49 3b 3f 45 42 44 40 44 47 41 46 49 4a 41 47 42 3e 4d 45 3f 3b 3f 46 3a 43 46 40 4d 4c 4b 4d 43 4b 46 48 4d 48 44 43 48 46 43 4c 42 49 4c 47 4a 4d 39 43 3f 3b 3f 36 2e 39 30 30 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 2d 3c 47 39 3f 39 3e 38 3d 3a 43 38 41 3c 3b 3d 3e 41 41 41 4d 3f 4d 50 4d 49 44 39 41 3f 41 3f 3b 42 39 3b 39 3a 38 41 46 3a 40 35 42 47 47 42 42 43 44 40 3e 3f 48 3d 43 3e 43 3d 49 39 44 35 3d 3e 37 36 39 35 37 37 38 32 2c 19 15 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 05 06 0f 1e 24 34 3c 3f 3c 41 3a 41 38 3b 33 2f 3b 3e 42 39 3d 39 37 38 31 41 3f 37 3b 48 3a 43 3b 3f 3a 3b 3f 3c 3d 37 45 43 44 3c 3f 3f 4a 3a 41 3a 41 45 4c 40 3c 46 3c 43 45 45 3e 41 47 3f 3e 3f 44 40 4a 50 4e 47 46 3e 45 49 4e 48 4a 45 4b 42 49 4c 49 4d 53 4b 44 46 3b 3b 36 30 3c 39 2f 45 31 22 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 36 3d 3d 37 3e 3e 41 3c 3c 36 38 40 41 41 3d 41 44 45 40 43 43 40 46 48 45 3c 43 44 47 45 42 40 41 3f 3d 37 3a 3c 3a 33 42 42 44 3e 42 3f 3e 43 4a 40 44 4b 47 4c 41 43 46 44 45 3c 37 3f 42 3a 39 3e 3c 2f 3a 33 35 35 34 30 2a 20 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 07 17 1e 2d 2f 3b 43 39 37 3e 3a 38 35 33 41 3e 42 33 3b 38 37 3c 35 3c 3e 3d 37 41 3b 3e 3b 3f 45 3f 3d 3e 45 3e 3f 3e 43 40 45 3c 42 43 42 41 45 44 39 44 48 45 46 46 44 46 42 4f 45 3e 49 43 4c 50 43 49 47 44 44 51 45 3f 3d 4a 4e 4f 4d 4e 4c 4e 4c 4d 4d 3f 43 43 41 3b 40 38 3c 3c 37 37 3b 23 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 32 32 3f 3d 41 36 46 39 3d 3c 4e 3f 3c 42 44 3b 41 41 44 47 4b 49 4e 40 47 48 43 47 45 42 43 43 44 3e 3c 3c 34 3f 3c 3c 47 3e 3c 3d 46 3a 44 48 41 4e 44 40 46 42 45 3c 42 42 41 3e 3f 42 3b 41 3e 42 3d 34 3b 31 39 30 30 25 1e 15 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 13 15 2b 28 36 42 3a 3f 3a 41 35 3b 38 41 3a 3b 35 3a 3c 38 3b 34 40 3f 34 36 3c 3b 40 41 41 37 41 44 3d 3e 3f 3a 3a 43 39 49 43 40 45 44 41 42 49 4b 51 3e 38 40 3f 47 45 43 42 3e 41 42 41 4e 3e 3b 41 42 4b 46 4b 43 49 4d 45 42 42 45 42 47 4b 52 56 4a 4b 3b 42 3f 3e 32 41 40 3b 41 3a 23 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 2b 30 3b 3c 45 39 38 38 36 3a 40 3f 3f 3b 46 3d 41 45 49 45 49 47 47 40 46 39 46 4e 4c 50 4d 42 4f 43 39 40 3d 41 42 41 40 3d 45 45 3f 4a 45 3d 41 43 48 39 3c 3a 43 3d 3b 3d 3b 39 3d 37 3a 37 36 36 41 34 36 36 2e 35 2a 1d 22 0a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 0d 1d 2d 29 37 33 36 3a 3a 3b 3b 38 30 40 39 42 32 35 38 39 36 34 34 34 3a 3c 31 3d 3a 3b 3c 40 3e 40 41 37 3c 3b 3c 4d 3e 3a 45 40 42 49 42 4d 3e 3e 41 42 40 40 3f 4a 3f 40 46 47 3d 42 49 47 3c 47 3c 3b 46 3c 48 45 40 48 4c 50 47 48 49 51 46 45 4a 4a 4b 3f 45 41 47 43 3e 39 32 36 34 28 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 29 36 43 36 44 44 41 37 3d 40 40 4b 43 46 43 40 4c 40 44 43 45 4d 55 51 4a 47 40 4d 47 41 4b 51 5a 55 45 35 3d 4a 3c 3f 40 37 44 41 39 48 3c 46 42 43 45 39 45 41 41 3f 3f 45 3d 39 38 35 36 39 3e 2e 37 33 33 33 2b 24 23 27 19 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 08 11 10 1e 2a 37 2f 38 38 44 32 33 38 2f 38 3a 41 3d 3d 3b 38 38 36 33 3b 3e 38 3f 3b 3c 3d 3d 3a 3f 45 3e 3d 44 3e 3f 3b 39 44 46 40 4b 4c 45 45 41 43 42 48 3d 42 40 43 3f 3f 42 41 41 43 47 46 3e 45 48 44 44 43 4d 45 4a 44 4a 43 52 4a 46 42 4b 4a 4d 4d 4b 47 49 42 3c 41 45 48 40 3f 3b 23 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 2f 37 3f 38 39 3a 3c 42 44 46 3f 44 4b 43 45 3d 4a 44 4f 3f 46 5b 5c 52 4f 46 4e 4d 46 4d 52 57 59 50 50 43 50 43 47 48 43 47 43 4a 43 40 42 49 42 46 3c 3b 42 36 45 3f 3a 49 3b 31 34 36 45 41 40 37 35 2d 35 2f 2b 2a 1d 18 13 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 0a 1e 26 2d 32 2d 3e 3b 37 37 2f 39 38 3b 3b 36 3e 39 38 37 3f 33 33 43 39 3c 3e 3d 3a 3d 42 42 43 4b 49 44 3c 44 3c 37 3b 3b 38 42 40 46 41 3f 49 44 41 43 3c 42 49 47 49 48 4c 40 3f 42 42 42 4d 43 46 40 42 44 43 48 4a 47 43 4a 3e 47 43 42 43 47 47 44 46 48 45 44 43 3d 3e 41 4a 43 2e 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 27 3a 46 3f 3e 40 3f 49 3e 45 46 43 49 43 46 3c 45 40 45 44 44 5b 54 4d 42 3f 48 3e 4f 46 53 4f 52 52 4f 55 56 45 46 45 47 47 47 3f 3a 4a 45 44 47 42 3b 3f 41 3d 3c 3d 33 30 3d 37 46 34 3b 3a 3a 33 3c 30 29 26 25 2f 1b 15 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 14 1d 29 30 36 2f 3f 35 37 32 3a 38 35 3b 36 3d 3c 3b 38 32 39 42 3b 37 3b 37 40 3a 3c 3a 3a 49 4e 3b 3b 41 4a 3b 41 3e 44 39 43 40 41 43 3e 40 45 43 3e 3e 42 40 43 41 43 3e 3d 41 44 42 45 50 4c 46 44 43 47 48 44 4c 49 44 45 4c 42 42 42 45 48 44 48 37 42 3b 42 43 3e 38 3f 38 3c 32 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 2a 3c 40 40 3a 3e 41 40 4f 45 52 39 42 40 3e 3f 38 3b 39 3b 4b 49 45 45 43 3c 3a 38 39 47 40 42 44 49 4d 5b 50 4b 4d 46 41 43 44 47 45 45 44 42 3c 37 37 35 41 3b 3c 44 3d 3d 3f 33 33 31 36 3a 3e 39 37 35 2d 23 29 22 12 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 1d 22 2c 35 37 3b 37 39 3c 3a 37 39 33 30 39 3a 37 38 39 42 38 36 38 34 35 3b 39 3a 3c 45 43 3d 39 45 46 44 44 38 3e 47 3e 3b 45 3e 3e 43 41 46 40 41 3e 4b 43 44 3b 3c 40 3f 3e 45 47 48 54 54 52 57 42 4d 4b 49 4d 56 51 4d 4a 40 3a 44 3c 45 41 44 43 3f 40 43 3d 43 3e 43 3e 38 2b 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 40 48 3c 39 3d 3d 45 4c 48 44 3b 41 37 3e 3c 3b 41 35 3c 43 43 46 3f 4d 34 3a 3b 3e 43 44 3d 3c 47 47 4d 51 4f 4e 4b 4d 3f 4f 4d 4c 4f 47 42 46 44 47 3d 3b 3c 44 40 34 39 39 34 3b 38 3e 41 43 3a 40 2f 27 2b 1a 0e 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 09 1d 21 31 30 34 41 43 3a 37 39 3b 31 39 37 36 39 32 35 3f 42 44 34 37 3c 3d 37 38 3b 42 3a 44 44 41 44 44 44 41 41 45 3b 42 44 3c 40 3f 3e 46 44 4a 49 44 41 43 44 3c 3d 3c 3f 45 46 44 53 61 5e 61 4b 50 4b 4a 4d 52 45 52 43 49 40 47 45 44 49 40 39 36 3b 39 3e 40 43 47 3f 40 33 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 25 3c 42 3c 39 41 43 40 45 3b 41 3a 3e 42 3c 3a 37 3c 42 37 3a 42 3d 3a 42 3a 3c 38 3f 39 43 35 41 43 40 46 46 44 4c 45 4b 53 4f 4e 48 4c 47 3c 42 41 3f 40 3e 3b 37 40 3c 3c 3b 35 45 42 3b 45 3e 32 35 2b 28 20 20 10 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 10 21 27 30 39 3d 45 37 38 35 38 33 30 34 39 3a 37 3a 35 31 3c 33 36 34 37 38 3b 3d 45 3e 3c 3f 3f 3f 3c 3b 3a 47 46 3f 42 43 3c 39 3e 36 3f 3c 44 3d 40 3e 3c 3d 3f 3c 44 3f 46 42 42 4c 57 53 59 52 4b 46 41 49 45 49 47 40 40 43 44 4b 40 44 47 48 3b 40 36 46 37 40 46 43 34 2a 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 20 31 43 35 3c 38 41 41 3c 41 3e 41 41 39 3f 3e 38 37 37 35 3a 38 36 3c 3b 30 40 39 38 33 39 38 3a 3e 40 3d 40 4b 43 46 46 4f 4f 4a 46 3d 4f 3f 3a 40 43 38 3b 3b 42 42 3d 3a 36 3a 38 46 44 3e 3c 31 2b 1e 1f 1a 11 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 1b 1a 27 35 3e 43 48 3e 3b 3c 36 33 3b 3d 31 34 35 2d 37 3a 32 35 33 36 3c 34 3e 36 39 39 39 3d 3d 39 3c 3b 45 42 44 3f 40 3d 3f 3d 44 3f 3f 43 44 39 44 45 44 46 36 40 42 43 44 45 4e 4f 47 4c 52 48 4f 3f 47 46 47 43 3f 39 3f 4e 48 47 4b 45 42 43 3b 37 42 3d 43 49 40 3b 28 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 27 43 42 39 39 48 3d 40 42 43 3d 3e 37 39 41 37 39 39 38 37 38 31 36 33 33 3c 2f 3a 34 41 3f 31 39 37 44 3a 3b 47 44 47 44 51 51 54 4d 44 44 43 40 3e 3e 3d 48 3f 43 3c 36 3f 39 3a 45 44 40 43 3f 31 2d 1d 1a 17 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0e 29 28 32 3a 38 39 3f 3b 41 33 31 3e 34 3b 3d 32 36 35 3c 32 3e 37 36 37 3b 3e 46 33 39 39 3c 41 43 40 3d 3e 3c 3a 45 3d 3e 43 40 47 3f 3d 39 3d 47 3e 42 49 3c 44 3d 3c 3c 42 4d 43 4c 41 44 49 41 42 47 3f 44 43 4b 42 42 3f 38 45 41 44 4a 43 47 40 41 3e 3d 3b 40 37 3b 25 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 2b 42 41 3d 40 37 3c 3e 40 3c 35 2f 3e 34 3c 38 3f 3d 3f 36 3a 34 38 31 3b 37 36 3b 37 39 34 3b 3f 36 3e 3e 42 4e 43 42 4b 47 4a 47 42 45 46 41 3d 3b 3f 36 3e 41 3c 38 35 3d 3d 42 4b 44 3e 36 3f 31 28 1c 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 11 0f 0e 1a 22 31 2e 3a 32 36 3b 32 33 2e 34 2e 2e 36 35 3c 33 3c 36 3b 3c 35 38 35 30 3d 40 39 39 37 39 49 36 43 3e 40 39 3c 43 3d 42 44 3f 3b 3b 39 3c 40 39 3e 3f 3a 3c 3c 3e 43 4b 4b 44 42 3c 3e 3d 3b 38 3f 3e 3e 47 3a 39 37 3b 36 4b 4b 4c 41 43 41 41 42 3e 43 3a 33 38 36 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 44 49 4a 44 3a 3f 3e 3b 32 3d 3b 30 39 35 3b 3d 33 35 30 39 3b 34 3a 3a 35 31 34 36 35 3d 31 2f 3c 3c 3e 3b 46 48 4c 41 4a 46 40 46 44 40 41 46 3a 3c 3c 3a 34 41 37 41 3e 3a 42 43 3a 38 26 2a 28 1d 12 10 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 0a 1c 2c 2b 32 2d 35 36 38 2f 32 39 34 3b 39 34 32 39 33 3c 3a 34 37 3a 35 34 41 3a 34 3d 3e 3d 3c 3e 3e 42 3c 37 45 3f 42 42 3b 46 4a 3d 3f 48 40 44 3e 41 42 42 3d 49 4a 41 42 46 3f 45 43 40 46 3f 43 43 3d 41 46 3b 41 41 42 40 49 49 4e 51 46 48 41 3f 3b 38 3d 45 3a 33 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 3b 3e 3b 45 3e 39 3b 36 3a 3c 3e 40 33 3d 3b 37 37 35 38 3c 36 3b 39 3e 37 36 37 3f 3a 36 2e 3a 38 36 42 3e 4e 4c 4e 4f 40 44 46 3f 45 48 44 42 41 38 3e 44 3d 44 3a 34 46 44 3e 37 30 30 3a 2a 1f 16 11 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1f 1e 25 27 2e 2e 2d 35 34 2e 32 32 35 35 34 38 39 35 3b 35 3d 34 39 33 3e 3d 38 3c 41 38 45 39 39 3b 48 35 38 48 3f 43 4d 3e 4d 44 40 3a 40 48 3c 4a 45 3d 41 3d 44 47 43 45 41 3d 40 3d 48 40 42 44 38 42 43 3d 39 40 40 41 4d 46 5a 58 4e 49 42 3d 35 39 33 42 3d 3a 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 39 42 40 3e 45 3c 3e 3a 3a 39 36 3a 3a 3d 39 34 33 39 32 3c 36 3b 3b 3b 3b 36 40 40 3a 40 35 36 40 3e 39 37 44 45 46 48 43 3d 4d 4a 48 49 41 3c 43 41 30 47 3f 40 41 37 3a 3e 37 34 30 31 2c 23 1d 0e 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 15 0f 25 24 2d 2a 26 30 2b 2d 2a 28 2a 32 36 34 3b 30 32 32 3c 3b 36 31 38 39 3a 3a 3a 3e 42 40 3d 3c 3b 3e 31 45 3c 3f 3c 42 44 43 42 3e 47 41 39 41 41 41 4c 42 40 44 41 45 42 48 3f 3d 45 45 44 3c 41 44 3d 3e 3f 40 40 3e 41 45 48 53 55 52 4c 42 3d 3f 42 3b 44 40 38 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 36 42 3c 3a 45 36 37 42 36 39 3c 37 40 38 35 39 38 3a 2b 31 3a 3f 32 3d 37 35 39 34 36 38 33 35 37 3e 40 3c 40 4c 45 4f 49 45 43 4d 51 4d 4d 41 3e 43 3c 3c 42 41 41 38 3e 35 2f 37 2f 28 24 1c 1d 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 17 18 23 20 26 28 2b 2d 30 31 33 32 2e 2b 32 38 3a 36 2d 30 35 36 37 37 36 3a 31 3b 38 3f 40 3b 3b 33 42 38 45 3b 35 35 38 36 3f 3b 3e 38 41 40 3c 43 41 48 48 45 44 43 38 4b 3c 47 4a 47 45 46 44 3f 44 45 3c 42 41 49 46 47 46 47 4c 4f 4c 4a 42 51 4a 44 3e 41 41 3f 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 33 3f 31 36 36 39 3d 39 38 44 38 36 2f 36 37 37 2f 38 37 3c 34 3b 35 38 36 3c 3b 3b 36 3e 34 34 42 3e 41 3c 47 44 45 47 44 48 44 46 4e 49 4e 41 43 45 40 3a 3d 3e 3d 39 3e 36 2f 31 2a 23 29 1d 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 14 1c 20 23 2a 29 2d 2f 36 31 30 31 39 35 34 31 3c 39 33 30 34 35 38 38 38 3a 40 37 38 3f 42 39 3d 3b 3d 3b 3e 3c 39 3e 39 43 3c 3a 3e 3f 44 3d 3e 45 47 41 42 43 49 4a 47 45 50 45 41 4c 4c 51 4a 4f 50 4e 46 49 51 4d 4f 4f 4a 51 4d 49 4d 4f 48 44 3d 41 3b 41 41 20 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 29 3f 32 36 31 33 3a 3e 36 3c 33 30 39 3b 42 34 3e 3d 34 34 34 40 3f 3c 39 36 36 38 3b 3d 37 35 42 3f 38 41 3f 4a 4d 4a 4c 45 43 51 48 54 4a 4a 41 44 40 44 47 46 45 47 36 36 2f 30 29 27 12 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0b 19 1b 23 25 25 2b 39 35 30 39 2f 32 39 3b 32 38 3b 32 34 3b 34 3c 3d 3b 39 3b 37 37 3d 43 3d 39 41 3d 40 36 34 44 3b 40 3e 36 41 3e 3d 41 44 3c 43 3e 46 42 47 50 44 47 48 4a 4f 52 5b 52 5f 5d 5b 66 5b 64 6b 61 61 5b 5d 61 5f 59 55 54 5a 54 50 4b 3b 46 40 36 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 2c 37 3d 39 3f 3c 35 3f 37 3d 31 34 36 39 3d 37 3f 36 3b 41 38 3a 38 41 3b 36 3d 35 39 3a 33 34 33 37 41 47 41 4b 47 44 47 45 4e 4f 4e 50 46 50 4b 49 46 4b 40 47 3f 39 39 2d 2d 27 22 17 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0e 13 19 20 29 32 31 2d 3d 2a 2b 37 29 36 34 30 33 38 2e 37 37 33 39 36 3f 31 3f 3d 41 39 3e 42 3b 3c 3c 41 3b 3f 3c 32 3d 38 3b 3e 40 41 3e 44 46 46 48 4a 4e 54 52 63 62 62 6e 67 6c 68 6b 68 6e 72 74 73 72 76 6f 76 76 6d 6b 6c 66 6b 5f 5e 50 50 4b 45 41 32 28 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 25 2f 35 35 3a 3b 37 38 3f 37 3c 38 42 38 35 37 35 3d 42 41 35 35 39 3a 36 35 38 41 39 34 39 35 42 3c 3e 3a 42 48 46 46 51 4f 4e 45 4c 48 48 54 58 55 53 4e 49 53 41 41 36 2f 2a 27 1a 10 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 10 15 23 25 27 32 34 3b 38 36 2f 34 33 38 39 37 35 35 37 36 35 3a 3d 3c 34 44 3a 43 3e 37 44 3f 36 3e 3b 39 42 38 3d 46 33 3e 43 41 47 4a 4a 48 4e 4d 61 63 67 6b 6e 6d 6a 79 7b 76 7e 7c 77 7e 71 7d 7f 75 79 83 85 7c 7c 82 7d 79 77 79 75 70 67 5b 59 54 46 35 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 2f 35 2e 39 39 37 3f 36 47 43 3d 38 2f 31 3c 33 3e 42 38 38 31 35 39 3d 40 38 38 38 38 38 39 35 37 38 3a 3e 4a 46 4d 45 45 49 4c 4f 54 4e 50 57 5b 50 55 4f 50 4e 46 40 39 36 28 26 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 19 1c 33 28 2d 36 31 29 2d 3a 31 3a 2b 31 31 36 2d 38 38 33 3a 37 3c 42 40 35 37 3e 36 39 3e 3d 40 3b 3c 38 36 3f 3f 42 47 49 41 53 56 5d 5c 67 70 6e 73 6e 7b 73 78 7d 7a 79 7f 7a 7c 81 7d 80 80 7a 82 7c 85 7d 7a 82 81 80 81 7c 75 7a 73 6c 70 64 58 33 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 26 3c 36 3d 38 3b 45 3d 3f 34 3b 36 32 39 3a 40 36 34 35 38 35 3c 43 2f 38 36 41 37 36 3d 31 3d 3c 35 3a 47 3e 4a 44 46 49 56 4e 4e 52 56 57 5b 54 5b 53 4c 55 51 52 46 3e 2c 24 1f 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0a 19 2b 28 2b 34 2f 39 33 2c 37 37 37 37 32 3b 2f 36 37 35 34 35 3a 3d 36 33 33 32 33 3e 3d 3b 40 2f 3c 3c 3d 3e 40 42 46 51 55 5d 6a 6e 6c 72 7e 75 79 7e 85 80 7a 7b 80 80 78 7d 7e 82 82 84 85 7d 84 7e 83 86 89 7d 81 81 80 7f 7d 72 7a 70 76 74 6e 43 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 28 38 3b 44 43 40 39 42 47 3d 3f 36 31 3b 34 43 36 3b 36 34 3e 3c 3b 3e 2f 38 37 34 30 3d 3f 3d 39 3c 43 41 41 3f 45 4b 49 54 51 50 55 54 5a 58 5e 60 59 59 54 59 52 4e 42 32 1d 0c 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0e 10 1d 2b 2b 37 30 31 36 34 3f 3b 37 35 33 3a 39 38 34 35 33 37 35 3e 39 34 3a 33 3c 3b 36 3b 3c 3b 3f 47 37 43 48 46 57 5c 62 66 6d 78 73 72 78 7b 7d 7b 76 79 87 7c 81 84 88 7e 7d 7e 82 82 82 7c 7f 79 8c 85 88 7e 7d 80 79 7f 7e 7c 72 78 7b 72 6a 49 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 2c 3b 3d 43 40 37 3e 43 3e 42 3a 3b 42 38 3b 3b 33 3a 38 35 41 38 3f 3c 37 3a 43 3f 47 45 43 38 44 45 42 3c 41 41 49 4e 4d 54 56 55 62 5a 5c 5a 63 61 64 5d 5d 5c 58 48 3f 2f 1f 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 11 1b 20 28 2a 35 37 2e 3f 39 42 33 32 2f 3e 35 3c 35 3c 2d 35 30 39 3c 32 3a 3a 36 44 3e 33 3b 3b 40 3b 41 45 48 5a 60 6f 7a 72 7c 7b 73 85 7c 7f 7f 7f 7a 83 86 80 75 78 7f 7b 80 7f 7b 7e 7d 74 83 77 7d 82 84 87 83 7c 74 7c 7c 7a 79 75 74 6d 6e 4f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 32 46 3e 47 41 44 43 3c 43 45 3b 3a 35 37 3a 3e 39 44 36 41 37 36 32 40 33 34 3d 39 3f 3a 3e 3e 47 46 44 41 41 49 40 4a 55 3c 62 5d 57 64 5a 5d 5f 6b 65 66 62 5c 51 4a 43 2e 12 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 19 21 2c 2f 2c 30 32 3b 33 32 38 34 38 32 30 38 36 36 3d 34 31 37 34 3e 3c 37 3b 40 3a 3a 31 3b 3c 45 50 52 5f 6c 6d 73 73 78 7f 7d 76 76 7b 7e 7f 7a 7b 7f 7a 79 81 82 7e 74 7d 74 7a 7a 6f 79 82 82 84 7f 78 7c 7a 7b 75 7a 79 78 70 70 6d 66 51 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 3b 43 40 41 3e 31 38 37 3f 42 3b 3a 39 3f 3e 3a 3a 33 36 3a 3d 3a 3e 3f 3f 45 37 42 3e 43 38 3c 45 3c 42 4e 42 44 4f 4d 56 5e 52 5a 5d 5e 5a 66 61 69 6d 67 60 62 54 4a 42 36 1b 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 15 19 21 2c 2b 35 35 31 35 3b 36 35 41 35 3a 34 3b 38 37 31 38 33 38 3d 40 36 36 39 41 3f 3c 38 3e 49 4d 61 6d 78 70 73 77 78 7f 7c 7b 80 7c 7a 7c 73 81 7f 78 76 78 7e 76 7a 7c 7b 7c 78 7d 76 7b 7a 78 74 7d 7c 7b 76 6f 72 7b 6f 70 7a 75 6e 4f 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 3f 58 50 41 43 33 40 36 30 3f 37 3b 3c 3a 3d 37 3e 3f 3b 44 3c 4a 40 4d 40 46 45 47 3e 42 45 42 46 44 42 49 4c 44 4d 49 57 55 55 62 61 6f 71 6a 77 72 73 76 66 5f 51 41 37 2d 21 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 13 24 2d 2c 35 2f 31 39 37 35 34 3c 31 35 34 38 34 3c 3b 33 33 34 39 37 36 3b 33 39 3e 3b 45 3e 4c 59 6a 76 7d 7c 77 79 7a 83 75 76 75 7b 76 75 79 7f 81 81 73 7a 78 78 74 7b 7d 76 7a 7b 75 74 82 75 7b 7c 7b 75 74 75 6b 6f 69 76 71 70 5c 55 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 3f 6a 5e 52 48 36 33 37 34 36 3b 3d 35 3c 3a 3d 40 45 42 46 47 4f 4f 52 59 49 54 54 49 44 3b 3e 41 3e 4d 4b 48 47 47 52 54 62 62 69 6e 6b 79 7e 80 82 7e 7b 6e 5c 57 3f 35 2a 22 1d 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 12 1b 23 28 29 33 30 3b 33 3a 35 2f 39 3d 37 31 3c 2f 2f 34 34 32 32 36 40 32 38 3d 31 3d 43 54 5d 6a 6b 6e 77 7d 72 72 79 73 71 79 75 76 6f 7d 75 75 7a 70 7a 77 76 6d 6e 74 75 74 75 7a 74 75 75 77 76 75 7d 73 73 67 70 6f 6b 6e 70 62 4f 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 43 63 60 60 51 3f 2e 34 31 34 36 39 39 36 43 40 40 4a 50 52 57 5c 5e 5f 58 60 57 51 49 3a 3f 3b 3a 3f 3c 41 4d 50 52 4f 55 5d 65 66 72 79 91 94 9d 96 92 83 6c 62 53 49 48 3b 2b 26 0b 08 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 16 0f 25 26 31 31 35 37 38 40 34 39 2d 2e 44 3b 3b 38 36 37 36 36 32 3b 37 3c 2c 37 3a 44 47 62 70 74 6b 73 72 73 70 75 7c 69 71 6e 69 6e 75 73 78 6f 78 70 78 6e 6f 7a 70 6f 76 77 75 71 6d 78 77 77 72 6e 72 6d 6b 70 71 69 6d 71 65 64 56 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 3d 64 62 64 50 47 34 36 38 41 35 41 36 41 4a 47 54 50 5d 5c 5d 6e 6f 73 65 69 65 56 51 49 39 41 33 44 41 44 4e 53 59 4b 5b 5c 69 75 8a 93 a4 bf c4 ca b5 9f 82 76 5d 4e 41 3e 2e 22 15 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0e 10 1d 28 2f 2d 38 35 38 3b 35 3a 31 2e 36 35 2f 3b 3a 38 36 36 3b 3d 36 3b 3b 40 3f 56 5c 67 6b 66 73 6f 71 72 76 75 72 73 72 75 7b 77 78 73 74 79 69 73 74 70 6d 75 6e 71 75 70 73 71 68 71 6f 71 74 75 73 6a 6f 64 66 6b 67 65 5b 4f 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 3a 64 60 66 48 44 3d 36 38 3c 3c 44 4f 4d 5b 56 61 6a 66 6f 70 6d 70 71 65 6b 65 56 54 45 3b 3b 3c 45 45 47 4b 4c 52 52 5c 60 6e 85 8e a8 cd d9 f3 fa e2 c0 a9 89 6e 56 49 44 34 30 26 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 17 1d 23 2b 2b 38 39 33 32 2d 34 2f 2d 29 32 3b 39 30 37 36 34 34 39 2d 3d 43 50 59 65 70 6b 6f 71 6f 70 78 76 6d 6c 71 70 75 74 6b 6d 6e 71 72 72 70 6c 6b 6a 71 72 6f 72 6d 67 73 63 71 6a 6d 6c 6c 6c 6b 6d 65 5f 62 69 58 5a 49 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 37 56 4b 5b 4a 37 32 38 3d 44 3f 41 4b 59 64 67 68 71 73 74 73 75 6a 65 67 60 5a 4d 4d 4c 39 3a 3b 41 42 47 43 51 5c 60 63 64 73 84 a6 c2 e4 ff ff ff ff f6 d2 ac 86 7b 54 48 42 3c 2f 18 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 11 1d 27 26 32 32 3a 2f 3a 33 36 36 3b 32 32 35 34 33 34 3e 2d 34 35 2a 40 47 54 60 65 6a 6f 73 77 6e 72 6d 6e 6f 74 6e 71 73 6a 6f 74 69 6d 73 6a 6d 66 64 6a 68 6e 68 6b 6d 6d 70 73 63 6e 64 69 6c 63 63 64 68 5e 64 5e 61 4f 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 31 4d 57 4f 41 35 32 35 47 47 50 53 61 5f 65 6d 6b 6c 6c 74 70 75 6d 63 63 4e 51 4d 4c 3f 3b 3d 37 39 40 48 55 58 62 59 5f 6a 6e 86 a8 d6 f4 ff ff ff ff ff ff d4 a4 75 5f 47 43 40 2d 1b 0d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0f 12 1e 25 2b 2f 31 38 37 34 36 2d 33 31 39 37 34 3b 37 34 38 3e 32 35 40 45 55 67 65 69 6d 6b 66 6e 6e 6e 72 6c 6f 6b 68 71 6f 6d 6e 62 72 65 6b 73 68 6a 71 71 68 65 6d 62 6c 67 64 63 63 6c 69 72 67 6a 62 5c 5f 5d 5a 5a 4d 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 28 4e 51 49 40 36 40 45 4f 52 5a 61 68 6c 6b 73 6b 70 67 64 5e 63 64 5c 5d 50 4a 51 40 3b 43 32 3b 3b 3c 4d 49 4f 5c 5f 61 6f 74 89 aa de ff ff ff ff ff ff ff ff cd 9d 78 5f 48 45 31 20 12 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 05 12 20 24 33 34 32 32 33 32 30 31 2e 3a 35 30 38 33 37 37 30 35 37 3f 43 58 57 63 6b 72 6e 6a 6a 70 6b 65 67 68 6c 6a 70 69 6b 66 66 6e 63 65 6a 65 65 6d 5e 67 72 62 67 69 67 67 61 6a 66 64 69 62 5e 64 5c 5b 5f 5d 55 4c 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1e 45 41 3e 42 40 45 4a 52 44 61 64 69 6e 66 6e 68 64 6b 6e 61 6c 5d 5c 53 4c 4e 45 41 3d 3a 36 2e 35 41 4c 52 4c 53 5a 67 6a 72 7f a5 cc ff ff ff ff ff ff ff ff ff b6 85 71 4e 47 3c 26 1a 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 12 16 26 2b 2e 2e 3a 2d 31 3a 35 34 32 34 39 34 3a 39 35 31 3e 42 48 4b 57 62 65 69 69 66 6a 67 66 6c 66 66 64 66 6a 63 67 65 67 6a 60 65 60 60 61 5d 64 65 65 65 69 5f 67 6c 62 63 68 5f 5d 5d 64 60 5a 62 5c 56 55 4f 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 42 42 46 3d 43 3b 47 51 63 5f 62 6a 67 6b 64 60 67 67 5f 62 5b 50 51 50 43 40 44 3b 2e 35 36 3a 34 3d 45 42 54 5e 61 64 65 70 77 8b b7 ef ff ff ff ff ff ff ff ff ec b1 83 61 49 31 28 1d 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 0a 17 21 2b 29 31 34 3a 3d 32 3a 32 31 3f 37 3b 3a 36 3a 36 37 4c 53 61 61 65 64 69 73 72 70 75 69 6c 65 66 69 60 61 66 61 67 61 5e 62 69 67 69 68 63 61 5e 66 5c 65 68 67 5e 65 66 64 5c 5e 65 5c 59 5c 60 60 59 4b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 15 3a 36 3b 44 3d 49 55 63 64 60 61 62 66 61 65 66 62 5c 59 52 5d 50 46 3f 39 40 32 36 36 39 35 34 34 45 3c 4d 53 53 50 62 67 65 6b 70 90 d1 ff ff ff ff ff ff ff ff ff d6 9b 73 58 3a 2d 23 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0d 1d 25 2a 2c 30 2f 37 34 39 36 39 2e 30 33 38 32 31 42 38 49 4e 55 58 5d 6c 6b 6b 71 66 65 6c 60 62 63 61 61 5c 66 61 60 60 62 66 62 66 66 5f 67 65 6a 5d 62 63 63 69 62 67 62 5e 61 5e 60 57 5e 53 62 5a 54 44 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 18 3b 35 38 36 38 4a 55 53 5b 5b 57 5a 60 4d 5a 5c 55 58 4a 4f 50 49 46 42 35 3c 35 35 37 35 36 35 3f 3a 2e 4b 4e 5b 54 54 5b 60 51 69 71 a6 ea ff ff ff ff ff ff ff ff ff b9 7f 61 3f 24 1a 0a 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0d 0e 11 25 24 35 32 32 31 36 3f 36 34 2d 36 3b 3b 3b 37 3e 44 4d 5d 63 61 67 66 6b 6b 6b 68 62 5e 63 62 5d 5f 60 5e 63 5e 5a 5a 62 5d 5c 59 56 5d 61 63 64 5f 60 5f 5f 66 63 6a 5f 5a 57 5a 58 4f 59 57 4f 4f 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 38 3a 41 35 32 43 48 45 50 50 56 55 57 57 52 53 50 45 46 44 44 46 3e 30 3b 2c 36 31 2f 3c 31 39 30 38 37 3e 44 4a 52 58 54 44 4b 4d 57 83 b5 ff ff ff ff ff ff ff ff ff d3 91 6f 4d 33 1c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 13 16 21 29 2f 2f 31 30 38 36 38 37 35 39 3b 32 3c 3c 42 52 57 58 63 65 6a 6b 65 6d 70 62 64 65 5d 66 55 60 5b 57 5a 55 5c 62 5e 5f 59 5b 5d 5d 64 61 5c 62 63 5e 6a 60 5f 57 54 5c 5a 58 5a 5d 55 5b 4c 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3d 32 32 3b 39 39 3d 42 43 4b 46 44 4c 4a 54 4a 48 44 3d 44 3b 3b 3a 32 36 35 39 36 39 3c 3a 39 36 38 39 3d 3c 47 47 49 44 48 44 47 5a 67 91 d8 ff ff ff ff ff ff ff ff f6 a7 75 4c 33 1e 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 1e 1b 24 2c 29 3b 33 31 39 30 35 33 3b 39 36 37 44 4a 54 53 5f 60 62 6d 6a 63 68 6a 66 64 64 5d 5b 5c 50 55 5c 58 55 54 56 59 5a 53 5d 56 58 60 62 58 5b 61 62 56 59 5c 5c 57 52 56 57 53 58 4f 48 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 35 30 2f 39 32 36 3d 36 3e 34 3e 42 44 47 45 44 36 39 38 35 37 30 36 35 32 34 2c 34 32 3b 32 38 3b 3d 3d 3b 31 36 32 31 37 35 36 45 4e 58 79 aa e5 ff ff ff ff ff ff ff ff b7 81 55 39 26 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 0d 1b 1e 2d 33 29 32 2e 3a 36 36 32 26 36 3a 45 41 40 52 52 5a 5e 62 65 63 60 6a 63 5d 60 5e 60 5b 5f 5b 50 53 53 56 4e 4d 4e 4d 4f 58 53 4b 52 5b 5f 53 5f 61 54 57 58 56 57 51 54 50 52 4e 42 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 2b 32 3b 34 31 25 2f 33 33 33 33 3b 37 34 3c 37 37 34 32 35 39 32 34 31 32 2d 38 34 36 38 36 3d 39 37 2a 22 23 20 21 25 2d 32 3a 39 46 57 62 84 b4 f1 ff ff ff ff ff ff ff c0 88 53 35 16 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 0f 1a 21 24 29 2a 31 39 33 32 33 32 36 40 3a 3e 3f 3d 4f 51 5a 61 5c 62 64 64 61 5f 68 56 5c 5b 57 52 51 4d 50 55 51 57 4d 52 50 4f 56 50 4e 59 54 54 5d 56 59 55 59 55 4e 53 4b 52 52 4d 49 2c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 33 33 39 35 33 31 2d 36 2f 34 32 34 39 3c 3d 37 30 35 32 2b 37 35 33 31 35 32 36 35 3a 3c 31 33 25 23 21 19 16 12 0d 18 17 26 27 34 3e 4c 53 67 97 c4 fb ff ff ff ff ff eb b7 83 4f 28 10 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 16 1f 20 30 2a 31 2f 33 36 38 3a 36 40 3c 45 47 4b 52 54 56 5f 64 54 61 5f 58 56 5f 5c 5c 54 5f 4f 53 4f 4f 56 53 49 53 49 4e 51 4c 51 51 52 4e 4d 5b 4a 55 54 57 4c 50 54 4b 41 46 28 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 31 2f 36 2c 2f 32 2d 32 2e 35 37 3b 3b 38 36 39 36 2f 2d 2e 31 3b 35 31 31 31 33 3f 33 2d 26 25 20 14 0e 05 03 06 06 0f 1b 21 2f 3a 3c 45 53 64 87 bf ec ff ff fe ed c7 9c 79 4a 25 0f 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 13 0d 14 24 2a 31 30 39 35 31 40 3d 3f 3a 3d 3f 3c 49 48 56 4f 56 5d 51 51 58 53 57 58 56 59 56 51 54 51 4f 50 4c 4f 47 4c 49 49 45 52 4f 4a 51 4b 4d 4e 4c 52 4c 4e 4b 49 49 44 46 26 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 29 2d 36 33 34 38 36 30 2e 2e 31 33 35 39 32 32 34 2e 33 2e 2f 33 30 32 2a 31 34 2b 35 2d 22 19 10 0a 00 06 05 03 00 06 05 09 16 25 2b 37 2f 41 4e 68 87 b0 c4 d4 ca bf a6 7f 5c 3d 1b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0d 0f 13 1e 2a 27 2f 2c 34 39 3e 39 35 37 3c 3b 43 3b 40 49 52 4a 4d 52 50 59 4f 53 51 4b 55 4d 51 53 4a 51 4d 47 4a 4b 4d 48 40 4c 4f 55 49 4a 47 47 4d 48 49 42 4b 44 51 46 38 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 26 26 32 3a 38 30 35 2b 2e 2d 34 36 3f 34 3a 30 2f 36 37 27 31 27 34 2e 31 31 2d 2f 2e 26 1e 13 05 03 00 06 05 03 00 06 05 05 10 15 1a 2a 2b 34 3b 4a 60 77 95 a3 9d 93 7c 5d 4c 2d 0f 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 07 0c 14 19 1f 24 2f 31 3c 35 38 32 34 3b 36 3e 41 44 43 3f 45 48 48 42 4a 48 49 4b 4c 4c 43 44 49 4a 44 46 4d 44 4a 42 49 46 45 4d 4c 4f 46 44 47 45 40 43 45 44 49 42 3d 31 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 2a 2e 36 3a 39 2f 3c 34 25 2e 3a 33 36 38 33 38 37 2e 2e 32 2f 2d 31 27 2c 35 23 21 17 11 06 05 03 00 06 05 03 00 06 05 03 02 0c 13 20 22 25 30 34 3e 4f 60 6f 6c 68 56 46 34 1a 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 15 16 22 28 2f 37 2b 33 34 2f 33 36 38 38 37 3b 41 41 3a 45 41 3b 38 44 3f 43 44 46 41 3e 3c 40 44 4e 40 3e 48 3c 3f 3c 44 45 43 44 40 3e 3b 40 3f 34 40 3a 34 35 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 2b 35 3a 39 3b 3b 39 37 2d 29 32 36 35 34 29 31 2f 2f 2a 2d 2f 30 24 21 20 27 1f 15 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0d 11 18 24 25 28 2e 36 3c 3d 41 3c 26 1c 11 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 0d 11 0f 1a 27 26 25 27 28 31 38 37 34 33 35 37 40 44 38 36 3c 3c 3c 44 40 3e 31 3d 44 44 48 4a 3d 45 3c 40 42 43 3a 38 3d 3f 42 43 3f 3d 3b 44 32 33 41 30 2d 26 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 28 33 37 45 40 40 38 3a 2f 35 34 33 30 36 2c 25 26 33 32 29 28 22 2b 23 1b 1b 1b 11 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 11 17 18 1b 1e 1e 27 21 27 1e 12 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 11 16 16 1c 23 2e 30 2f 2e 2f 39 35 3c 35 3d 3a 39 43 3b 3e 3a 3a 44 44 3e 4a 41 41 43 3d 3c 40 3d 3b 41 42 43 41 44 40 35 3e 39 3a 38 36 32 3c 3d 2a 2f 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 23 2e 34 44 46 3b 4a 3b 3b 35 2e 32 36 2f 2f 2e 2a 28 26 2d 28 1d 18 15 18 0d 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 0e 0d 12 0d 14 13 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 17 15 1d 1b 20 24 2c 2a 30 32 2c 23 39 30 38 36 33 38 3a 3d 38 40 3c 44 44 44 48 3e 3d 3e 32 39 33 33 39 3b 39 2f 31 3a 37 3f 32 35 29 34 35 24 29 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 22 42 44 35 3a 37 35 3c 3d 33 30 31 30 2d 28 2b 2c 21 1f 23 14 12 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0f 12 19 18 22 23 2c 31 34 2d 28 2a 33 35 3d 33 2d 32 30 3f 44 44 44 4a 42 40 3d 3a 2f 35 38 3d 41 35 33 37 33 32 32 30 2f 27 2e 2d 23 26 1c 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 2b 2e 2b 35 2c 2c 32 28 2b 34 28 29 2f 26 2b 2c 20 1e 10 13 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0e 1d 1d 1f 26 2a 2a 29 30 2e 31 2a 35 33 32 3b 3e 3c 3f 40 43 3e 3e 3d 36 29 35 33 3c 39 32 37 31 35 30 30 2c 2b 2e 2f 2f 23 23 1d 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 24 2e 2b 27 2b 2c 2a 2a 28 24 2e 29 2a 16 23 1a 15 13 10 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 16 1f 1f 17 22 24 2b 33 2c 29 33 30 2e 33 38 3d 40 38 37 36 35 39 34 30 2f 36 33 2d 3d 30 2c 32 2a 25 28 1e 2a 23 28 21 2b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 1d 26 28 1d 24 29 22 25 23 22 1d 21 20 1a 15 0f 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 04 09 0b 15 19 1a 17 1e 24 23 23 2a 2d 35 2a 33 2d 33 2e 27 2e 31 30 2f 32 30 2a 32 33 38 2c 36 27 25 27 26 2b 24 1d 26 1b 20 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 14 22 20 12 21 22 18 24 1d 13 12 11 10 05 06 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 07 05 05 13 1a 19 1e 21 20 1e 29 28 31 30 2c 27 27 2b 2e 2f 29 34 28 33 32 2a 30 2c 32 25 2a 23 26 28 1f 25 20 1c 1a 17 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 19 1b 1d 19 16 1d 1d 1f 0f 14 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 05 0a 0a 12 15 19 1c 15 1b 29 23 1d 25 23 2d 2b 2b 31 30 22 2e 29 2c 2d 25 25 21 2a 26 1c 23 17 1d 1b 1b 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0f 0a 05 08 06 11 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 03 07 06 0e 0f 0f 13 18 1e 23 28 22 27 1f 22 25 19 24 27 25 21 1c 1b 20 18 18 1c 17 17 12 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 11 1b 16 1d 20 17 20 1b 1d 1b 20 25 1d 18 19 14 13 15 16 15 16 14 0b 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0c 0f 10 09 0b 0e 0b 05 13 0c 0a 14 0f 0e 0b 0e 06 0b 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 04 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
