 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 01 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 06 07 03 00 06 05 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 06 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 08 03 00 06 05 0c 05 0a 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 01 07 05 06 01 06 05 05 05 06 05 08 02 06 05 04 00 06 06 06 00 06 05 03 07 06 05 03 06 06 05 03 00 06 05 04 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 00 06 05 08 04 06 07 03 00 06 09 03 09 0b 07 03 08 08 05 08 02 06 0c 07 00 06 05 03 05 07 05 03 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 08 05 05 00 06 05 03 07 0d 0f 0d 06 06 05 04 07 06 0e 07 0a 06 05 0b 05 06 05 04 0c 06 0d 0d 0d 06 0c 04 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 03 06 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 03 09 08 05 0c 04 06 05 04 0e 15 0c 16 0f 0d 16 16 0b 11 11 0d 0f 0b 0f 0c 0b 0e 0b 13 16 22 1b 1e 1f 16 19 14 0c 0b 07 05 00 06 0e 03 07 06 05 05 07 06 0b 08 0e 06 0e 04 07 06 05 0a 05 06 05 03 00 06 05 05 03 06 05 03 00 06 09 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0f 07 06 07 08 06 0c 06 08 0f 0f 17 23 21 35 2c 27 21 1f 24 1c 1f 17 13 15 17 15 20 34 3b 3a 33 3a 27 2b 24 14 14 09 11 12 11 14 0c 0d 0e 06 09 05 0b 0d 08 05 0c 08 12 13 0a 09 08 0a 0e 06 05 05 06 06 05 04 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 00 06 13 0c 01 06 05 03 00 06 05 03 00 06 05 09 0b 09 05 03 12 14 0c 1a 25 36 3b 52 67 7b 69 53 3e 39 3e 2c 29 38 27 2a 30 29 31 33 3e 42 38 2e 3c 35 39 29 1f 10 0e 12 13 19 14 10 11 0f 12 0b 11 0f 0e 08 0f 10 15 11 11 11 0c 18 13 0f 07 07 04 0d 0b 0a 06 06 0a 05 06 06 05 05 01 06 05 0b 05 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 0b 02 0f 05 07 01 07 05 07 0a 0d 0f 07 0b 06 14 0b 11 23 26 41 45 5a 5e 66 83 b7 a5 77 68 51 48 3c 3c 4c 48 4f 4f 3e 31 2d 2b 2e 26 2b 30 2e 3c 32 37 29 1f 20 1f 1b 19 17 1e 1e 17 14 1f 16 17 17 1b 14 1a 18 20 1e 20 0e 1c 1c 18 14 12 1b 15 0d 12 0a 09 0c 0b 0f 07 08 0c 06 16 21 0c 06 05 03 04 06 05 03 01 06 05 03 07 06 05 03 06 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 0a 06 04 06 05 03 0e 12 14 14 23 15 19 22 20 31 3e 4f 5e 62 6b 70 78 81 7a 70 6d 61 5d 4d 59 6a 63 62 4b 3c 2f 32 2b 2b 2b 2a 35 2c 34 3e 31 32 33 30 36 2e 2a 30 3d 35 27 20 20 2a 2a 28 20 21 31 33 39 2e 2b 29 29 2d 33 26 27 22 1d 19 21 22 19 13 16 14 14 12 0e 06 0a 13 18 10 08 0b 00 06 06 03 00 08 05 05 02 06 06 03 06 06 05 03 03 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 0a 0d 06 0c 05 0e 0d 09 10 10 17 1c 20 29 2d 28 31 3d 4a 5d 62 64 5f 61 5c 5e 5e 5d 6a 67 60 55 65 63 5f 6a 62 55 4e 4c 44 3f 3a 3d 3b 49 4a 3f 49 57 4c 50 43 41 42 36 46 45 4c 44 38 48 4a 59 42 44 3e 49 4b 56 50 3b 43 48 40 3e 46 3d 3b 3c 2a 2c 24 25 2d 28 26 22 15 14 0a 06 14 10 12 06 03 09 07 06 06 0c 0b 05 10 0f 06 06 03 02 07 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 0a 15 16 19 18 18 15 18 18 28 2d 31 33 3f 4d 43 4e 5f 73 8f 85 71 62 50 4e 5f 52 54 52 56 5c 69 6e 6e 6b 6f 6d 72 85 8a 79 75 66 5e 54 5b 59 60 66 66 69 58 43 41 42 46 42 4d 4b 48 4d 5b 67 66 6c 6b 5e 5e 67 72 83 6d 70 67 66 64 67 70 64 59 48 44 4a 49 49 45 35 34 30 28 17 21 1f 18 1e 1d 11 16 0e 0c 0a 0d 0d 0f 0b 0e 06 0a 08 06 08 06 08 0a 06 05 06 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0f 00 06 05 03 05 06 05 05 09 06 0c 0a 04 0b 14 19 17 1c 1e 24 25 17 21 2a 39 4b 56 4a 65 7d 6d 73 7c 8c 8b 78 6b 62 58 4b 5c 59 5f 64 62 71 71 7b 81 7e 82 7b 88 9b a5 a9 9e 92 7d 70 6f 73 76 72 69 68 56 44 43 48 45 49 56 5d 64 62 65 6c 65 7b 80 7b 84 81 88 87 86 7d 79 80 7c 7b 79 72 74 66 50 53 52 51 49 4b 4a 47 3a 2d 29 2b 2f 2a 25 1f 24 21 17 12 20 0f 0e 18 0b 12 0b 08 02 07 05 0c 10 07 09 0a 01 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 04 01 06 05 04 03 06 05 03 0d 08 23 31 2e 35 2f 2b 2b 22 29 29 39 52 5b 59 6c 84 8c 81 86 7c 70 6c 5a 5d 5e 64 6a 79 7c 73 76 78 76 7c 7c 8e 88 8d 8d 88 9a 98 96 91 94 84 7c 76 73 72 6f 5c 54 4d 48 4b 4e 55 5b 66 69 6b 6e 77 72 68 7a 78 83 78 8c 8b 84 83 88 85 87 80 87 87 88 7e 69 67 67 5f 51 47 55 59 63 60 57 50 50 51 45 3c 3b 35 32 20 20 26 15 1a 17 16 17 0f 0c 06 0c 05 07 06 05 03 01 06 0b 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 0b 03 04 06 05 05 00 06 05 04 11 0a 05 0b 0a 0d 12 0c 19 2a 2a 3c 3a 48 4c 4c 3f 3e 47 4c 55 5d 7c 83 87 86 88 85 79 80 77 75 7b 7a 7d 8c 80 83 81 7b 84 7e 78 78 80 83 87 8b 87 83 8c 8e 93 88 8a 83 81 81 7c 6a 5f 60 58 57 59 53 62 6a 73 82 76 78 70 78 7d 79 7d 80 89 87 8e 8e 93 95 95 96 95 8e 94 95 8c 83 7e 81 83 78 69 5d 62 67 6e 6c 6e 71 7d 83 78 77 75 6e 5a 45 31 32 30 21 1e 1f 22 20 1c 15 0f 13 13 0c 09 0b 0a 08 05 0a 07 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0a 08 05 0d 06 07 12 0e 0a 12 1c 14 0f 16 13 27 38 3f 40 40 4f 5a 5d 5f 5d 56 5e 60 67 72 87 90 88 92 84 83 84 88 87 8b 88 8b 8f 92 83 85 84 81 7c 85 82 76 7d 7d 7e 7f 7b 7d 7f 84 89 8b 8a 84 84 74 67 64 60 63 63 64 65 73 76 7c 83 93 8b 7b 85 82 8a 83 91 92 92 9a 9f 9d 9a 99 a1 9a a1 a5 9b 95 95 95 8d 91 90 88 84 73 7f 76 7c 7e 79 79 87 8d 94 9b 9e a4 92 80 71 63 5a 4d 4e 3e 41 2a 27 1e 1f 14 19 19 14 0a 07 08 13 08 05 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 0b 06 05 0c 00 08 05 08 0b 0c 0d 13 0f 12 1c 1a 1b 1d 28 2b 39 46 50 5a 69 6a 64 6a 69 68 6a 6e 67 76 7d 7d 89 8d 8b 91 8f 94 90 91 93 8d 8e 85 8a 8b 8e 8c 8b 89 75 76 7f 84 86 7b 7d 67 7a 74 75 76 7c 72 6d 6b 63 62 6d 69 73 76 81 89 82 90 90 8f 98 8a 92 8d 9b 95 9d 9d a5 a1 a6 aa a2 a4 a6 a5 aa a1 a1 92 91 94 90 9a 95 92 94 90 90 8a 85 88 84 78 7e 78 90 99 9f b3 b8 b5 b9 b6 ad 93 76 74 5d 4b 3d 3c 2c 2a 20 16 1c 13 18 0f 18 0e 0c 06 05 05 03 06 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0d 05 09 00 06 05 0f 0c 0d 05 0e 0e 14 11 16 18 10 1c 16 1d 20 28 30 30 39 40 48 52 61 60 67 65 6e 68 61 65 67 72 77 70 75 74 76 81 89 86 90 96 95 94 8e 95 91 94 92 90 9a 91 8f 89 81 79 6d 71 7c 82 87 86 7c 79 78 76 78 75 72 71 70 68 73 76 77 89 9a a8 b2 a8 a5 a5 aa 9c 9a 9b 99 9b 9e a5 ab b2 ab af b3 a9 a6 af b0 b3 af a1 a4 9f 9e a1 92 99 9b 9d a0 98 a1 98 8e 97 94 8e 93 97 a0 a0 a5 ad b0 be dd dc e6 cd b2 9c 7b 70 62 50 3c 2a 28 23 24 2e 21 1a 20 10 10 19 11 11 09 07 0e 05 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 03 0a 09 05 04 10 08 0f 09 0a 07 0c 1b 19 1c 1f 1c 21 28 2e 2f 40 3d 44 4a 44 4e 59 5c 6a 66 6a 71 6b 6d 69 6b 69 70 6c 82 88 89 84 7f 78 78 81 87 8d 99 98 9c 9e 98 94 8d 8b 8d 8c 8d 8d 87 7c 7b 79 85 8a 8a 98 8a 84 83 7e 85 81 83 85 82 87 85 8d 99 ba d6 ec de cb b6 b0 af a6 9e ad ab b7 b6 b4 b8 c1 b6 be b5 b9 b7 bf bb b9 b3 ac a6 a9 a6 9f a2 aa ac ae a5 aa 9e a4 a7 a6 a5 a4 aa a7 a5 ae ac a7 a6 a2 b1 cd e9 f1 f9 eb cd b5 9c 98 76 60 47 3e 32 2a 2d 2b 23 26 25 20 15 17 18 08 10 10 07 07 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 04 07 05 03 09 06 0b 0c 05 15 0d 0c 12 19 15 1b 20 2a 35 3c 3b 57 59 6e 6d 5c 44 4f 50 56 54 5d 70 64 72 6a 6f 74 76 6c 72 70 7e 85 7e 83 7f 7f 86 86 7c 76 7e 8d 85 92 94 90 8d 7f 7f 8e 81 8b 86 82 84 83 89 89 88 8e 9a 91 93 8a 90 8b 94 8a 86 92 9d 9e ba cd f7 ff ff f8 dc c0 ba b7 b5 b5 b8 b6 c6 cb c6 bb c8 c1 be c1 c3 c1 c6 bf bb b6 b3 af ae b3 a9 aa b3 b8 b2 b2 b2 ad b2 b5 b7 b2 b0 bc b5 aa af b3 b2 b1 b0 a8 b6 ba c4 dc f7 fd f1 ec d1 bf b2 91 79 5c 51 42 47 40 3d 37 31 22 21 26 1d 20 16 10 08 0e 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0c 05 03 07 06 0c 0e 0d 0c 10 1c 1f 1c 2e 34 49 56 58 66 71 84 99 95 8d 80 5c 51 4f 51 5b 61 5b 5d 5e 70 68 6a 82 84 7c 85 88 80 6e 75 77 74 87 86 84 83 87 82 79 7a 84 85 8b 87 89 85 86 8e 8f 8c 97 94 93 8b 95 9b 9e 9d 99 98 9b 9b 94 9f a4 a9 be d8 f7 ff ff ff ff ff e5 ca c2 c2 c4 c0 cc d3 d8 d1 d3 d4 d1 d1 cc c8 c4 c7 c4 c3 c9 cb be ba c3 bc bd c2 c1 bc b9 be bd bf ba bb c1 c8 bf c2 c2 ba b3 b5 b6 b8 af ad b4 b9 b1 b8 c5 d4 d9 e9 e4 e3 d7 c8 b4 a0 91 87 7b 69 5e 55 45 35 30 2d 2c 23 1e 16 0e 0e 08 06 12 0a 0b 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 07 06 05 08 06 06 05 0d 09 09 0d 06 0e 0c 0c 18 16 23 30 32 3a 51 61 70 7c 8f 86 87 87 99 a5 ab 9e 96 7f 63 5b 5e 5e 5b 5e 5b 61 61 5f 63 75 7a 7d 86 8a 86 7a 7b 79 7a 7b 83 83 83 8e 98 99 8c 87 87 86 91 8c 8e 8e 98 98 97 98 90 9a 9b 97 a3 a5 a9 ab 9b a7 a3 b1 c0 d0 ed ff ff ff ff ff ff ff ff e4 ce c4 c9 ce d5 db e7 e4 df e0 e3 d8 d8 d8 d3 d3 d8 d9 d1 d5 cd cb cf d4 d8 d0 ce cc c5 c8 c8 ce cf d0 c9 c5 d2 ca c6 c6 c8 c4 c3 b4 b9 b3 b6 b5 b7 b8 b5 b5 ad b1 b8 b6 b9 be c3 bc b4 ac ae a6 9d 89 78 61 4c 4d 3b 3b 30 27 25 1e 12 1c 0f 17 0a 0f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 07 01 06 09 07 02 0d 0f 10 17 17 1b 22 3d 4b 66 6e 78 87 8e 93 9c 9c 94 9d 96 96 97 a6 a6 b0 a7 89 6c 65 60 5e 60 59 63 61 5f 65 77 69 78 7b 7c 87 7d 80 84 7d 85 83 81 7e 81 90 95 9c 9b 9c 9e 97 96 93 9a 95 a1 a6 a6 a4 a0 a4 a4 a5 a8 ae ad a7 b0 bf dc ed ff ff ff ff ff ff ff ff ff ef e0 d9 df da e0 e5 e6 e7 f3 f3 e9 e1 e6 db d9 e1 d5 d8 e0 e2 e2 de df df e2 e1 db d7 d4 d1 d1 d6 d4 d4 d4 ce d3 ca d0 d1 cf cd c7 c2 be bb b7 ba b5 b4 b3 b3 b7 ab af ab a6 a9 9f a3 9f a5 9a a2 af bf b5 a6 88 73 6d 5f 4e 44 38 32 2b 19 26 1e 24 16 12 10 0f 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 0c 10 06 09 06 0e 14 25 32 36 4a 57 65 80 86 93 97 9e a2 a2 a1 a4 9c a3 9e a4 a4 a8 b8 c0 c1 b3 9b 7e 72 65 6b 63 61 66 69 66 68 64 63 7e 7d 7c 87 84 84 8d 8c 8a 81 8e 8e 91 9d 9f ab ab a7 9e a5 a5 9f a9 a1 b6 b3 a9 a1 a8 a0 ad b4 b4 b9 c6 cd d6 e4 e6 fd ff ff ff ff ff ff ff f4 e6 de e0 e1 e3 eb ee f3 fe fd fb f5 f0 eb e5 e0 e6 e0 ea e6 db e2 dc e9 e6 e3 eb e9 e3 e2 e3 df d8 dc d8 d9 dc d0 d5 cc d0 cc cd c9 be c4 b6 b8 b4 ba c0 ab b1 b3 a7 af b3 aa a5 a2 9e a1 9c 9a 93 9f a1 b3 c9 be 9f 92 70 6b 62 55 4e 3e 38 32 2a 24 25 1f 0b 0e 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 03 00 06 05 03 00 06 0d 08 0e 0e 0c 14 24 2c 3c 4e 66 6d 7a 89 94 93 a4 a1 a3 ab aa ae af ab aa a5 ab aa b1 a8 a7 ba c8 d9 cd c9 b9 9e 90 88 7e 77 7a 77 80 7e 82 83 90 92 91 91 9c 8c 94 98 a1 95 98 9b a9 a7 b1 b5 ab bb af b1 b4 ad b4 c1 bc bb b8 b4 b4 ba c0 bc c8 df cf d7 d6 de ea fb ff ff ff ff ff f3 e9 de e8 ea f4 f1 f5 fd f9 ff ff ff ff fc f1 f4 f3 ee f0 e8 ee e4 ec e9 f1 f2 eb f5 f0 e5 ee eb ee e8 e5 de dd dd d4 d7 de d0 c9 cf c7 c3 c6 c0 b6 b6 b6 b0 b7 b0 a9 b1 b6 b0 a1 a4 a1 a6 9d 92 95 92 9e 8d 90 a4 c1 c6 b9 a5 90 84 76 66 5d 51 4f 47 37 30 26 16 10 06 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 06 05 06 00 06 0b 03 02 06 05
 12 10 12 10 26 31 49 68 80 8a 90 97 9f a1 a6 ad af ae bc c4 b1 ba b6 b2 b7 b2 b0 b6 b4 b5 ba bd d1 dd e6 e3 d7 d2 c5 b5 a9 98 99 9f 9b a1 a7 9c ab a2 9f a3 af b3 b5 b2 b3 bb bb c5 cd da d2 db c9 c7 cb bd c2 c0 cc d6 d1 cd d3 c6 c9 c7 cd dc ef ef e6 dd d7 de f2 f6 ff fe f4 f5 eb ea f0 f0 f4 fa f8 ff ff ff ff ff ff ff fe fb f3 f6 f1 fb f8 f3 f8 fb f5 f2 f9 f5 f7 f6 ee ee ee ea e6 e7 e0 e1 df e0 d9 d4 d9 d4 cb cb c3 c1 b6 b9 b8 bb bc ad b9 b4 b3 b2 b2 aa a3 9d 96 9e 9c 99 91 9b 94 91 94 a0 ad be c2 b2 a3 99 8d 81 7b 62 53 45 33 22 13 15 0d 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 1e 0e 03 09 06 05 03 0d 07 09 0f 1d 20 2d 45 4f 70 85 90 96 a3 a2 ac ae a9 b4 be bb b9 c7 c9 bc c4 c4 bf be bd b9 c0 c4 be c2 cc d2 d4 e7 e8 ec e4 d6 db c6 cd cb d6 da dd e4 d2 d0 cb c4 c6 cf da e0 d7 de d1 d2 dc ed f3 ed dc cc d5 d2 d4 d4 df e3 cc d9 d2 d4 dd df ef fb ff ff fb ec dd df e8 f3 f0 f2 ee ec ef f3 f1 f6 f7 f7 f8 ff ff ff ff ff ff ff ff ff f8 f9 fb f7 fb f8 fd fe f8 fd fd f6 f3 f7 f7 eb f0 e6 e8 e1 ee e4 e4 da db dd d0 cf cc c8 c0 c2 c1 be b4 bb b4 b2 b5 b2 aa ad a7 9f a1 99 99 9b 9a 98 95 8a 92 8f 8a 8e 90 98 a1 ad b7 b9 ab 99 8c 7c 68 4d 38 2b 1c 0f 12 1b 07 09 09 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 1e 30 2b 28 12 07 14 09 0b 0f 07 1e 33 3f 52 73 8d 8d 9a ab a0 ac b0 b8 bd bd b9 c0 c5 cd c8 ce d2 d1 cd ca c4 c5 cc c1 c7 ce d1 d4 dc d8 da de e4 e7 e4 e4 e1 e1 e3 e3 f4 fe fd fe f1 e5 e4 e3 ec e9 ed f5 f0 ed e2 dd e5 ed eb f0 e9 e2 e4 e6 e2 e6 ec e1 e0 de d9 eb fd fe ff ff ff ff ff ef e6 e9 f4 f3 ea ed fb f5 f9 fb f1 fc fb ff ff ff ff ff ff ff ee ff ff ff ff ff fc ff fe fb f7 fc fb fc f6 fa ff f5 f8 ef f2 e9 e7 e2 e6 e6 de de d8 d8 d5 cc c7 c0 c2 bb bb b7 b5 be b9 b5 ae a8 a6 a9 a8 a2 95 95 93 9a 93 95 95 8d 8d 92 94 94 98 98 9d a1 b0 b6 b2 9a 89 6b 65 4f 41 25 29 16 19 15 15 14 10 0f 0f 08 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 2a 39 31 34 22 0f 17 10 0b 1c 29
 33 44 5f 7d 92 95 9a 9c ac b6 b6 bf c1 d0 bd ca d5 d6 de dd df e1 db e0 e4 d6 d5 dc da dd d7 e8 ea e4 e7 e5 e8 ef f5 eb f8 f0 f5 f9 fb ff ff fd ff f6 fb f0 ff f8 fe fc fe fc fe fa f2 f7 fb f5 fc f2 f9 f3 f9 f0 f1 ec ed f1 f2 f0 f7 ff ff ff ff ff ff ff ff fb fa fd fc f4 f6 f6 fb ff fb ff ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fe ff ff fa f9 f6 ee ea f3 f1 e1 e2 d9 de db d8 d1 d0 c8 ca c0 c1 c6 ba be ba b3 ae a7 ab a4 9f a6 9e 97 9b 9c 9c 99 95 93 91 93 8d 90 91 90 91 92 8f 90 9e a5 a5 93 85 74 66 4d 3c 29 2b 1f 24 13 1c 12 16 10 0c 08 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 10 20 26 23 20 0e 0c 17 10 1a 24 31 43 5e 80 9c 9d 8f 9f 9e ac b8 c2 bd ce d4 dc d9 e7 e8 e2 e6 eb f2 f2 ee e9 ea ea e5 e3 e4 e8 fa fc f1 f5 ee fb f7 f9 ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff fc ff ff ff ff fd fa fa fb f8 ff ff ff ff fe f8 fe ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f9 ff fe fb fa f4 f4 ee e8 e7 e4 e6 db d9 d4 d3 ce cc be bc b6 be be be ac b3 a4 a1 96 a5 97 9d 98 93 98 8e 8a 8d 90 8f 8b 95 87 89 85 83 87 85 81 83 84 8c 8b 8b 7b 76 65 55 46 31 26 1e 23 1c 0f 0f 16 10 04 09 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 1c 17 16 13 0b 0a 1d 1f 20 37 38 58 78 90 a5 92 93 99 a2 a7 bd ba c2 cc d3 e1 e9 f1 f2 fc fb fd fe ff fc fe f7 f4 ef f9 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff ff ff ff ff ff ff ff ff f6 f0 f9 f2 ec e3 e5 dc da d4 da d1 c4 d2 c6 bc c2 bd b9 a7 ab 9e 9a 96 9a 92 93 92 95 96 92 8d 89 8f 86 84 83 85 81 85 7f 77 7a 75 70 7a 74 7d 7c 80 7e 76 73 68 46 34 28 22 1b 1b 0f 23 20 16 0d 0a 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0c 06 0d 13 0e 11 15 16 24 2b 34 3d 4e
 6a 80 98 aa 9f 9b a1 a2 a4 ab a8 be c3 c7 dd dd ec f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 ff f4 ef f1 e9 ee eb e5 da d5 d6 d4 cb cb c4 c0 bc bf ab a5 a9 9e 9f a0 9c 9b 87 8d 94 8c 8f 90 87 8a 88 82 83 86 80 7b 81 74 76 6d 64 68 75 6b 72 7a 7f 7e 77 58 58 3c 2f 28 1d 1c 15 1e 1f 1e 1b 11 09 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 07 05 08 15 0d 12 1c 24 2e 30 42 43 53 7a 92 a4 af 9c 9a 9e a1 a1 aa a9 b0 b0 b7 be cf e4 e5 f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb f4 f6 f9 f2 f3 ec ea e5 da de d1 c8 c6 c3 b7 af b0 a9 a9 a9 a1 9f 9d 98 99 86 89 82 84 8d 8c 8c 89 82 86 7b 73 7d 76 77 6c 6d 6e 6f 62 62 6e 67 66 74 6f 70 6e 60 51 3f 30 24 27 1c 1e 2b 31 22 18 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0d 06 10 17 18 1a 0f 28 2f 3c 45 52 69 81 93 98 a6 a8 9c 90 9e 9d a0 a9 ab a6 b1 b4 ba c6 d2 d8 ea f0 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 f3 f5 f0 f1 ef eb e5 db d6 d2 cf c4 bc b6 b5 b4 ad a8 ad 94 9e 97 95 95 92 87 8a 8f 94 8b 90 8a 7d 81 7d 71 77 79 74 6b 6a 6b 6c 61 62 5d 5a 65 64 73 6b 72 70 65 56 3a 32 2d 2a 2e 3a 31 34 2a 1e 0f 0d 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0c 05 08 0c 0a 12 1c 1b 24 22 31 2f 53 6f 7c 97 a7
 9a 9f aa 9d 98 92 99 8f a1 b1 ae ab b6 b0 b8 bf ce dc dd ec ed f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff f7 fb f5 ef e8 e3 d2 ca c4 c5 be b4 b2 b3 ad a2 a5 a4 9f 98 98 94 95 93 90 97 95 94 92 81 81 85 7b 75 76 77 6b 73 6a 69 62 60 60 5f 5e 5b 61 64 6c 6c 6e 71 65 45 3e 38 40 44 43 3a 36 2d 24 12 0f 12 09 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 05 0e 0d 0e 1a 13 1c 17 25 28 37 3c 5c 7c 9a b2 ae a7 a1 9e 92 90 94 95 99 a5 a2 a5 b2 b4 b7 be c0 c7 ce de df ea fa f6 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe f4 ec e4 e0 d2 cb c8 c7 ba b7 ac bc ae a7 a7 a0 a1 a5 9c 9e 96 9b 95 93 95 97 8f 8a 82 81 7e 72 6f 71 74 6d 68 6d 63 5b 58 5a 5e 5b 5a 61 5d 6b 6b 77 6f 64 55 52 4d 58 52 41 3a 33 26 1e 17 13 06 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 08 0b 0f 12 12 19 15 26 35 40 47 53 86 9e b3 c6 af a6 9a 9c 8c 91 9d 9a 9b 9e b9 ae b4 ba b5 b8 c9 ce cf dd df e7 ef f9 f2 f6 f4 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f5 f8 eb e0 d2 cd c7 bb bc c1 b8 be bd b4 b1 ae a9 ad af a5 a1 a2 9a a5 95 92 94 90 8e 81 87 81 6c 73 6d 78 71 62 65 65 5c 59 5c 59 5a 5a 56 59 60 5f 5e 70 73 77 7a 73 68 60 52 41 41 29 21 1c 11 15 10 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0f 11 14 0f 1b 1b 1b 1f 21 31 3c 47 62 87 a4 b2 b6 a5 9b
 9f 90 93 9a 97 a0 a1 a1 b1 b0 ba bf bf ce cd cd da d1 d4 e5 eb ed f5 f7 ef f4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f0 e1 dd d0 d0 c6 c2 bf c0 c4 bb bd be b7 b6 bc b3 b2 b1 b8 b1 a5 aa 9e a0 9d 9e 91 86 7e 7f 79 7a 79 6f 6e 67 6f 6d 69 71 5a 5f 5a 5f 56 60 5e 58 63 6f 82 82 87 77 74 6f 5a 50 45 3c 28 22 21 14 0e 0e 0e 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 03 06 08 0d 16 1a 18 21 1e 1e 19 24 2c 34 4c 65 81 9e b2 b0 a3 97 95 96 93 93 9b a7 a2 a7 b4 be c6 c2 c6 c7 cd cd d7 dd da df ea ea f6 ee eb ef ed f5 f3 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f0 e6 e0 db d2 ce ca cb c0 c7 c7 c4 ca c6 c3 c0 c4 bb bf bb ba b7 b5 a5 a9 a2 9b 94 89 86 85 7c 78 73 74 71 71 6e 6f 6c 64 65 57 67 5a 60 5d 66 62 5b 59 63 69 70 7d 74 6c 60 67 64 52 49 33 2d 21 1b 15 18 14 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 05 03 10 11 0b 0e 1b 16 1d 24 23 29 27 2f 3c 51 63 83 9b a7 a3 91 93 90 8e 97 92 95 9d a4 a7 b4 b9 be c1 bf cc ce d4 d6 db de e2 e6 e6 e8 ef f0 ee ef ee f1 eb f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f4 eb ec df d7 cc cf c6 cd d8 c9 d3 d2 cf cc d1 cb c8 c5 c4 c4 b5 bb b8 ab a5 a4 9d 99 93 85 83 7e 7e 7a 79 77 6e 7b 74 6a 66 65 68 6d 67 6e 63 5d 6b 5f 66 60 67 5f 5f 5c 5b 5f 71 6c 61 4b 3b 35 20 1b 21 18 1a 10 10 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 03 0c 0a 13 14 13 0d 1a 16 1f 20 2d 36 3c 3d 53 61 76 83 8c 9c 9b 8c 8c 8c 94 8c
 94 9c 9f a2 ad b4 b5 bf c3 cb c8 d0 d5 db dc da dd d9 e2 e7 e3 e4 e3 e8 e7 e9 ed f5 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ef e7 e4 d9 d6 d8 d4 d1 de df e1 de df da d9 d4 d1 cf c9 c7 c5 bc b9 b2 a6 a1 9b 95 91 85 86 89 7b 7e 7c 7f 71 78 7b 70 70 70 75 70 69 6f 61 69 69 67 63 67 60 58 61 5b 5e 5c 71 79 75 64 5d 49 3f 33 27 24 1e 17 07 07 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0e 08 0b 13 15 10 11 15 1b 1f 29 26 38 4d 6b 72 81 88 94 93 8f 8b 89 90 92 95 98 9a a4 a1 a6 b0 b0 b6 ba be ca c6 c5 d4 d6 da d7 d4 df e5 e6 ec e9 ea eb f8 ef f7 fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 f1 e0 dd dd e1 de e7 e1 e3 df e6 ea e7 e0 d7 dc dc d1 d1 ca cc c7 ba b8 ae a2 9f 9b 94 91 8d 83 7d 82 7d 81 82 7d 7e 75 74 7b 82 7f 78 73 70 7e 72 6b 6d 66 66 62 65 5d 61 5e 71 87 87 79 65 52 47 3b 31 36 30 27 1c 0e 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 08 07 11 0c 13 1a 15 1c 24 29 33 56 6b 70 89 89 86 89 80 8b 88 8f 95 8c 98 95 a2 9a a7 a8 af ad b1 b1 c1 c3 c6 cd cf d6 dc e2 e0 e2 ed ea ef f2 f4 f1 f2 f5 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f3 ef ef e8 eb e7 ed ed ee ea ea ec e9 e9 e3 dd da cf d7 ce c7 c4 bc b8 b0 a6 a5 97 9c 94 8f 8d 8d 88 82 89 8d 82 89 85 7c 79 7b 85 7b 72 7c 79 77 6f 6f 6a 6b 6b 6b 65 62 55 5a 6b 84 8f 86 6e 6b 50 52 48 41 3a 2f 27 15 0e 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 12 1a 19 1a 23 20 28 30 48 5d 7a 74 77 7e 84 86 86 8b 86 8b 87 8e 8f 8f
 9e a1 9a a6 ae b0 ae b6 bc c9 ca cc da d7 e5 e2 e9 e3 f4 f9 fa f9 ff ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fb f7 f0 f3 f0 f9 f5 f5 f4 f0 ee f3 f3 e4 e2 db d2 d4 d6 ca c7 b6 b9 ab ac a3 a2 a5 a1 96 91 94 86 83 8d 90 92 95 89 80 7d 86 84 7a 84 80 81 81 78 75 72 69 70 71 61 60 62 54 5e 77 8d 8d 89 7b 72 66 5b 4c 44 38 35 2f 10 0a 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 01 06 13 17 1f 17 1c 1f 27 32 3d 4e 62 6b 73 74 78 85 85 8a 87 88 86 8b 90 8d 94 95 9f 99 9c a4 af b2 b5 bb c6 cf d2 d7 e4 dc f0 ef ee fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fb ff ff ff f6 f6 f3 fa ec ed dc dc dc d6 d0 c7 c5 c0 b9 ad af b3 a5 aa a5 9c 9e 92 95 8e 97 92 8c 92 8e 91 94 88 89 8e 80 82 8a 7d 84 77 78 80 74 74 67 68 6a 5d 61 5e 64 7a 83 8b 8f 84 7c 64 5e 53 41 3b 34 2c 1d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 15 18 19 15 1b 23 2e 39 44 53 5f 64 73 79 82 81 83 84 82 82 8b 91 89 82 92 97 99 9a 9b a0 ab a8 b9 bc ba ca cb d1 dd e1 e8 f5 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fe fd f1 f2 eb e9 ef dd de d4 d1 ce c4 c5 b8 b6 b0 af a9 ab 9c a6 99 9f 93 8f 93 94 95 90 92 97 93 91 8e 8a 85 87 85 8c 80 83 7a 7c 70 79 6f 72 66 6a 64 5e 59 5d 69 6d 7b 91 8c 7e 76 6d 5a 53 45 37 30 28 1a 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0a 1a 2a 1e 26 2d 26 32 32 52 62 5d 75 70 69 79 7f 81 82 82 86 87 8a 8e 8c 92
 96 97 9a 98 ae a5 ad b7 b5 c5 c9 cb db e3 e8 f7 f6 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff f5 f5 f2 ee f0 ef d9 de d3 c7 c5 cb c5 ba b9 b7 b4 ab a7 aa ad 9b a0 9f 9e 97 9b 9b 8f 94 96 95 93 91 95 88 8e 81 84 76 7e 7b 74 73 6c 6b 69 6b 6d 60 5d 6a 5d 67 65 73 8a 91 99 8b 76 6b 58 4d 39 34 2e 1a 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 06 09 0e 19 21 24 25 25 36 36 46 49 65 61 6a 74 6b 71 75 7d 78 7a 7f 82 87 88 8f 85 9c 9b 9b 9a 9d a8 a4 b0 ac bd c2 ce ca df e4 eb f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe fb f8 f7 f5 e9 e3 ea d6 d6 d4 c6 c2 c4 be bf bd a9 ab ad a5 a8 a2 ab a0 9c 9e 9e 96 97 a2 98 8d 97 94 91 92 8b 82 85 87 85 84 78 7c 73 6f 6e 6f 67 69 66 63 5f 65 66 71 6c 83 96 8d 8d 84 6d 61 58 45 3d 2e 20 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 0c 18 1c 1e 27 33 38 45 42 4f 58 5d 66 60 6a 69 70 7c 71 7b 79 7a 81 80 92 8e 91 9a 9c 9b a6 ae b1 ad b6 bc bf bd cd d6 db e3 e7 f9 f8 f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f8 f1 e4 ec e5 d8 d4 ce d2 bb c7 bd b6 b3 b4 b4 b1 ad ae a9 a8 a6 a0 a7 a1 97 94 99 97 a2 94 92 94 8a 90 8c 8b 87 87 81 79 7d 7c 7a 73 77 69 69 6d 6a 6a 65 73 70 6f 6b 7b 8a 98 93 83 76 69 59 52 45 3c 1b 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 07 08 06 1c 25 23 34 33 49 44 44 5a 69 61 63 68 73 74 6f 71 6a 79 79 7a 79 78 90 8f 9c a5
 ad ad ad b3 bb bb c2 bf c8 ce cd e3 e0 de ec f1 f3 f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 ec f1 df e8 d8 d9 cc cd c9 be c1 bb b2 aa af a7 b2 aa a8 a6 ab ae a9 a4 a6 a0 9d 95 93 9a 8c 95 85 83 8e 8c 8c 80 8b 81 87 81 7c 79 80 73 6d 75 6e 65 69 73 6e 75 66 6f 69 87 9e 99 9b 81 6c 62 58 49 3a 1f 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 02 08 11 11 27 2d 26 38 3e 40 49 48 5f 70 6b 69 6f 6f 71 75 74 71 7b 7b 7a 88 91 96 99 a7 9e ab b5 af b1 c3 c0 c4 cf d5 c6 da db dd dd e3 e2 e4 ef ed fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fb f4 ea e2 df da d3 cf c2 c9 c0 b7 c1 b4 b7 b6 a9 b0 a5 a9 a5 ab af 9f a8 a0 a0 9c 92 9a 9e 99 97 8f 92 83 8e 85 8d 92 7e 85 88 7f 80 7d 7e 7c 7d 7c 84 6f 74 79 73 6e 76 68 6f 6f 8d a4 98 8b 7f 6a 60 51 44 30 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 07 04 0a 07 19 24 30 2f 46 46 41 46 59 61 72 69 6f 72 6b 64 6e 78 76 7b 7e 84 89 98 99 a9 ac ad b7 b2 b9 b8 c6 c7 c7 d0 cf cb ce d3 d7 dd d8 dd d8 e8 e6 ef f8 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f6 f6 e8 e2 d9 dc cc d5 d2 c5 cb c0 b4 bb b3 b6 af ac ab a6 aa aa a9 a2 a5 a9 a3 9a 95 93 94 8f 92 92 8c 93 8b 8b 87 8b 86 8e 8d 87 82 7f 7d 84 7f 85 7a 79 74 74 7b 7a 70 69 68 69 64 82 a6 94 93 7d 74 5e 43 3e 29 15 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 15 13 22 34 39 3e 3f 4f 50 4f 61 7c 7b 74 70 6b 6b 69 66 72 78 87 8c 97 99 a3 a8 ab b6 b1
 ba b5 bc c3 be bf bf c5 bd c7 ca cd d2 d2 d9 d3 e1 df da ef ed f0 fc f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e9 e9 e4 e2 e0 de d0 d4 c5 c4 c4 be b8 b6 b9 b5 ad aa af ab a6 a8 a5 9e a2 a5 99 9f 9a 95 92 98 94 90 90 8d 83 8c 8c 8b 92 8f 86 8f 8b 84 85 8a 80 84 7f 7f 79 75 71 6f 6a 5f 62 65 6b 7b 98 a5 95 8e 72 64 55 40 2f 1f 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 06 0a 12 1e 27 30 32 42 52 54 5c 64 68 7d 88 86 70 71 6d 66 6a 7f 85 8d 92 9d 9e a3 a9 b2 ba ba b6 b2 b2 bc be b6 b8 be c2 c0 ba c2 c6 ce d6 cd d8 db e2 e4 e3 e6 f1 ef f7 ff f8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f8 ed e9 e5 e1 e1 d9 cd d6 cb cd c5 b8 bb b6 b6 b2 ba a8 b0 b0 a7 a0 a4 9e a5 9c 96 93 93 9c 92 97 8f 8d 8e 8f 8b 90 91 8e 92 91 90 84 8a 85 89 83 86 7e 7e 7e 74 6c 73 73 6e 66 69 63 6d 69 7a 8c a6 a6 87 7f 63 59 50 37 28 15 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 06 05 10 0e 15 26 2e 37 37 46 50 5e 63 60 69 7a 87 86 77 70 6e 75 7b 7b 85 97 97 a3 ad b2 b0 aa a6 a5 b4 a6 ae ad b7 a9 b6 b6 b9 c4 c7 c4 c6 c5 c9 d5 d5 d8 dd da e3 e1 ea ed f7 f6 f2 fc f8 f8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f8 f1 ec e2 dd d8 d3 d1 d3 cc c5 c8 c0 bb ba ae b4 ae ae a9 a6 a7 a9 a3 a6 99 a5 9b 97 9f 9c 93 92 93 92 8c 93 94 9a 99 96 92 8b 89 8a 87 84 83 86 7f 7e 7d 74 75 72 6d 6b 5e 64 6a 69 67 6c 63 6f 7d a6 9d 92 85 73 65 55 37 28 15 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 0a 14 21 2f 3d 44 4a 55 59 65 72 71 75 7c 85 80 6f 6a 6c 74 86 8c 9b a0 a8 a7 b4 ab a3 a8 a4 9b
 9e a1 a6 a7 a4 b4 a9 b3 b6 ba b8 c0 bd c6 ca cc cb ce d5 db e3 e0 e0 e5 ea ee e8 f0 f0 eb f0 fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f8 f2 ed ea eb e1 de d2 d0 d3 ca c7 bf c4 c1 b6 b7 b3 ab a9 a8 aa a5 a5 a2 a0 9c a0 9c 9a 9d a1 9d 94 91 9b 90 98 91 90 95 8d 94 89 88 85 8b 88 84 78 7a 79 7a 7a 74 77 70 6c 6d 6f 68 6e 6a 6b 65 6f 6f 7e 9c a1 90 8c 72 63 50 3f 30 18 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 0f 12 1d 2a 31 39 43 54 60 69 6f 73 71 7b 7d 77 6e 6c 71 77 81 81 90 96 a5 a7 a4 a5 9f 9d 9e 9f 98 99 9a a5 9c ad a3 a9 b0 b7 b3 b9 b9 c1 be be cc cc d2 d0 d7 d3 dd df e6 df e2 e6 ed f0 f0 ee f5 f7 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f6 f2 f1 e9 e5 e3 d8 cc d2 c3 c7 c7 b8 c4 b6 ae b5 af ab a7 aa a5 a6 a6 9b a4 9a 99 9d 9f 9a 9f 93 9b 9a a1 97 a0 9b 9e 98 94 90 8e 81 81 86 7c 86 7e 81 77 67 76 73 77 71 6d 6e 6b 6a 73 67 67 72 6f 6b 80 97 a4 9c 8b 7a 62 5c 41 2d 1a 09 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 14 2d 3e 45 4c 4c 5b 64 73 80 75 6d 6e 71 6c 65 67 68 72 83 87 8f 9d 9b 9d 93 96 94 8c 8e 98 97 98 93 9d a4 a8 a1 ae ab b0 b9 ae b6 bd c1 c5 c7 cf d5 d3 d5 d1 d8 d6 df e2 e2 e3 ea ee ea ee f3 fb f4 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe ee ed e8 e7 dd dc d3 d7 d5 cb c7 bc b6 ba c0 aa b2 b0 a7 aa aa a5 a2 a7 9d a2 9f 9f 9e 9e a6 9c a6 a0 99 9b 97 97 9e 93 91 8f 85 8d 81 81 85 86 84 84 73 7f 7f 74 73 6d 6e 6d 6e 72 6d 72 66 77 72 71 74 76 76 85 a5 a1 98 7c 6d 5e 4c 3c 13 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0a 13 28 30 46 47 4d 5d 67 74 7d 81 7d 6d 60 59 64 6a 64 70 78 76 87 82 95 91 8e 8e 86 8f 90 8b 86 8f
 8d 8e 95 96 9e a3 a2 ab ae a9 b2 b7 bc c3 c2 c4 c9 c7 d4 d0 d1 d6 d7 d9 dc e3 db d7 e1 e2 de e4 eb e5 f6 f4 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f5 f5 ed e4 e0 e3 d3 d7 cf cf c9 c8 c6 c1 be ae ba ac ab af a1 aa a5 a0 a4 a0 9a a1 9e a1 9f 9e a6 99 9c a3 a1 9c 9c 9c 99 8f 89 86 84 85 8b 80 87 85 7d 77 7d 74 71 6a 6f 69 68 6d 6e 65 6d 73 6f 6f 71 73 77 72 72 7d 96 a8 98 82 6e 66 43 34 1f 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0e 21 35 41 4e 54 4f 5e 6f 7d 82 8f 7c 61 62 5f 5e 65 6e 72 78 82 85 89 90 83 89 8a 8d 89 86 7f 85 84 8a 90 8a 95 9d 9a a4 a8 a9 ad b4 b6 bd bb bd c9 ca cb d2 d2 cf d8 d8 d2 db cd d9 d0 d9 db db df e8 e4 ec f2 ed f9 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 ec f6 eb e6 e1 e0 e1 d7 cc cc cb c5 bc ba b8 b2 ae b4 af ae a7 a7 9e a0 aa a5 9e a7 a0 9f 9c 9d a5 9e a2 a1 a2 99 9f 91 96 90 8e 8e 85 89 7d 7c 76 7e 7a 7a 79 77 72 72 6d 6f 6b 71 6f 6a 6d 74 74 73 72 76 75 73 78 84 90 ac a5 90 78 69 50 35 15 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0f 35 3a 42 59 55 5a 6d 79 7d 92 91 7b 65 59 5e 5b 64 6a 6e 7b 78 7f 85 7f 82 87 85 80 84 78 78 7b 7c 89 8a 8b 91 95 9d 9f 9c a4 ae ac b5 b8 c1 be c9 c2 bb cd cd c6 c9 cb cb d2 d1 cb d1 d3 d2 da d9 dc e6 e4 ea df ec f6 f1 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f6 f0 f4 e8 eb e5 db de d6 da d6 d0 cd c8 c5 c0 bb b3 b5 b9 af ad ae a9 aa ac a0 a7 a0 9f a3 9f 9d a3 a4 a6 9f a4 ab 9a 96 97 98 95 8a 86 88 83 82 82 7f 7a 75 74 73 73 72 77 79 6a 73 76 75 76 78 6b 74 79 78 74 7a 78 78 75 74 8d a5 a5 8e 83 63 47 31 11 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0b 1d 2b 46 4d 4c 53 64 78 77 84 8e 8f 7e 5e 61 5f 67 66 66 71 7a 77 84 7f 7d 83 80 74 75 76 76 79 7b 7d
 8a 84 8e 8b 8d 9b 9b a6 ac ae b3 b7 bf b6 bd c3 bf c0 c6 c4 c1 c7 c4 c8 c5 c7 ce cc ca d6 d5 d6 d6 df e2 e1 e2 e4 ed eb f5 ec f1 f9 f8 fc f8 ff f8 ff ff ff ff ff ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f8 f0 ed ed ee e6 e5 dd db da d5 cc ca c4 c4 c3 bb b5 be b9 b2 ae ac a9 a0 a7 a5 9f ad a6 9b a3 a2 a3 a0 a5 ab a2 a3 a0 99 9b 91 92 97 90 87 83 74 79 7e 73 78 70 74 7a 6e 78 6c 74 77 78 75 6a 77 78 76 6f 7b 78 75 74 73 75 7a 80 91 a3 ac 99 74 5e 47 2a 15 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 21 34 4c 54 56 66 73 7c 80 87 93 92 85 65 62 64 5f 68 69 6d 73 71 7a 7b 75 73 78 6f 74 7d 72 7f 86 81 86 87 8f 93 95 9b a2 a6 aa a6 b1 b6 b1 b5 b2 bb c5 b7 c0 bb ba c0 c7 c4 c4 c2 c4 cc d4 d1 d1 d1 db e0 db e2 dd df e3 de e6 e5 e5 f3 ef f6 f4 f2 f8 ff fe ff f7 fb fc ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 ee f6 e9 e9 e3 e3 d9 e4 e3 d9 d4 d0 c4 c4 c6 bd c1 b4 ab ba b9 ae b8 a9 ab a4 ac b1 a6 ac a6 a2 a9 a9 a9 aa ab 9d a0 a5 98 9b 96 8a 8e 82 85 80 78 79 75 73 74 73 71 77 74 71 7a 74 7b 74 72 81 75 77 76 7d 81 76 7e 79 7b 7e 80 7f 92 a1 a9 95 76 60 45 28 15 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0f 1e 3d 49 56 62 65 75 7d 84 8a 96 9b 8a 69 66 66 66 67 6d 71 74 7a 78 7a 6a 6a 67 6a 71 76 7b 7a 7d 81 8e 8a 90 91 99 97 9e a5 a8 ab a9 af ad b7 b2 ae b3 ad b5 b5 b3 b5 ba bc b6 bd c6 b9 c3 cd c4 d9 d9 d8 d8 e4 dd df e0 dd e6 e1 e8 e5 e0 e5 e6 f3 ed e6 f1 ee f9 fb f9 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa fa f3 f1 ef f0 da e9 d7 ce d3 d2 cd d2 ca ca c2 c1 be bc ba b6 bb b1 b0 b1 b2 af b1 ad ac ae a8 ad aa a5 ad a5 aa ab a4 ac 99 8f 8e 90 83 8a 80 7a 75 7a 73 79 71 75 76 7e 75 78 7b 6f 75 7c 74 7c 85 7a 7c 7d 7d 79 7a 7f 7c 81 7f 82 88 a2 ae 93 77 60 42 26 15 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 08 10 17 35 46 50 65 66 75 7a 81 8d 96 95 90 7e 6a 68 6c 6a 6e 75 6d 71 71 73 71 6c 69 6f 73 72 70 6e 7b 73
 87 87 87 90 96 99 a1 a0 9f a5 a1 9e a3 a7 a6 a6 b0 ae aa a7 b4 ac b5 b5 bd bd b5 bd bc be c3 c7 c6 ca d2 e1 dc dc df d9 d7 dc d7 e5 dc d4 e0 e2 e2 e7 ee e7 e8 ed f0 ef fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fa ee eb ea e4 e4 e2 e0 da d1 cd d1 ca c9 c7 c5 bd bd ba b7 c3 b9 bc b1 b0 b3 b2 af b4 a8 aa a9 a9 aa a8 a1 a3 a1 9a 9f 8e 8f 8a 88 87 75 7a 74 7a 77 71 74 74 6b 71 77 7d 7c 7c 75 7a 79 7d 80 82 7d 77 78 7e 7a 7e 7d 7c 7c 78 78 80 76 8c a0 a6 91 74 5f 3b 2b 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 06 14 24 40 47 47 59 6f 74 81 84 84 8e 93 93 84 6b 6c 65 66 61 6e 67 6b 65 6c 6d 6e 6f 6d 70 71 70 78 87 83 86 84 87 89 95 96 95 98 9b 97 97 a4 9f 9e a2 a6 ac ac 9e aa 9f a9 b1 ad b6 b5 b0 b2 be bd c1 c2 ce cb d3 d4 db d5 dc d9 d5 d5 da d3 da da d1 d9 d3 d0 df de e0 e5 ed f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f7 eb e7 e6 df d8 d3 e3 d9 d6 cc c8 c4 c0 c7 c7 c0 c4 bb b6 b4 b2 bb af ad ab ae a6 a5 a0 aa a2 a2 a7 a1 aa 9c a3 99 8e 8e 84 83 81 80 80 83 70 76 75 70 74 70 75 78 78 78 7e 86 7f 79 82 7b 7e 80 81 78 82 80 88 7e 80 79 82 79 82 80 80 93 ab a2 8e 76 54 41 2b 13 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0b 19 2d 43 42 4e 59 5f 6b 79 79 85 8a 8f 8b 71 60 5d 58 64 69 67 6a 6b 6b 6d 77 74 6f 70 79 75 6f 7d 7d 7b 7e 84 8c 8d 93 94 9a a1 98 96 9d 9b 98 9b 9e 9d 9e a8 a7 a8 a7 ab b2 ac af aa b2 b6 bd b8 bc c5 c0 ce cc d0 d9 cf cf d4 dd d6 d6 d7 d6 d2 cf cc d3 cd d1 da de df e2 ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 f7 f0 ef e4 df db da dd da d5 cb ce c5 c7 ca c1 c5 bd bd c3 b8 af bc bb af a8 af a8 a6 9a 9b 9b a0 a2 9c a2 9f 9a 94 8e 90 90 8b 7c 89 7d 7d 7c 7f 7e 79 7e 71 75 79 7d 79 7f 7b 7a 81 84 7d 7d 7e 89 85 85 84 86 85 85 87 85 86 85 80 86 88 a1 a3 a3 90 75 5f 38 25 12 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 04 06 05 0b 20 2a 47 56 55 56 55 60 62 70 6e 79 82 7c 63 5c 54 56 61 60 5e 67 66 5e 61 71 6c 70 73 75 77 7c 79 82 82
 8b 87 89 90 92 91 8e 95 96 9d 9d a1 96 9b 93 9d 9e 99 9c a3 a7 a2 a8 ae ac a4 ae b6 b5 b8 c1 b6 c0 c1 c2 d2 cf cd cd d3 ce ce d2 cd c8 c9 c9 c7 c4 cb c2 c8 cf d6 de eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 f4 eb e8 ef e2 e0 dc d2 dd dc db c7 ca d1 c0 ca b7 bd bc bc b7 b9 b2 b4 b2 aa aa a6 ab a7 9e a3 a4 a1 a1 9b 99 9b 94 93 8b 87 87 82 7d 7e 85 84 78 7d 7c 7a 7d 71 7b 75 79 76 80 85 7d 85 7c 82 87 8c 85 8a 85 86 84 84 88 86 81 8b 85 85 89 89 9a a3 b3 90 6e 5f 36 20 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 06 1e 2a 45 5a 54 57 59 57 60 63 64 6f 69 61 5e 57 54 5a 5b 62 63 64 67 6d 69 6e 6c 71 70 78 89 77 7f 85 7e 8a 87 8b 8c 92 91 9d a4 a4 9b 9c 94 9a 8f 95 9a 96 98 97 9f a5 a3 a5 9d ad ad a3 ae ad af b1 bc bf c1 c2 ca c9 c5 c6 d3 d1 cb d0 d2 c8 c8 c5 c3 c0 c2 bc c6 c6 c6 da f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 ff fb f3 f5 ea f0 e4 e6 dd dc d9 dd db d2 cd d0 ca cc c6 cc c3 bb c2 bb b2 b3 b5 b8 b4 a7 b0 9e a3 a6 9d 9f 9c a5 9e 9f 9b 9e 97 8c 8d 80 89 88 8a 89 8b 86 7b 8d 77 82 74 7d 80 7f 87 7d 7f 83 85 87 84 81 87 7e 88 8a 87 87 8d 8e 82 82 83 84 83 8a 86 8a 9e ac a5 8d 76 58 33 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 05 06 05 0c 16 2d 4d 61 5f 64 60 5d 5a 5e 54 5e 5f 5a 57 55 59 59 5e 5b 60 62 68 67 61 6a 6c 70 74 76 82 7c 7a 82 87 87 86 94 96 91 9c 9c a8 ac 9a 97 93 90 89 94 97 9c 98 98 9d 9f 9a a1 a7 a5 ab ad ad b2 b4 b4 b7 bc bc c0 c9 ce c7 cf cb cf ce d2 c1 ca c1 c0 c3 bf c2 bb bd bf cd e1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff f7 f9 ff f8 f5 f8 f1 fe ef ef ef e4 e6 e6 e7 e5 e3 df dc d7 d5 d3 cf d6 ce c2 c1 c2 c0 b7 b5 b9 aa ad ae aa b4 a6 a1 a9 a8 a1 9e a6 a0 9d 9f 9b 94 9c 97 94 91 89 92 88 88 89 81 83 86 7f 85 8b 79 8b 7e 7e 84 8a 8b 85 7f 89 87 8d 8d 86 8a 8d 8f 89 8d 90 91 88 86 8c 81 90 89 8e a4 a7 af 92 6c 57 2d 15 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0f 10 14 2a 41 56 66 6e 6b 68 66 60 5e 5a 58 55 55 59 60 5f 5f 65 60 60 65 64 6e 70 6c 72 7b 79 81 79 81 81 89
 88 84 8a 90 95 a0 a3 97 99 93 94 8f 92 90 8e 92 90 8f 9c 9e 9c 9a 9c 9e a7 a9 b0 aa b3 b2 a6 b5 bc be b9 c4 bf c6 c6 cb d7 ca cc c2 c6 b6 c6 c6 c0 c1 c1 bb c4 c6 e5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f9 fc f8 f5 f4 f5 f0 ec f4 eb ec ea f5 ec e9 f2 eb e4 e4 e2 da db de db d7 d3 da d6 d1 cb cd c9 c9 c0 c5 c0 bd b8 b6 b3 b0 b2 b2 ad ae b0 a6 9e a6 a1 a5 a6 a0 99 a3 91 99 90 97 9f 90 8a 87 87 8b 85 81 85 85 86 84 86 81 85 83 83 83 8c 82 8b 86 88 88 90 8d 8a 93 8f 8d 8b 87 8b 8d 8c 8c 85 8a 8a 8f 99 a9 a4 84 61 47 1f 18 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 0b 29 40 53 68 6f 73 72 6b 5e 53 59 59 51 57 59 57 5b 61 62 61 6a 66 60 6b 6d 6f 70 6e 70 76 81 75 7e 84 81 80 8c 91 93 96 96 88 8b 86 8e 8d 88 91 94 92 95 94 99 9b 9f 99 9d a2 aa 9b a6 ae b1 a8 ae b9 b2 b7 ba c8 c6 c9 c4 cc ca be c0 be ca be c0 b8 c4 bb ba bb ba cc ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e5 e1 d5 d2 d2 d7 ce d1 cd dd dc e9 f0 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f3 ef f3 f8 f3 f4 f0 ee ed ee e2 e6 e5 e9 e6 eb e5 e0 df d8 e5 d9 db dd d8 d8 e0 d0 d5 cd cc cd cd cd c6 c1 be ba bb c1 b8 bb b3 b1 ae b4 b2 a9 ac ac a4 a2 a7 a3 99 99 9f 9a 9e 94 95 97 97 8e 95 90 8a 87 86 84 85 82 83 7f 86 88 85 83 83 89 86 8c 8b 86 82 8b 8d 8a 90 8a 83 89 8a 94 8d 7d 8b 88 8a 8b 80 8a a3 9e a3 84 62 47 1e 10 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 0b 0f 1f 3f 4e 64 6d 7a 7a 75 5f 57 4b 5b 58 5a 5f 61 60 61 67 66 67 6e 71 6c 6d 6f 75 71 6f 72 7a 79 85 88 87 88 8b 93 92 8a 7d 85 81 86 88 8c 89 8c 8d 91 9b 9b 8f 97 99 9f a0 a1 a7 a4 a5 ab ac a6 b3 b8 b7 bb c0 c7 c4 be c7 c7 d0 c6 c2 b9 c6 ca bd c1 bf b5 ba bc c3 d2 ff ff ff ff ff ff ff ff ff ef f1 f1 e8 d9 c0 aa aa a2 a3 94 95 96 9d a1 b0 b8 bf c4 d1 d3 e0 e9 f9 ff ff ff ff ff ff ff ff f8 f5 f1 f4 e5 e7 e4 e6 e8 e4 e4 e2 e0 db de db e1 d6 d7 e0 d7 cd d1 d2 d5 d3 d2 d0 da c7 ca d1 d0 cd c3 ca bf bd c0 be bf ba bc b5 b6 b5 a8 af ac a9 ac af a9 b0 a0 9f a2 a6 a0 9d 9f 98 99 94 94 9b 92 93 87 8d 8a 91 91 83 87 82 88 83 8a 88 8c 8b 8a 75 88 82 85 8d 88 8b 8e 8d 8d 8f 89 89 8f 89 87 89 8f 8c 8a 81 8c a6 ac 9a 7e 58 39 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 1c 20 3c 53 67 76 79 7a 7f 6a 63 5c 56 57 5d 5d 62 60 69 6c 68 71 6a 71 6f 69 73 78 70 77 80 7b 7e 80 86
 89 90 96 92 8e 82 7c 7f 85 87 87 85 88 8a 89 8e 8f 93 96 a0 9d 9e a2 9e 9f aa a4 a4 ac aa ae b4 b7 be bf c2 bb c3 c6 c1 cd c2 c8 c6 c0 be bd b3 bd af b7 c1 c3 e6 ff ff ff ff ff ff ff f7 db c6 c0 c5 c2 a0 93 85 82 7b 72 74 76 75 7b 75 7f 8e 88 91 9c aa b4 c7 d3 e1 f5 ff ff ff ff ff ff f2 e9 e5 e1 e5 dd dd e3 d7 dd d9 d6 d1 d7 d0 d6 cf d1 d4 ca d2 d1 cc d6 cc ce cb cc cd c6 c8 c2 cc ba c4 bf be c0 be bc be bc bd b5 ab b1 a2 ae b3 b0 a7 ae a8 ab a0 aa 9e 9f 9b 9c 94 9c 9d 91 9c 95 90 94 8d 86 8d 85 86 85 8d 85 82 84 8a 8a 8a 88 8f 89 8a 84 8a 86 8d 8e 87 8d 92 91 95 8f 8b 8f 87 86 8d 86 85 86 9e a4 a0 93 76 5b 36 15 0b 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 06 0c 0b 20 38 4c 68 77 7d 84 7e 79 66 62 57 59 65 5a 5d 61 62 6b 66 66 70 6c 6d 76 74 75 71 6c 77 75 7d 7d 82 7e 81 89 93 90 84 7c 79 6d 75 79 84 79 85 92 8a 91 91 90 9b 9c 9d 9f a2 a5 a0 aa a9 ae ae b2 b3 c2 b2 b7 b8 bc bd c4 c8 c5 ce c2 c1 c0 c8 b6 bb ba b9 ae bc c5 fb ff ff ff ff ff ff ff ef bf ae a8 96 89 79 69 61 6a 64 5b 5c 5e 58 58 5f 5c 65 63 64 7a 8a 8c 91 9e b6 ca ed ff ff ff ff ff da df dd dd df d9 d0 d7 d1 d0 d0 d1 d4 d2 c9 cb ca c8 cb cc cf c8 cb c4 c5 c8 c3 c6 c6 be c0 c2 c1 c3 c2 b5 ba b8 bc be ae b7 b1 b9 b4 aa a4 a9 ab ab ab a9 ae a0 9f 98 a4 a1 98 95 8b 94 96 95 97 92 8f 95 84 87 80 89 88 86 8c 82 8c 86 7b 87 7f 82 88 88 89 8b 88 85 89 86 80 8e 89 92 89 93 8d 91 84 87 84 86 8d 87 9a a3 a1 91 75 4a 24 20 08 0a 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 07 15 20 45 52 6b 79 82 80 89 8d 83 69 67 57 5a 58 62 63 6b 66 6e 6d 70 6f 6c 70 6d 7a 76 70 7a 75 7f 80 7b 84 83 85 a0 9a 88 7f 7c 77 80 79 7d 7f 84 8c 8c 96 95 8a 9b 9a 97 9f a3 a8 a5 a0 af ae b2 b4 b4 be b1 bb be c4 bc c5 c4 c2 ce bb bd bd b6 c1 be b5 be b7 bd cc ff ff ff ff ff ff ff e9 c6 a2 90 88 78 64 60 5f 55 56 5f 50 4f 51 4a 53 52 56 51 4d 3e 60 6c 6e 72 82 8b a6 bb e1 ff ff ff ff df d8 dc d2 d9 ce cf d5 c4 d0 d0 c8 cb c6 ca c8 ca c8 bf c4 c1 c3 bf c7 c6 c4 c8 be b7 c8 b9 bf bf bf c2 b0 b9 ba b0 b2 b5 b8 b6 b2 b3 ac ab ab ac b8 ae a7 ac 9d a0 a1 a2 99 9d 9a 96 94 94 95 90 8b 87 89 8a 86 84 87 86 80 7f 80 82 85 82 87 7e 7e 7f 83 86 86 84 82 84 87 89 89 92 94 8c 96 8f 8a 86 88 86 86 84 88 9c a9 a7 94 72 53 32 1b 0c 07 06 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 08 1a 1b 38 5f 63 71 7f 83 97 92 91 78 64 66 58 58 62 6a 66 70 6a 6d 75 6c 6e 71 70 76 6f 78 79 71 7d 82 76
 7e 7f 87 99 9d 89 7e 75 6f 80 75 79 82 8c 89 90 8a 94 8d 96 95 9a a0 a4 a7 a1 a4 ad a8 a6 b4 ba ae b8 ba bf bf c1 bc c0 ca b7 c2 c0 bc bf b6 b9 bc bd b3 b9 d3 ff ff ff ff ff ff fe cd ac 8a 82 69 62 5e 50 48 4b 4e 49 4b 47 40 3f 3b 47 4c 44 41 2a 49 55 62 59 68 74 7e 8d a3 da ff ff ff e1 d9 cb ca d1 ce cd cf cc c3 c1 bf bf c3 c6 c6 c4 bb c6 be c4 c7 c4 c0 ca be c9 c2 be b9 b9 b8 bc bb b4 b0 ad b7 b2 af ac b0 af b0 b1 a8 ae ab ae ae a4 a9 a8 98 9c 9c 97 99 98 90 96 93 91 91 8e 90 8b 85 84 7f 7d 87 7c 79 78 7e 8a 7b 77 79 7b 80 80 7c 80 7f 7a 7b 85 86 84 87 87 88 8b 8a 8b 8f 8e 8a 84 88 85 8e 94 b0 99 92 6b 4e 30 21 0c 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 11 0b 21 38 5a 61 77 86 84 95 96 98 91 6e 68 5c 5c 5e 5e 6a 6d 6b 70 6b 6b 6f 68 6d 67 6f 71 6d 72 6c 78 6d 76 7a 85 85 8a 82 7b 75 79 7e 76 7c 84 81 87 8a 86 90 8d 8e 8b 99 9a a3 a0 a0 a6 a5 a3 a5 b2 ae b9 b5 b5 c0 bb bb be bd ba bf b8 bb b9 bb b9 be bb b7 b5 be cf ff ff ff ff ff ff f5 b2 90 70 5f 53 56 47 4f 43 3e 40 36 3e 36 2b 34 35 32 33 3b 3a 37 40 42 45 47 53 5e 6a 79 87 ae e0 ff ff de d0 c9 c9 c4 be c1 c2 c5 c2 c2 b4 bf b3 be c2 c3 b9 bc b7 bb bd bf b7 b7 c2 b9 ba bc b1 af b3 ac ae b0 aa af b4 ae aa aa a7 a4 a9 a6 a9 a6 a9 a8 9f a5 9e 9f a0 9b 8e 93 8c 8f 90 90 86 81 7c 8f 85 85 89 79 7a 7b 78 7b 7d 7f 7c 7e 6e 70 74 70 7c 76 76 84 73 7a 80 7b 7d 82 80 84 8e 87 95 89 8d 8a 89 8e 7d 82 8c 9b a5 9e 91 6b 58 3c 22 16 11 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 0c 18 26 40 53 66 72 82 92 94 9f 9c 9e 7a 67 62 60 5f 64 5f 66 67 67 6e 63 6c 6c 70 74 72 76 74 6c 70 72 73 73 70 74 82 85 85 78 75 6f 6f 78 76 7a 80 83 81 87 8a 95 98 92 93 9b 94 aa 9f a6 a9 aa a9 a6 ae ac b1 b9 b7 bd ba b6 c0 bd bc c1 bc bc b6 b9 bc b9 b2 b8 bd d3 ff ff ff ff ff ff da 91 7a 66 55 41 49 3e 39 3b 39 3a 36 2c 27 27 2f 2d 2d 2e 34 34 33 39 3a 45 42 45 52 5d 67 70 94 be f5 ff db c3 bf c0 ca c3 c2 bb c0 bf bd b4 ba b8 b9 ba b5 bd ba b3 b5 b4 bc ba c2 b9 b3 ab b6 b9 aa ad b1 aa a7 a1 a8 a2 ab a8 a9 a6 a2 a5 a6 a9 98 9d a4 9d 99 a1 98 90 95 99 8a 93 93 89 86 80 84 8d 80 7e 78 77 77 78 7b 7b 77 6f 74 7a 79 77 6f 7c 6d 76 72 7b 76 75 7b 7c 85 81 83 78 7e 83 8b 8b 87 87 82 8c 86 80 84 80 9d b0 a1 91 6e 5a 47 2a 1b 07 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 10 1b 2d 44 51 6e 7b 88 92 99 a9 a5 9e 8b 6a 64 5e 62 68 6a 6d 64 6b 68 65 6a 68 6b 6c 6e 76 71 78 68 70 76
 72 77 7e 84 87 6f 76 6d 73 72 76 78 75 81 76 83 85 87 95 8c 8f 9c 9e 94 9c 9e a0 a2 a8 b0 a7 b4 af af b0 bd b8 bb bf be c2 ba c1 b8 b9 b9 bb b9 bd af ba bc d1 ff ff ff ff ff ff bc 75 63 54 4a 3e 40 3b 28 31 2f 33 28 23 20 23 26 24 22 1e 2a 2d 29 2b 35 34 3a 41 45 4d 51 5a 81 ab d9 ff dc c2 c2 b8 c3 bc b5 b9 c5 bd bc b3 b9 bc b5 ba ba b8 b7 b1 af bc bf ba b9 b3 b4 b1 b4 b0 ac ab a9 ae a1 aa a3 a6 a4 a8 a5 a3 a4 a3 a1 9d 9f 9c a1 a0 a3 9f a0 96 90 96 89 8f 87 7e 83 80 8b 86 86 82 7c 7b 77 77 70 76 7b 69 7d 72 75 74 73 6a 74 70 79 73 76 74 79 73 70 75 7c 7c 81 81 7f 8b 82 85 83 81 82 84 7e 8b 9f b2 a2 87 79 5e 49 2f 20 11 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 18 31 3d 53 6d 74 86 8f 98 a5 ab a3 89 69 58 51 59 63 68 6e 66 63 5f 62 64 62 64 69 64 73 6d 66 71 6d 73 7b 83 86 78 72 71 6d 70 7b 6f 7a 78 74 74 75 84 7d 83 85 88 86 91 96 91 97 93 9d 9e aa a2 a0 a9 ae af b3 b1 ba ad ad bb b6 b7 bd bd ba b1 b8 ba b2 b3 b5 bf c9 ff ff ff ff ff da 94 70 5d 49 41 3f 3d 30 27 24 21 1e 1c 23 20 20 1d 16 1f 21 1d 23 23 22 2a 30 2c 34 3a 3d 44 61 6f 8c d0 ef db c6 bd ba be b7 ba c4 c2 bb ba b6 b9 b5 b1 b1 b2 aa b4 b1 ae b3 ac b5 b8 b8 af ab ad ab a5 a9 a8 a9 a7 a6 9a 9f a5 a6 a0 97 9e 9d 95 91 9c 93 99 9a 92 8f 98 8c 8d 8e 85 86 84 85 80 7f 7b 85 7a 7d 7b 72 72 71 74 72 69 72 6f 77 76 67 72 66 73 73 6f 7b 70 6d 6f 71 75 75 77 81 83 81 7e 7f 85 84 85 81 82 7f 7c 85 97 b0 a3 97 7b 5b 48 2a 1f 14 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 09 16 1e 38 4f 5b 71 78 88 94 9f a8 a9 a9 91 67 67 59 5c 61 61 63 5f 68 64 61 62 6b 69 68 66 6d 6c 6d 74 7a 7a 81 7f 76 6d 76 73 6c 6d 73 72 76 73 6f 77 73 7c 7b 7f 85 87 88 8e 95 96 92 92 96 9d 96 9b a4 af af ad af b4 b0 b4 ae bb b6 b5 b0 b6 b0 b5 b6 b6 b9 af b5 be cc ff ff ff ff e3 b5 89 65 4e 40 30 30 2c 22 25 1d 1d 24 21 1e 1b 12 15 11 17 1b 23 1b 1a 1c 21 28 22 31 31 30 42 4f 62 83 ca eb d3 cb be bc bb ba b9 ba bf b8 bb b2 b8 af ba b4 af ab aa ab b5 ab ad ab af ad ae aa ab a9 a6 a9 a8 9f a4 9d 98 9d 9c 9b a0 97 96 9e 9a 99 99 9a 9a 9d 8d 8e 96 8b 84 8b 84 87 81 7b 7c 71 7d 76 7e 78 72 78 73 6e 6f 70 70 6e 6c 69 6c 6e 6f 6f 70 77 73 73 6e 6d 6b 6a 6d 73 7b 76 7f 79 77 81 83 84 7b 88 7d 73 7e 7d 9b ac a7 98 89 69 4f 3b 26 19 04 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 07 06 05 1e 24 34 53 67 6a 85 86 91 a0 ad ab ad 95 6a 5e 61 60 64 66 62 5c 65 62 5f 5a 66 67 67 68 6b 74 74 76 82 82
 79 78 72 6b 74 6f 72 7d 72 7a 76 70 73 7a 81 7f 7e 7c 86 85 87 87 86 8b 8d 8e 97 94 90 9f 9a a5 a7 a1 aa ae a8 ae ad b2 b1 b0 af b5 b8 b3 ad ad b4 b4 b7 bb c4 ed ff ff f1 c5 9b 7d 59 51 36 31 2f 23 21 1c 1e 17 15 17 1a 16 12 14 0d 14 1a 0e 0f 16 18 1b 24 24 28 21 32 36 49 61 7b bd e1 cd c4 bf c0 be bd b9 b0 b7 b1 b4 ac bc ad b8 b6 a9 b3 ab ad a6 ae aa a8 ad a6 a0 a4 a9 a0 a0 9e 9f 99 9d 9e 96 94 9b 9b a3 99 98 93 95 93 95 98 94 9b 89 8b 8a 83 8f 7f 7f 7c 7d 7d 76 74 7d 78 78 74 75 71 79 69 70 72 75 6e 72 6b 72 69 70 73 6f 68 6b 72 79 70 6d 6d 6f 76 76 76 77 81 7a 85 7b 7a 7c 7e 89 7c 7e 7a 9a b5 ad a0 89 71 52 47 28 1a 12 06 05 06 04 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 1a 29 33 54 65 7b 86 90 92 a0 a7 ad b0 91 63 60 5d 5e 64 68 65 59 60 61 60 64 66 6a 61 62 74 72 79 7a 76 73 76 6b 78 67 6f 71 7a 75 6f 75 70 70 76 76 75 7d 76 75 85 84 88 82 8a 82 88 8e 95 8e 96 95 9c aa a6 ac 9f b1 af ac a5 ac af b1 a9 b3 a8 b4 b3 ba b4 b3 b9 bd c0 dc ff ff de b5 8b 70 51 48 2c 20 26 1e 15 17 0d 15 0a 14 0d 10 0c 09 15 0c 11 13 11 10 11 13 15 24 24 24 26 21 38 5e 80 ba e2 c9 c3 bb b0 be ba ae b6 ad ae b7 ae b9 b4 aa ac b0 ae b2 a6 aa a4 a6 ac a5 a4 a2 9d a5 9c a2 9a 9d 99 97 95 97 99 97 8e 90 97 92 95 95 8e 91 97 8b 8b 8b 8a 90 85 86 89 82 7a 79 79 72 7b 76 72 78 73 78 75 6e 6e 6b 6e 65 6a 6c 6b 73 6b 6b 66 6f 64 6b 73 6a 6a 6f 6d 6d 6d 70 71 7a 78 73 7a 7e 7c 78 7e 7e 7f 7b 80 93 ab ad a4 84 71 5a 44 35 1f 13 07 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 12 14 20 25 39 53 67 73 80 96 91 a1 b0 b1 ad 94 64 5e 52 5b 5e 5d 61 60 5c 5a 5c 5e 68 68 6e 71 68 70 6e 6e 6c 6e 69 6c 70 69 6e 79 75 78 77 7c 77 73 78 78 77 7b 73 7f 78 84 79 86 8a 8c 93 8e 85 8d 8f 95 94 94 a3 a9 a2 a1 a1 a2 ac a5 b3 b0 ae aa b0 b0 b0 b4 b9 b8 b6 b1 bc d8 ff ff da ad 88 69 4b 34 2b 23 15 15 13 15 12 14 0f 12 0f 10 0b 0b 0d 0c 06 11 0c 0f 13 11 1c 1e 1d 1d 20 27 35 54 80 be d5 c4 b7 b6 b6 b1 b8 b2 b5 b8 b0 ae ac af ac ab a9 ad a6 a6 ae ad 97 a0 a3 9f a1 9a 9a 97 9c 92 95 98 96 95 94 94 98 95 95 91 93 9a 92 93 8f 93 94 90 8f 8b 86 82 80 87 7f 7c 76 6f 76 7a 74 74 75 77 6e 6f 6b 74 69 6d 76 71 69 65 63 6d 6f 73 6b 6b 68 6d 6c 6b 6a 61 6f 6e 70 6b 73 75 73 78 76 7d 72 7b 7e 7b 7c 78 84 89 ac a5 a6 8c 70 5f 3b 33 1f 18 0f 09 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 0f 1a 27 34 4c 64 6a 74 8b 94 9e ac ab ba a4 85 66 5d 60 60 62 5f 5f 66 64 64 5e 65 65 6d 6d 6f 6c 6f 6c 6c 67 66
 6e 6c 6b 72 66 6e 77 71 76 75 77 7a 78 7a 76 79 7f 79 81 80 7d 81 8b 88 8c 85 85 87 95 8f 93 98 9f 9e a5 ae ad a1 a7 a4 b0 a9 ab a6 aa ae a8 ae b7 af b9 b3 be c2 ff ff d6 a9 85 66 49 3a 1b 15 0f 16 11 08 0f 0b 0f 0d 05 0a 0a 06 09 0b 0d 11 05 02 0d 0d 16 1f 1b 22 22 20 2d 4c 81 c0 c4 bd bc b8 bb bb bd b6 ae b4 ae b6 ac b0 aa b1 ae ac ac 9a a1 a1 a9 9a a3 9d a1 9e 96 99 9d 97 94 9c 92 9a 99 94 90 90 95 8a 91 8c 91 8b 93 90 8e 8c 89 8b 8f 8d 89 7d 7f 75 79 75 6c 79 73 75 68 70 72 74 73 6f 69 71 6e 66 6a 6e 70 75 67 6e 70 6b 7a 6b 72 6b 69 70 70 6c 74 6e 70 75 7b 7a 80 72 74 7d 81 79 78 7a 7b 81 a5 af a5 98 79 69 52 3a 30 21 15 0b 05 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 07 0c 09 24 23 38 4f 5b 6d 81 91 95 a5 a7 ac b5 a3 76 61 5f 53 5f 61 63 61 65 65 6e 6d 74 69 6b 5f 58 62 64 64 66 62 66 6c 6d 6c 69 65 69 68 71 6e 74 7b 78 74 80 78 7d 84 7d 82 77 80 7c 84 7c 88 85 85 8e 84 8c 92 99 9c 9d 99 9a a1 9b a6 a9 ac ac a6 a7 aa a7 a7 ad af ac b0 b2 b6 c3 e2 ff e3 b6 8f 6c 3e 28 13 0e 0f 11 11 07 10 08 13 09 07 06 06 05 05 0c 06 05 07 0a 0c 12 14 13 1a 1c 21 15 2c 47 8a bb c1 b9 aa b2 ba c5 b2 b9 aa b2 aa b7 a9 ad ad ad a5 9c a3 a2 a2 a5 9f a0 9e 9b 9b 90 94 94 8e 90 86 97 8e 92 93 8c 94 98 91 94 8c 92 90 8f 89 8a 8b 89 8a 83 87 85 84 7f 7d 74 68 6c 6e 76 6a 6d 6a 6a 67 69 6e 69 69 69 6a 6b 6d 6c 66 6a 6b 63 6c 69 71 64 63 72 61 69 6e 6e 6b 6b 6e 70 6a 6e 72 75 78 72 7b 74 73 79 78 7f a0 a9 aa 91 7b 67 50 3e 28 21 0f 0d 05 0d 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 12 15 18 25 3e 49 5f 7c 85 97 9b 9d b0 b1 b0 9b 70 68 52 5b 61 61 64 65 6b 6d 6c 68 68 61 61 5c 61 64 65 5c 66 67 69 68 63 69 65 63 62 5e 6c 71 6d 66 75 71 76 7e 7f 83 7e 7d 81 7c 80 80 89 8a 8a 7d 8a 88 8a 94 95 93 99 95 a5 9f a1 9c a3 aa a0 aa a5 a0 ab a6 b0 a6 aa aa b3 b6 bb c8 fc ee c9 95 75 48 2c 1c 08 11 0d 06 0e 03 04 08 0e 03 09 06 05 03 06 08 08 05 09 06 08 0e 0c 14 1b 17 1c 25 45 84 b7 b7 b5 b3 ba be bd be b9 b0 b5 ac af a4 aa a3 a9 9b 9d 9d a6 a1 a1 9a 9d a0 9e 9c 90 92 92 93 91 8f 8e 8d 8a 8f 89 8c 86 89 8c 8e 8c 85 94 8d 85 86 77 86 7d 83 7e 82 80 7d 6b 64 74 6e 6c 65 6b 6d 6a 6e 61 6f 6b 67 6a 65 69 65 67 68 63 61 6f 69 67 6d 6a 71 69 6e 6c 6f 67 70 68 6f 6c 68 6d 6a 6a 6e 6d 76 7c 7a 74 73 7d 90 ab a5 94 7d 68 55 45 3b 2d 19 12 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 05 0e 1f 25 31 41 4b 62 74 82 a3 a4 a5 b2 ab a9 8a 73 66 5f 5f 5d 56 62 63 6f 75 6b 70 5f 5c 58 5f 58 5d 62 5d 66 5e 66
 65 62 62 68 66 68 71 68 65 70 71 72 74 73 78 84 7c 77 7f 83 7b 7f 86 76 84 81 85 84 8b 86 8a 93 94 94 98 96 97 9e 9e a6 a9 a2 a8 ab a2 b0 a5 a9 ad a5 aa b2 ab b5 b8 de f1 df ae 7b 49 25 0d 05 03 08 0d 05 07 0c 07 07 0c 03 06 05 03 09 06 05 06 0c 06 07 0e 17 19 19 13 10 22 52 84 ac b4 b3 b3 b4 be ba b6 b0 b2 ae b4 ae a6 ab a9 a3 a1 9e 9b a0 9d a2 96 9a 96 9b 95 94 96 86 91 91 8c 8f 88 8a 83 86 8f 92 90 8d 87 8b 8f 8a 89 87 89 87 8d 7a 86 88 7c 7e 76 76 70 70 6f 70 66 6d 6a 6a 6f 68 6d 64 60 66 6f 6d 67 68 63 6b 69 69 6a 68 6e 68 69 72 68 68 67 65 6e 68 67 63 67 5e 72 6b 73 70 7a 74 72 77 79 74 89 9d 9f 98 81 74 61 4c 40 2c 2d 18 12 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0b 11 09 1c 30 2a 43 59 6b 7b 87 99 a8 a8 af ae 99 7b 65 5a 54 5c 62 5f 6f 68 6a 72 64 57 5c 59 5c 65 61 62 63 61 5f 61 6c 69 6b 69 63 68 6d 6d 64 78 6e 66 6e 76 74 79 80 77 7e 85 84 7d 7e 80 80 84 7d 7c 83 84 89 8a 8d 91 91 8d 97 98 9c 9b 9c a7 af a4 a8 a8 a3 9e a7 a7 a2 a7 a5 ac b2 ad c6 f1 eb c3 8b 53 29 12 0d 0e 09 06 0a 03 00 09 09 03 06 06 08 03 0a 06 08 07 02 07 07 0a 0a 0b 0b 12 12 1e 4b 88 a0 b2 b7 b3 b3 b1 bb b4 b5 ac a5 a8 a6 a5 a9 9c a2 9e a3 9f a4 9b 93 95 95 8b 95 92 94 91 93 89 84 92 8a 8d 8a 86 8b 89 84 88 81 86 81 83 88 84 8a 87 7d 80 7d 85 7f 6f 70 7b 74 70 6b 63 6b 6f 60 65 6e 6c 6d 65 64 64 67 66 6a 6c 60 6b 69 68 6b 6e 6a 6b 6b 6f 68 6b 6f 71 65 67 6e 64 6d 6c 62 70 72 6b 6f 69 78 72 76 76 78 86 93 9c 94 7a 72 5f 51 3f 37 25 1d 14 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 08 09 1e 25 2b 40 49 5b 71 7c 89 94 a5 a6 b1 a1 92 6f 56 62 60 61 68 61 76 6f 6c 61 61 5d 5a 5c 5d 53 5d 5f 63 5d 5e 63 5d 64 68 5e 67 6d 65 62 65 68 6d 67 6c 6e 71 73 71 72 81 7d 84 82 82 84 7f 83 7d 7e 81 7e 82 88 86 8f 8d 8d 96 8a 97 9e 9d a1 9f 99 a2 9f a1 a1 a5 a6 a6 a4 a8 a0 a5 af b9 dd f1 e2 a2 63 2a 0f 05 05 09 06 05 03 0b 0a 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 0b 11 0e 10 1b 15 4e 7f 9d b0 b1 b8 b9 bc b5 b1 b2 aa a9 aa a9 a2 a1 9a a0 a1 9a 99 9f 96 9a 96 95 99 90 8a 8f 91 8e 88 8c 8a 8b 8a 8f 8c 8c 87 8a 88 84 89 83 83 88 82 7d 7f 7c 88 78 82 7e 76 71 72 6f 6c 6c 65 66 67 65 6a 6c 60 5e 65 6a 68 66 68 63 62 65 64 65 5f 65 66 66 6b 5d 67 6e 6c 67 65 63 6e 61 69 70 64 67 65 6a 62 70 6b 68 76 6f 73 71 76 8c 92 98 7f 73 63 54 53 36 29 1e 0f 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0b 19 14 1f 2c 38 50 62 74 86 9a 9e a4 9e ac 98 84 61 5f 60 59 67 6a 70 71 6d 64 60 5b 55 56 61 57 5e 64 62 5c 66 5d 68 64
 64 67 64 65 6c 6f 65 71 6a 65 6e 6f 70 70 71 72 6e 79 82 76 81 89 83 7d 7b 80 80 82 87 88 85 89 87 90 8e 8e 8e 91 94 95 9c 9d 97 9c a0 9f 95 a2 a4 a0 a2 a5 9e a7 ac aa ba ce ed c4 75 2d 12 07 09 04 06 16 04 01 0b 05 03 00 06 05 03 01 06 05 03 00 06 05 0c 0b 11 0a 13 1d 1c 41 79 a7 b6 b4 b5 b5 c2 b9 af ad a0 a2 a3 a5 a4 9f 9f a3 a1 9e 98 9a 8f 95 8e 9a 90 93 8f 8e 8b 8f 86 89 84 89 8c 8f 8a 8a 8c 87 8e 86 8d 83 80 84 80 7f 85 7c 85 7b 76 83 7c 74 6b 6a 6e 64 73 6e 61 64 66 72 63 68 68 61 63 6a 69 63 66 6b 6a 65 64 60 67 6e 65 71 67 6e 6a 64 68 60 6f 6a 6d 63 62 61 6d 61 6c 6b 74 70 6a 74 74 6b 73 7d 86 90 81 76 6b 55 45 3e 2e 1d 0f 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 08 0d 10 14 1f 35 44 52 64 78 82 92 aa a5 a3 97 7a 6c 66 5e 64 5a 66 74 6c 6c 63 59 5e 58 5a 5f 57 56 65 59 65 60 5a 5f 67 66 61 6a 66 69 6b 61 63 69 73 6e 6c 71 70 6a 70 73 6e 79 75 84 81 81 81 7a 80 78 82 82 7a 87 83 86 8b 84 89 90 8d 98 96 99 9d 92 8d 99 92 9f 9b 97 98 98 9a a7 9f a3 ab a6 aa b6 d5 d4 8b 34 0d 10 03 01 06 07 03 00 06 09 05 00 06 05 03 00 06 05 03 00 06 0a 03 07 06 0e 14 18 1f 32 7e 9e b6 bf bb c2 b3 b2 ad ad ad a5 a3 a2 a0 9e 9c a4 9a 9b 98 a0 95 98 92 91 9a 90 90 8b 8b 8f 84 8d 8c 88 81 8b 85 80 8b 85 89 84 81 84 85 86 89 81 82 79 81 7c 7b 7b 71 6f 70 70 66 67 69 67 68 69 69 69 62 61 69 69 65 61 5e 65 62 6a 64 66 62 70 62 6b 68 64 6a 6c 69 64 65 64 67 69 5e 64 64 60 6a 5b 63 65 66 6e 71 6d 72 72 71 74 79 84 85 7b 67 67 5a 4c 36 28 16 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 07 06 13 1d 31 36 40 54 68 80 90 99 9f a6 91 82 6d 5a 69 62 5d 68 6a 72 6c 68 63 5c 62 58 55 55 60 69 57 62 61 62 57 5f 6f 68 65 6c 6b 65 66 6a 6b 62 6d 6b 68 67 6d 70 71 6c 72 70 78 7a 7c 84 76 7d 80 81 7e 81 76 72 7d 7e 85 85 82 90 89 8d 99 95 91 91 89 8a 97 8b 96 9b 9c 9c 9c 9e 9e 9f 9e a5 a0 a8 b1 c2 9e 3a 0d 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 0a 0b 14 2d 78 a4 b7 bd b9 b1 af b3 a9 a5 9b a0 a1 a1 a1 9e 99 97 99 9f 9b 95 98 95 8b 91 8d 8c 8f 86 88 87 86 89 85 8b 80 86 80 80 80 8a 7c 81 84 81 7d 76 78 77 76 80 75 7b 76 7c 6e 70 70 63 63 66 60 65 62 62 66 64 62 62 68 5f 5b 64 61 67 6c 61 67 69 64 6c 63 68 67 6e 67 67 60 62 64 66 66 6a 65 5b 5d 63 5f 64 68 69 67 6a 69 6f 75 70 6c 6a 78 78 79 78 6c 60 51 4e 39 28 1a 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 06 13 1a 25 34 42 56 6b 84 98 9c a4 9b 74 67 5d 61 66 62 64 6d 6d 6c 63 65 63 60 63 59 57 5b 5f 60 59 5d 58 67 63 65 72 5f
 63 69 67 62 71 61 6d 6c 6c 7a 64 69 78 72 75 6a 6d 73 74 77 79 77 81 7a 7d 7d 7f 84 7c 84 7e 77 84 82 87 8b 8c 90 94 8c 99 91 90 90 95 92 8d 90 96 9e 9a 9d 9a 94 97 a1 a3 9f ab 9b 88 3b 0c 06 0c 06 06 05 06 00 0b 05 04 00 06 05 03 03 06 05 03 00 08 08 04 02 06 0e 15 10 0f 35 6d a9 bc c3 c0 ab ac a8 a7 a1 9d 9a a8 9e 9d 9e 9d 9e a3 91 97 99 9b 8f 92 89 8a 8f 8c 90 89 89 8e 80 7e 85 86 7d 85 84 81 80 81 84 88 83 82 7d 80 7b 74 7c 77 77 7e 76 73 69 69 6f 67 61 65 64 64 65 6a 5e 6b 61 5d 5f 59 5f 62 69 64 66 60 63 5f 60 68 64 6a 63 67 74 67 67 65 58 67 5f 66 62 61 66 61 65 63 60 69 69 69 6a 70 70 6c 66 68 71 73 76 77 65 5d 54 42 29 18 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 08 14 17 1a 2b 37 49 5a 76 84 97 9f a4 8d 74 65 5f 58 66 63 70 73 68 6b 67 63 66 5c 56 5d 60 5c 66 62 68 60 5e 66 62 61 68 67 68 6c 69 68 64 6c 64 69 6f 6b 71 6f 6e 6f 70 6b 73 76 79 6f 72 78 76 7f 7a 78 7e 7d 7e 77 7a 7b 81 82 88 8c 88 8d 94 93 92 89 92 8f 89 92 8f 8e 97 87 9a 93 a4 9d 99 97 a0 9c 9a 93 7f 45 12 0d 09 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0f 07 0e 10 11 22 66 9f b6 b5 b0 ab a6 a3 a8 a0 a3 a1 9d a3 a3 9c 94 9c 9e 95 95 98 8a 97 8b 8e 8f 86 90 8f 84 8a 82 8b 83 86 83 81 89 84 82 85 85 84 81 7f 85 7d 84 7b 75 7a 7e 78 76 7a 67 60 6d 66 62 67 61 64 68 64 63 6e 69 64 65 64 62 5c 65 67 62 68 63 5d 66 6e 60 68 64 6d 5d 63 60 65 67 63 60 60 6c 65 5c 5e 5f 5e 65 60 65 5e 65 6c 6a 6d 6e 72 62 6d 77 79 77 6c 62 4f 4a 33 20 19 09 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 07 15 25 2a 3a 54 5a 70 7f 93 a0 96 79 6b 60 61 67 69 6b 66 6f 66 5a 66 63 5f 66 61 5b 5c 5d 5c 5c 5e 61 65 69 67 5d 65 6a 68 64 65 69 65 6b 66 6f 67 6b 6f 6d 6c 6e 73 6e 72 6c 6b 6e 6e 7a 79 74 7a 75 72 75 73 79 7b 80 7e 7a 81 84 89 8c 88 88 91 81 86 87 83 8c 8a 91 97 90 8e 96 92 90 95 93 93 90 94 8a 7b 42 0d 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 0d 06 04 0f 13 1b 5d 98 af b3 b1 a1 a0 a3 a2 96 a3 94 a2 96 93 94 8d 9a 95 95 96 92 91 85 8a 87 89 91 88 81 82 7d 83 85 80 84 7d 7c 7f 80 7d 7b 81 84 7e 76 81 82 78 79 7c 72 7a 72 6b 75 68 6b 6a 65 66 62 64 66 5c 6f 62 62 64 5f 63 5e 56 5f 5b 65 5f 5f 65 67 62 65 5f 60 63 61 65 62 60 64 5c 56 58 5c 5f 62 58 5d 5c 5f 58 5f 61 5d 63 65 6a 69 66 69 5e 63 6b 70 7d 71 65 59 4c 3b 21 10 0d 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0f 11 19 2a 40 53 5d 6d 84 9d 9c a1 7f 6b 6c 65 6b 7a 6f 6c 64 61 5d 63 5d 6d 65 5e 61 5f 63 5e 64 5d 60 5b 64 5f 6e 6c 65
 68 6c 6c 68 6e 61 6d 63 65 6f 66 6a 6f 6a 67 71 6e 6b 75 6c 77 74 75 76 7c 7b 77 7c 72 7c 82 83 7e 80 81 86 8b 89 89 8d 89 86 82 84 86 81 85 86 8c 94 8f 8c 8b 92 88 8c 8a 8b 95 87 75 4e 0b 05 03 00 06 05 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 0b 11 13 20 53 95 b2 b0 a8 ab a1 9c 9c 9c 99 9c 97 8d 8e 96 8f 9e 94 92 92 8d 8b 91 88 80 86 7e 86 8a 85 86 84 7f 7c 82 84 7b 85 84 79 82 84 79 83 80 82 76 78 72 74 74 78 71 74 71 68 61 63 64 61 62 5a 66 67 68 60 67 62 68 61 59 59 60 5b 56 5f 60 60 61 5b 67 61 63 62 61 5e 62 5e 5f 5a 5c 5e 56 60 60 5e 5d 5d 56 5c 57 5d 5b 61 67 67 6b 6b 65 62 62 69 74 76 78 63 58 49 34 23 16 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 1a 16 22 34 4a 4d 67 76 8f a1 a7 90 79 68 70 71 79 7f 75 6e 6a 65 5d 5c 66 64 62 5c 62 5a 5f 6d 62 5e 6c 68 6f 68 6d 6f 6d 64 66 6b 65 6c 6a 65 67 66 69 70 67 6e 67 6e 6f 73 6d 6c 6f 64 6f 73 75 7c 7b 75 79 78 70 79 7f 7b 76 83 88 86 83 87 84 87 86 7e 84 83 8d 81 85 8d 8d 91 8e 8b 8f 87 8b 93 85 8c 84 78 4a 10 05 0a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 10 15 14 28 49 83 a6 a2 9e a9 99 a1 9d 99 93 92 9c 98 93 8c 8e 96 93 8b 92 96 95 92 8b 84 88 8d 85 85 7f 7f 81 83 89 7f 80 81 7e 84 75 81 7e 80 83 7d 83 7e 76 74 76 7b 7b 73 75 73 67 68 66 6a 60 5f 6b 62 65 5f 65 60 67 68 60 63 62 60 67 60 5c 61 65 5d 5f 61 5d 5f 64 60 5f 61 60 61 5e 60 62 5f 62 65 5f 5e 5d 55 58 5b 5e 64 5b 64 6b 64 66 60 5d 58 6a 73 72 76 6d 52 49 36 24 1a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 10 06 14 26 2e 46 5b 6b 84 90 a3 a6 8b 7e 70 7f 7e 87 85 79 71 69 61 5d 65 61 64 66 64 5b 5c 5e 62 68 64 68 69 6a 63 67 6d 65 61 70 67 61 6a 6f 64 69 6e 6d 61 62 67 69 67 69 70 65 64 6b 6a 6a 6b 78 7b 76 76 78 76 7a 7c 79 7d 82 7f 87 85 81 80 82 7e 76 75 7b 81 79 88 84 8d 89 86 79 84 8a 82 84 89 81 84 81 6b 4c 1b 10 03 00 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0f 0b 0d 10 11 1b 40 86 99 a6 a4 a2 9b a3 97 90 93 95 92 91 90 96 93 96 93 8e 91 8f 8a 89 89 8e 8c 87 8f 89 7e 7f 7a 7e 82 80 82 84 80 7a 85 80 84 80 7b 82 76 7b 76 70 7a 75 75 6b 6c 71 65 67 68 57 5b 60 62 67 58 5e 5f 62 59 6a 58 5e 58 59 65 60 5d 5d 62 5f 5c 5e 54 60 5b 61 5e 5e 5f 5e 61 5d 5c 59 5e 61 5b 5d 56 59 59 5d 5b 64 57 5e 64 66 68 5f 65 5b 62 70 77 80 6e 65 4e 3a 27 1b 0c 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 11 22 28 35 4b 50 6a 82 99 a2 a4 99 82 7a 7d 85 8b 88 79 6c 5b 5f 66 69 64 65 5f 61 60 66 62 66 65 65 67 68 65 67 67 61 68
 65 61 68 64 63 65 62 65 67 65 66 5f 68 6b 6a 6e 6c 60 66 6f 64 6d 6a 64 7a 6e 7b 70 76 78 76 79 83 80 80 82 75 7a 82 76 74 80 7d 84 7c 82 7e 75 85 82 84 87 87 8a 88 81 7e 81 7f 7e 79 46 19 0b 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 08 05 07 0b 06 14 35 7e 9a 9f a3 94 96 8f 93 91 93 8c 97 8f 87 8d 90 95 88 88 89 88 92 8a 8b 81 8c 8d 82 7b 83 89 7e 83 73 80 7a 81 7d 7c 87 77 7a 7d 7d 80 7e 7f 77 75 70 7d 74 73 6e 66 64 5b 5f 60 62 67 5a 64 5e 62 5f 65 5f 5a 61 60 5a 5e 62 5c 62 5d 57 5c 54 60 5d 5e 60 5e 62 58 64 4f 55 60 58 51 5f 58 4c 5b 60 51 58 5a 5d 5e 58 67 66 65 62 62 59 5d 64 73 76 78 70 65 51 43 2d 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0a 23 24 41 51 5d 6a 80 9c a0 a4 8b 83 7c 77 89 8b 83 77 6b 66 5b 62 68 64 63 64 62 63 61 64 66 65 65 64 68 64 61 68 68 64 66 67 68 63 6b 6d 71 66 68 66 69 68 67 6b 60 63 66 72 6f 69 63 67 64 74 6d 75 7d 74 74 7d 79 83 7b 81 83 80 7d 7e 7a 77 77 76 7f 7e 80 81 78 7a 84 7b 7e 80 84 8a 80 84 88 8a 85 82 77 4e 15 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 09 07 09 0c 10 16 31 6f 94 94 9a 94 93 94 92 96 88 85 8e 8d 8a 89 8a 93 8c 8a 8b 87 87 8f 83 86 86 84 84 7e 7e 7e 7b 7c 79 86 7d 7b 81 79 7f 83 80 79 7a 7a 74 79 77 79 78 7e 7d 72 70 64 5f 62 64 5b 63 5c 69 5f 5e 64 5d 60 59 5e 62 61 60 58 62 5c 61 64 5f 5e 4f 5f 5a 5c 56 5d 56 5a 56 57 5b 5c 59 5c 58 5b 5d 60 65 5a 5c 56 60 5c 5d 5e 5a 64 6c 64 67 64 5e 70 76 7c 73 60 51 41 33 27 0b 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 14 21 2a 3a 4f 5f 77 86 9c 9c a2 88 84 72 7a 7d 84 8a 7e 6e 64 5d 60 67 67 69 63 65 67 65 60 67 63 66 6e 64 68 66 5f 65 63 61 60 69 63 62 6b 61 67 6a 6f 6b 64 65 67 6a 65 69 63 69 65 61 66 68 6d 67 66 76 76 75 70 7b 7f 84 82 78 7e 75 80 6b 7b 78 71 75 78 79 7c 7c 80 82 7e 82 7b 81 84 87 8b 86 81 85 80 77 60 19 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 16 07 12 2c 66 8a 97 96 98 96 89 83 84 8f 89 8a 83 88 88 85 88 86 88 87 89 89 87 87 80 82 84 81 7e 7f 84 7f 81 78 83 77 86 83 74 81 7b 80 82 80 7a 77 7b 76 77 78 71 7b 71 6f 62 61 61 61 5f 65 5e 5c 55 58 60 5e 5e 5a 5e 5f 5b 57 56 59 61 59 55 5a 56 59 54 5f 59 5d 5b 5b 61 55 5f 5e 57 5a 5a 5a 57 5c 59 5b 56 59 59 58 5e 5f 60 61 65 68 64 65 57 60 6b 7a 7a 6d 61 58 43 33 20 0e 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 13 0f 1d 2e 3d 4d 5c 7a 85 9a a6 99 8b 79 79 80 6e 77 7b 77 6a 69 65 64 5b 66 61 5b 6e 61 65 5f 62 65 66 6c 66 68 6c 64 61 65
 62 6e 69 65 5e 66 62 5e 66 62 63 69 68 5c 6b 6a 64 6b 6a 71 65 64 68 63 66 73 6f 70 7c 7b 7c 7e 7f 77 7e 7a 72 77 74 6f 73 6f 76 7e 70 7c 79 80 75 73 82 87 83 8b 8a 7b 7e 82 83 84 74 60 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 08 05 06 0f 28 5b 93 96 9b 94 93 94 89 89 8a 87 8b 88 88 87 8b 7d 83 87 87 8e 8a 86 88 8e 84 86 7d 84 77 81 74 82 79 7e 76 80 85 7d 86 80 7c 83 73 7b 7e 76 7c 71 7d 79 76 71 71 64 62 61 63 63 62 60 56 5c 5a 5e 5d 67 5a 51 55 57 59 5f 55 54 5b 5a 59 56 52 59 57 55 5e 61 55 57 53 57 56 5a 56 5f 56 55 5a 57 56 59 58 5a 4f 5b 54 61 5d 61 63 60 5c 5c 5e 71 75 7e 74 63 57 45 35 28 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0f 14 22 2c 42 5b 64 7f 8c a0 a8 9e 7b 75 75 72 7b 7e 7c 74 74 62 69 5f 5e 60 62 69 68 65 66 65 5a 6a 62 5e 6b 68 64 65 6b 70 63 6d 64 60 65 64 69 64 5f 60 62 63 62 70 66 68 61 66 68 65 64 60 63 5c 68 69 6c 7d 78 7b 80 86 7f 81 72 6e 6c 72 6f 74 78 72 77 7e 6b 72 77 6b 79 7e 85 82 85 78 77 7b 7f 77 85 77 80 5e 25 08 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 0c 0b 14 26 56 87 96 96 8c 8e 87 87 86 7e 89 88 88 83 84 86 86 85 7e 85 82 84 89 81 80 7b 7d 81 7c 7b 86 78 85 80 7e 81 81 80 80 79 81 7c 7d 73 77 7e 78 77 7e 77 82 81 6f 69 67 63 64 65 5c 5d 63 5e 5f 62 60 59 58 59 5f 59 5e 54 56 57 5f 5d 5b 5d 55 54 56 5a 5b 5a 63 52 62 59 57 61 59 5e 5c 55 5c 5b 61 5c 61 60 58 59 58 5b 5c 5d 64 63 61 61 63 5a 69 80 78 72 68 5d 42 2d 2a 12 0d 05 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0f 2d 32 49 5d 64 7f 8c a6 a9 94 7d 7d 78 7a 83 84 84 83 77 62 62 60 5d 6a 6a 67 65 61 64 64 62 64 68 5b 5e 61 6a 65 6c 63 62 62 63 65 60 5e 63 67 62 67 5e 5f 66 62 66 65 63 6a 66 65 63 60 6a 5b 63 67 68 78 77 72 82 83 7a 7a 7a 74 6a 6f 71 70 6d 6a 73 76 7d 78 76 79 77 7c 81 87 7d 7c 7a 7e 7a 75 85 7a 73 66 32 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 03 09 13 1b 5e 81 8f 98 8c 89 86 81 84 85 85 81 89 80 84 7e 83 87 82 85 7b 85 80 86 86 87 84 77 7c 79 7c 7d 76 79 7b 7f 81 7e 7a 7d 77 76 77 84 7b 7f 7b 7a 75 79 70 78 6d 62 6e 56 64 5f 5d 61 5d 5b 5d 58 52 5d 5c 5a 5e 60 58 55 5b 61 5c 56 59 5a 51 4f 5c 55 54 57 5f 59 57 55 5b 60 52 5b 5a 57 5b 59 5c 59 5b 5f 56 5a 58 51 5f 5e 6b 5f 61 5b 61 5a 67 7c 80 75 67 59 45 30 24 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 06 06 18 1b 2b 45 5a 62 79 93 a5 a0 8a 7b 6e 6d 7b 78 80 7b 80 70 64 68 61 62 67 61 68 5f 62 63 5c 63 60 62 64 60 5f 66 63 64 61
 65 5f 5b 5c 5a 5f 60 64 5d 63 5b 69 62 5f 62 65 5e 5f 65 63 63 5f 65 64 6a 66 61 70 76 7b 7e 81 78 6e 67 76 72 6c 6a 6f 78 61 79 6e 69 74 6f 7c 75 76 7d 76 6c 71 70 71 7a 74 7c 7b 75 64 22 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 09 19 4d 7b 8b 92 85 89 86 7f 7f 7d 80 81 7c 78 79 7b 83 81 84 80 82 80 80 7e 88 7f 81 80 83 76 7d 7d 7d 72 74 7c 7e 7c 7c 7b 80 83 7f 78 71 7a 78 75 79 76 76 6d 62 64 61 5c 5f 63 5f 59 5d 5c 57 52 5b 59 55 5b 55 54 5f 4f 4f 5a 5a 5e 55 4a 54 4f 56 51 58 54 5e 54 62 4c 59 58 56 59 5f 57 5e 56 5a 5b 5a 55 50 59 5f 51 58 58 62 61 60 59 5d 5f 6a 74 7a 77 69 59 49 35 27 07 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0e 19 1e 2f 44 5b 6a 86 92 a4 a4 91 71 73 6e 7f 79 86 80 7c 75 6c 5e 64 65 67 68 61 5f 5c 60 60 60 66 61 5f 5c 5f 61 63 63 64 5d 64 54 61 62 5a 66 63 64 5f 60 65 62 61 6b 64 5c 63 61 60 5e 5d 5e 63 60 61 6d 70 75 77 73 77 78 75 77 74 6e 6c 6c 67 71 70 6e 6f 6b 76 7b 7b 7d 7c 71 7b 73 67 70 75 6f 73 78 79 6d 67 2e 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 09 1c 41 7f 8d 8a 8a 83 84 7e 7c 81 80 84 81 7e 7e 80 84 81 75 75 7b 7d 84 81 7c 7f 7d 7b 76 76 7a 7c 7f 7c 81 75 7e 79 84 7c 79 76 7c 7b 77 77 6e 74 80 78 72 70 66 66 64 56 59 59 5e 60 5e 55 59 5b 5b 59 5d 57 56 57 58 5e 58 61 5a 59 57 5a 5e 58 52 59 59 53 55 63 5b 50 56 58 5d 5e 5a 5f 5f 54 55 5a 52 55 51 5b 56 5f 5d 61 5b 60 5e 61 60 59 61 6f 76 7a 68 57 4a 35 28 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0d 1a 15 2c 45 56 67 82 8d a4 9e 8c 78 70 72 78 7d 7a 81 71 6d 65 5d 62 60 63 63 63 65 63 5b 61 62 62 65 62 5e 5e 61 58 5e 5b 5f 5f 64 58 57 5e 5f 59 5a 65 62 63 64 69 62 5f 62 62 65 61 61 5f 62 5f 5c 61 65 67 6a 72 7a 75 7b 72 75 70 6e 6d 70 71 71 6f 70 6e 6c 71 70 72 7a 75 75 6b 69 6d 70 73 70 72 78 75 6e 6e 33 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 06 0e 05 13 42 6f 8e 8e 8f 82 86 7c 78 82 78 7b 84 76 7a 75 78 7b 81 7b 7f 7d 7f 76 76 80 7e 75 7e 7a 7e 77 7b 7b 7c 75 7d 78 7f 80 7b 74 7b 7e 7a 7a 76 74 70 75 6e 6c 61 65 59 65 5e 59 60 5b 5b 5a 53 5a 5d 5d 58 56 55 55 57 57 60 61 53 51 5a 59 64 57 5b 51 54 51 5f 5e 64 5f 52 57 54 58 5a 58 63 5b 5f 5d 59 5e 52 56 5c 5a 5a 5a 5e 5c 55 57 5b 5b 60 6f 78 71 61 5d 4b 3a 2a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 03 06 18 19 30 49 55 6e 7d 9c 9c a7 91 72 65 60 6f 7e 80 81 72 71 5e 64 59 61 5d 60 69 63 64 61 60 64 62 5d 5f 66 68 63 60 66 5d
 5d 5a 58 58 5c 55 5c 60 5d 5f 62 5e 5b 63 5e 64 68 61 5a 63 5b 5d 62 62 65 5e 60 5d 68 70 71 6e 71 6d 6c 72 6f 71 65 6e 6d 69 68 6f 68 6e 6a 73 78 75 71 6c 62 6b 65 6a 69 6a 77 74 79 65 39 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 07 0d 3a 72 82 8c 84 7e 7b 71 79 79 80 7b 76 7d 7c 78 7b 7d 78 7c 7b 7e 7d 7d 71 77 76 7c 81 7e 7f 80 74 7a 81 73 83 79 81 7c 79 7c 7e 79 77 78 7c 70 71 6b 6a 65 5e 64 5b 5c 5a 5e 5c 5a 5a 54 56 5b 57 51 5a 5a 55 60 59 57 5a 55 54 58 59 51 54 53 51 4a 54 5a 55 56 55 52 57 60 51 57 56 60 50 61 60 56 59 54 55 59 55 51 50 5b 5d 5b 54 4a 55 53 61 6c 76 74 66 62 48 3a 2c 12 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0c 17 22 2e 43 54 6c 80 97 aa a5 90 7a 67 6b 6e 75 7e 79 77 64 63 61 64 6e 60 65 65 62 66 61 5f 68 63 61 60 61 63 65 64 5b 61 63 5f 63 5d 61 5c 61 66 59 63 5f 61 65 66 58 61 66 5f 6a 63 59 5c 5b 5b 61 65 5a 6a 68 6a 72 75 75 7c 78 75 67 6b 6d 6d 6b 6b 6a 6d 68 6a 6d 75 7b 74 72 6d 66 65 65 5f 6d 6e 68 76 71 67 39 07 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 0d 0f 30 6d 84 8f 80 81 76 74 77 75 75 79 74 75 75 71 7d 7b 77 7d 81 7e 83 77 7b 81 76 7f 74 76 75 79 7d 79 80 7a 79 7a 7a 74 75 6d 70 6f 70 7f 7d 7d 7a 6f 6e 63 64 66 57 58 59 54 54 5d 57 5b 58 5a 58 55 55 57 56 5c 52 51 57 58 54 5d 58 58 58 50 53 54 57 60 5a 56 57 59 55 5d 58 5c 5f 5c 55 58 57 5a 62 57 5c 5b 5f 54 59 59 57 57 55 54 55 4f 60 6d 72 7c 77 66 53 40 2b 12 0e 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 03 0e 0e 22 2a 48 59 71 86 8f 9c a8 92 7b 71 71 74 7b 83 87 75 6a 5b 6a 5d 69 5b 5f 66 6a 5f 5e 62 5d 63 63 62 61 5c 5b 5f 59 61 5d 61 5f 5c 5f 59 5d 59 68 60 57 60 5f 62 5b 66 64 64 62 65 5f 64 5e 5d 53 5c 65 67 6b 68 6d 75 6d 6f 77 73 76 7a 71 71 75 68 6f 69 6b 69 6f 78 6f 72 67 68 6a 6d 69 68 73 74 80 74 6f 6f 3c 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 05 12 26 65 88 8c 87 7e 79 76 6c 75 75 75 7d 72 7b 72 7e 7f 7c 75 7a 7e 75 75 75 7c 7b 71 7a 7b 7e 75 7f 7a 7f 79 7c 78 7c 72 75 7b 74 73 79 79 6e 75 6f 6b 67 64 62 5a 68 62 5b 5e 5f 59 5a 61 53 58 5d 5b 5e 5c 5f 57 53 50 58 5d 57 57 59 57 4d 52 53 57 50 51 5f 5b 64 5b 62 5b 5d 5e 5c 59 5b 58 5a 5c 5d 5a 58 53 5d 61 5c 5d 57 5c 51 5a 52 58 59 6a 77 70 70 5e 52 40 2b 19 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 14 1e 33 3b 5f 6a 79 96 a2 a3 96 87 7a 76 7a 81 84 86 72 6e 57 52 5a 5d 61 62 57 62 60 5e 5c 5c 63 62 5f 61 67 55 54 56 5d
 57 61 59 5b 5e 60 5b 63 60 5f 56 65 5d 54 64 63 61 62 60 63 63 56 60 5b 5f 55 5a 5e 5d 63 6c 69 6d 6d 6d 77 6f 76 75 71 77 60 64 66 6d 70 6c 74 74 6b 6d 65 65 6a 68 66 6f 67 6f 70 6a 69 44 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 06 05 0c 25 61 82 8a 85 73 73 68 74 6c 70 73 70 77 74 6c 72 76 75 7d 7b 6f 7a 79 71 74 6e 79 76 76 7d 7d 74 77 7b 71 7e 75 79 75 73 76 76 73 7b 71 72 6e 6d 60 64 58 63 61 5b 5b 5a 61 64 5a 5e 56 56 4b 56 55 53 53 51 52 60 52 54 5f 51 57 55 56 54 58 51 5e 54 55 5e 5a 55 5b 56 56 5a 60 5a 5e 54 5b 5b 57 5a 57 50 5f 57 5e 5a 59 55 55 51 55 50 51 5b 67 74 80 68 70 51 3a 2f 14 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 17 1d 2f 40 52 71 78 93 a2 9f 91 85 82 89 7f 90 8f 92 7e 70 65 60 5f 5b 62 67 60 59 5f 6b 60 5f 65 5b 62 61 63 63 5f 63 5f 5d 58 5a 5d 51 5b 56 5c 61 5f 5e 60 5e 64 52 60 62 55 61 5c 5b 62 56 5f 5a 61 5d 62 5c 62 63 62 62 69 69 72 6e 6f 76 74 68 6a 70 66 64 68 65 6c 73 6b 6c 6a 66 61 64 64 6b 71 76 70 6a 68 3e 17 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 06 22 62 87 8a 7e 73 70 70 6a 71 6e 76 6f 6b 7a 6f 79 7a 73 7a 75 76 77 71 72 76 75 79 75 71 75 72 7b 6f 75 79 7c 72 7e 71 76 72 72 6c 77 70 72 6d 6d 64 64 63 59 5d 56 52 53 5b 55 5b 5b 57 52 59 5a 56 59 52 50 57 51 52 57 57 57 5c 58 54 4c 54 4d 50 5e 53 58 5a 54 61 5a 55 55 57 59 56 56 51 53 5d 57 5c 4f 58 5e 5b 5b 5c 58 50 4d 49 4e 5b 5b 6b 7a 72 73 64 54 3a 28 17 09 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 09 0b 14 1f 2b 41 59 6e 7b 93 a0 99 9a 8a 8b 8c 91 92 9b 9d 9b 83 75 66 62 5e 5c 5b 67 67 5c 62 58 5c 63 62 62 64 66 5b 5e 5c 5e 60 65 62 5b 5a 58 63 60 5c 69 64 60 5d 5f 5c 58 5c 61 5e 64 5c 60 65 5e 66 55 5a 60 65 5c 5e 61 5e 68 63 70 6d 70 6b 6f 65 6d 66 6d 6c 65 6e 70 68 75 72 64 61 63 66 65 66 6b 75 76 6d 6d 4a 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 0c 1c 56 7c 92 83 7b 7a 77 76 64 6e 76 6f 6a 74 6d 77 7b 7f 70 7a 7a 78 72 79 7f 77 78 7e 77 75 7c 78 75 7b 76 70 81 7e 74 76 7b 7b 71 75 74 6e 67 62 5f 5f 5f 60 60 67 5e 56 62 59 5e 5b 57 52 4c 55 55 54 5a 52 52 57 51 56 5b 5a 5c 5a 59 57 5a 5a 63 61 54 58 4f 60 5e 5c 61 64 53 5b 5c 59 61 51 59 57 52 55 54 5a 5d 5a 65 58 56 5c 51 53 58 5f 6b 7e 74 6f 5f 4b 3b 24 16 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 19 1d 2a 47 53 66 83 91 95 96 87 8a 89 8d 96 93 98 a3 9f 8d 88 6d 64 5c 5d 61 60 5f 61 5e 5d 5e 57 59 5b 5e 68 58 58 56 5d
 64 67 5d 5a 60 58 5c 61 5c 5f 55 62 62 5a 5e 5e 55 62 5a 64 57 5f 5c 58 5a 53 5c 62 54 55 57 5e 58 5b 57 5a 65 67 5b 68 62 67 67 66 6b 6b 69 5e 74 6b 6d 71 65 64 65 68 6a 6d 60 64 66 63 4a 19 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 08 20 56 87 8d 8d 81 75 68 73 65 73 6a 7b 73 74 75 7b 76 6d 77 70 74 77 73 6d 74 69 75 76 79 79 76 72 70 79 6f 7a 77 7a 7a 74 75 75 72 6a 6f 68 6d 69 5f 5b 5e 58 62 5d 58 5a 5b 5c 57 54 51 4f 53 4d 55 54 55 52 54 56 54 4f 4d 53 5e 5b 5e 53 57 51 54 5b 5b 5a 5a 5b 56 57 61 51 57 5a 5d 5b 5d 53 56 59 5e 54 59 59 5b 59 5b 59 56 4f 56 4b 54 5f 60 7c 75 71 66 4e 3a 28 0f 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 11 10 28 3c 51 67 77 8b 96 9a 89 7f 86 86 94 96 9b 9f 92 96 88 7b 6d 5d 64 61 60 61 6b 5e 5f 5f 5b 54 5e 55 5f 5e 60 67 5d 58 60 55 5e 5e 5f 5d 5c 61 62 5c 59 59 58 5d 5e 5e 5a 5f 5d 5b 52 57 53 5a 52 59 59 59 56 56 53 5a 5d 5a 64 62 5d 5b 67 63 68 69 59 64 69 68 74 70 67 67 6d 65 66 61 65 62 6e 6d 67 66 67 54 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 06 16 55 82 96 90 91 84 74 6b 6e 67 73 74 6a 70 6e 6c 73 75 70 6e 70 6f 76 6f 73 73 75 75 78 76 7a 71 74 74 71 71 80 75 77 77 77 76 70 6c 74 6b 63 5f 61 5e 5e 59 63 56 57 58 5f 58 5a 52 55 5b 56 58 55 54 52 50 59 4e 50 55 5d 4e 51 53 5a 53 53 5c 55 54 58 56 57 5e 59 5e 58 57 5d 4f 57 54 58 56 56 57 50 5a 53 56 52 5a 5a 5c 57 52 55 4c 4a 5e 6f 76 73 70 5d 4f 38 2a 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 11 21 3f 58 6c 7b 8f 92 96 84 70 7c 80 8d 8c 9c 98 a0 8c 8a 81 71 66 5b 5c 62 62 5f 5c 5e 61 5e 68 60 5b 5f 55 5f 68 59 60 63 61 5d 57 57 55 5a 53 63 59 5b 63 5b 61 56 57 5f 65 60 5a 59 55 5b 56 57 62 5b 5f 5d 4d 59 59 53 5a 5e 57 5f 64 62 66 5c 5f 62 69 66 73 77 78 76 72 62 64 69 6d 62 6b 6e 69 6f 6e 6c 51 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 16 50 7e 87 92 88 85 7e 70 6f 6f 73 6e 73 6b 68 70 72 74 74 77 6b 6a 70 77 77 76 79 78 71 7b 6f 72 6e 7a 79 75 70 76 76 6f 7c 6a 6b 69 64 5e 5e 61 60 55 59 59 5e 57 57 5f 54 61 5b 5e 56 53 4e 54 55 58 5d 52 52 51 4f 51 57 53 56 5f 5d 5f 52 59 57 54 5c 64 5a 60 55 5b 54 5c 59 5c 59 54 57 50 5c 5a 58 51 5e 5d 4d 59 5a 56 5e 51 51 51 57 64 72 76 7a 68 5d 4e 34 26 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 11 29 36 4f 66 76 91 93 92 86 72 71 77 85 84 93 92 96 90 80 80 85 6e 6a 63 66 69 64 61 61 62 61 62 58 57 56 57 5c 5e 5f
 5c 61 5e 59 60 5e 5e 5a 61 55 5b 57 5f 62 58 57 63 5a 5b 58 5d 5d 55 5d 5e 57 52 52 5b 53 51 5a 5d 5c 54 5b 4c 5d 61 5e 64 5a 61 63 70 6a 74 7d 83 80 6f 70 63 60 66 5c 6a 69 63 63 63 6f 53 1c 05 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 08 03 0f 48 6d 80 8b 86 84 86 7c 72 73 6c 75 74 71 66 75 78 65 78 6f 7b 72 6f 70 6b 73 6d 68 70 6c 6c 6c 6e 74 6c 73 70 7a 76 72 6d 63 63 65 61 63 5d 5c 5b 5b 5b 5d 57 58 54 51 5a 5c 55 57 51 53 58 54 59 54 56 51 50 5a 50 59 57 5e 54 5a 58 4e 4e 52 56 51 55 5e 57 58 52 59 55 56 57 57 55 52 50 5c 55 59 53 57 58 5a 4f 54 5e 59 56 50 55 47 52 66 6a 7c 75 63 59 44 2e 20 0e 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 13 1f 32 51 5e 72 88 91 8a 85 6e 6d 67 71 82 89 8c 92 8e 82 84 8b 85 74 67 67 67 6a 5f 66 5e 57 5e 56 5a 5f 5f 62 60 53 5a 5f 59 52 5c 5b 58 54 56 5b 5f 52 56 55 52 5d 5a 5a 58 57 5b 57 62 4e 59 54 57 55 57 56 54 5e 5a 56 5d 52 5e 5f 60 5c 64 5c 65 65 60 6d 7e 85 83 7f 68 5a 60 5e 61 63 62 69 64 65 5a 64 57 27 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 39 71 84 85 85 84 8c 7c 79 75 74 6f 72 6e 6e 76 6c 70 69 73 6c 71 6e 72 72 6c 73 78 72 76 70 78 70 74 6d 6d 72 70 68 6c 6e 6e 67 64 5f 5b 53 5f 57 62 57 56 5c 5c 57 54 59 5a 53 4e 4d 4f 54 55 52 5a 52 54 4e 54 52 5b 4f 4e 54 55 51 56 52 59 5e 5d 60 58 59 55 59 5b 5e 55 57 59 53 56 57 50 59 50 51 4f 56 59 59 54 5f 4d 50 4f 50 58 59 6b 6b 79 73 5f 58 39 28 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 14 33 45 62 6f 7f 93 93 85 6d 69 6f 6b 6d 79 82 84 7e 79 76 83 92 88 75 70 69 64 5a 54 5e 5a 5b 5b 55 57 5d 60 5c 5c 60 5e 5c 5c 5b 5f 56 61 57 5a 55 55 59 59 53 51 5d 59 5e 55 57 5e 57 60 57 58 58 4f 4f 5b 4f 56 56 4e 4e 5d 59 5f 61 52 5e 62 65 66 64 74 70 7e 7b 6c 6c 6b 5f 5f 67 5f 63 5f 6a 67 5c 60 4f 20 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0b 2e 70 81 79 81 7f 85 7f 7d 7c 80 79 7f 7a 79 75 73 75 6b 75 70 71 72 69 6d 71 6f 74 6b 68 73 6d 6c 75 6c 70 68 78 67 71 6d 68 67 62 60 5f 55 58 56 5e 5a 5d 5a 55 53 5a 5c 57 52 57 53 5b 59 56 53 52 51 4f 4f 56 4f 5a 52 55 55 5a 53 53 58 55 59 52 5d 5d 53 5e 58 5b 59 59 5d 53 57 58 4e 5e 4f 58 59 53 57 57 4b 57 5b 59 54 50 54 4d 59 6c 77 75 71 63 50 3f 2c 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 10 10 2a 3f 57 75 84 87 88 83 74 71 6b 69 76 70 7a 86 79 77 79 7b 88 94 89 73 6b 5e 61 57 5d 62 60 5b 5f 5b 5a 59 59 5c
 5a 5f 60 5c 5b 5a 5d 5d 54 58 57 5c 5c 5a 55 4f 5e 56 53 5a 54 56 4d 53 52 55 54 5c 50 50 4f 50 53 51 4d 54 54 53 52 55 62 5a 60 69 67 5f 70 72 70 6e 67 6a 5f 64 6c 64 5c 66 66 65 5f 61 53 27 06 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 30 6a 7b 81 7f 7d 7b 85 89 80 80 81 7e 7a 73 79 7d 7d 79 79 71 73 71 6a 74 6f 72 72 73 72 6d 6a 70 74 63 6b 77 69 6b 61 5d 64 58 5b 60 56 62 61 60 60 5f 5d 5f 5e 56 50 5e 58 51 56 4e 5a 59 55 4a 5a 56 50 56 50 50 50 51 52 54 58 52 55 56 5e 56 59 5a 5e 59 54 62 55 51 52 5b 5c 58 5a 4e 53 55 55 5e 5c 55 59 52 5c 53 50 56 54 5b 57 5c 60 6b 6b 69 53 4b 33 1a 15 07 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 06 0f 14 1e 37 49 66 80 88 90 8e 7c 6e 65 6b 66 6d 6c 74 6f 79 6d 79 8b 91 92 80 6b 61 5d 52 5c 5c 58 4c 4f 5b 5e 58 59 63 5d 60 59 56 58 5e 55 50 58 57 59 4d 5a 53 64 58 52 51 61 54 5a 58 56 5a 5d 5b 4f 58 4c 50 51 4d 4c 4f 51 54 57 59 5d 56 5e 5c 63 5f 5e 66 6d 66 66 6e 6f 61 64 66 6a 67 5f 60 62 65 5a 60 53 29 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0b 29 5f 79 7c 80 7c 7d 84 7b 81 76 83 71 72 74 78 80 80 81 80 7a 7c 80 73 7b 77 6b 74 73 71 6f 6f 6d 71 71 66 6c 61 65 5f 62 62 5d 5f 5f 53 58 5a 58 5b 57 5c 57 58 5b 59 54 55 50 4f 54 57 57 4d 4a 52 52 55 55 4f 50 53 4e 55 55 56 4f 50 53 5b 57 56 51 58 5b 5b 5a 53 4f 53 59 50 53 54 4f 59 5a 53 52 53 4e 55 4a 52 54 54 5b 51 5c 50 52 5f 6a 6f 62 4d 33 2b 1e 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0a 0d 0e 1a 2c 4c 68 7b 7e 98 8e 7e 75 69 67 67 6c 69 6b 72 71 70 6d 79 82 89 87 79 6e 58 55 55 59 5b 58 5e 61 52 5c 59 5e 69 5d 5a 5a 59 5d 5a 56 5c 5d 54 5b 4b 61 56 57 5a 54 52 5c 52 50 5c 53 55 55 5b 55 52 54 4f 4f 50 52 54 53 4f 50 56 5c 61 5f 5d 5c 5c 61 65 5c 69 60 6a 67 66 5e 61 59 57 64 64 60 5f 62 5a 2b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 27 5b 81 7e 88 80 7a 86 84 81 81 79 7b 74 75 7a 76 76 80 7b 7c 7a 80 7c 7f 76 7e 71 6a 72 73 6f 70 6e 6b 6f 6b 6e 6e 61 61 5a 5a 56 54 55 5c 58 5a 5e 62 60 64 58 60 62 5a 55 53 50 4d 57 55 4a 55 52 52 4d 50 54 4d 50 51 54 56 57 5e 55 56 57 52 4e 55 68 55 59 55 60 5a 54 57 55 5a 51 51 50 58 53 60 53 4d 5b 54 59 5c 5e 5e 59 57 5c 53 5f 68 5f 50 43 33 26 19 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 12 2c 48 5e 79 83 8a 8f 7d 79 6b 6a 64 64 6c 6c 6e 6f 65 6b 72 86 81 94 87 71 5c 51 59 57 55 55 58 58 5c 56 50 5f
 5f 50 56 54 55 5a 4f 51 59 55 5a 5d 55 52 56 4f 56 56 52 5e 55 53 5a 4b 57 52 4e 54 50 59 5a 53 55 52 57 56 52 59 59 5c 5b 5a 58 5b 5e 57 60 5e 62 67 6b 64 68 68 5a 62 5b 66 65 66 5a 60 54 2f 0c 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 23 58 84 85 87 7c 87 81 80 7c 79 85 70 75 64 6b 72 70 73 73 79 76 74 79 7c 78 76 79 79 6f 70 6b 6b 72 68 61 5f 5f 62 5d 61 5d 55 59 5e 5a 5d 54 5a 58 5f 58 5b 5a 4f 5d 55 5e 51 52 56 50 58 4e 56 56 51 4f 4d 4d 4e 53 50 51 55 5b 55 5c 57 58 4d 50 5c 5e 61 5e 5a 5e 52 53 51 4f 52 5d 55 53 5a 56 54 51 4b 5c 59 59 52 5d 5c 55 56 56 55 56 59 53 4a 36 2c 1d 14 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0b 17 24 38 54 6e 81 88 85 7c 74 69 65 69 65 66 6d 70 72 73 6f 70 76 7c 95 8f 72 5c 4e 4b 5c 4d 50 56 53 53 54 5b 5c 56 5c 55 54 4e 50 50 55 4f 50 48 59 53 4e 4e 55 4e 54 52 56 4d 53 59 5f 5a 57 55 50 4d 49 54 51 50 56 4d 4a 54 4f 4d 51 56 54 57 58 55 61 62 5e 60 5f 66 6b 6a 60 62 5a 5b 5e 63 68 61 65 55 35 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 15 61 7d 86 96 8c 83 87 7d 77 77 74 78 77 73 6f 79 6c 75 74 72 70 6f 73 74 72 7c 72 76 6d 68 70 67 6c 67 5e 5d 64 57 60 58 53 5b 56 59 56 54 5a 5b 5a 5a 50 4e 5e 52 54 4f 56 53 4e 5b 59 4e 56 51 50 4d 50 4b 48 51 52 54 54 56 4c 4b 57 51 55 57 55 55 57 4e 58 54 5d 5b 57 5b 56 59 5e 55 5b 58 51 51 50 56 5e 5b 52 52 59 58 59 55 55 59 50 4b 41 3c 2e 1e 17 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 06 06 09 09 0c 12 24 32 52 65 72 8d 84 7b 71 67 64 66 6b 68 67 63 6c 6e 6c 71 74 82 8e 9c 76 62 5b 53 4e 50 5b 59 59 5f 4e 5d 5d 5b 59 57 53 53 55 52 53 55 50 59 4d 4d 4f 56 51 4c 52 56 57 52 56 59 58 53 50 50 4d 53 52 56 54 57 56 4c 50 4f 54 58 55 5e 52 57 57 53 5b 5c 5d 55 5c 63 6a 62 6f 61 5a 62 5e 5e 59 69 5e 60 3a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 19 5d 88 8a 94 8b 87 77 84 7c 7a 72 74 74 66 73 75 73 66 6b 70 73 6e 6f 76 71 79 80 7b 77 69 74 69 66 64 61 59 5e 5f 5d 5a 52 56 5a 5f 5b 4a 60 5b 57 5a 54 50 60 56 51 56 56 4e 50 59 50 4e 55 4b 53 54 51 4f 4d 55 4f 52 51 4f 53 4e 47 5a 5d 55 55 57 5d 5a 58 59 56 57 55 5d 52 5d 53 5b 55 5c 55 57 56 5b 5e 59 53 5b 59 5b 5c 55 56 44 51 4b 3f 3d 21 1b 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 03 0d 0d 1b 21 3a 58 75 7d 91 80 6a 6b 65 60 5c 62 60 67 69 66 68 66 64 7f 89 90 7c 58 51 54 52 5b 56 59 59 52 5c 5f 60
 61 5a 57 58 5e 56 52 59 55 58 50 4d 54 58 54 61 54 55 52 55 5a 56 52 54 58 56 4d 4f 51 53 56 4e 50 4e 49 59 4c 58 4d 54 58 57 59 57 58 5a 5c 58 62 5f 60 64 6a 66 5b 5c 60 5f 66 65 56 65 5b 3f 14 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 06 19 55 84 8a 91 84 7e 83 7d 7c 76 7a 74 75 68 6f 70 6f 72 6f 6b 71 77 6c 73 7a 7b 7d 79 7b 7a 7a 62 72 5d 66 5e 63 5d 5f 5d 5f 5c 50 59 5d 57 57 56 55 55 58 56 55 58 59 5e 51 5b 57 52 57 52 56 46 4b 5c 50 51 49 53 54 51 4a 52 50 56 54 4e 54 59 4d 59 61 51 5a 5b 57 5b 4f 59 5a 5f 55 59 55 5d 5b 56 56 60 57 59 5e 5c 60 5d 5e 59 54 50 4d 45 36 36 23 11 0d 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 03 04 10 0c 22 30 4d 67 7e 86 79 6a 63 5f 57 58 61 61 61 62 69 67 62 5d 66 74 7d 72 5c 52 55 57 53 53 58 4a 52 50 52 57 58 5e 55 58 52 4e 4d 59 5a 49 57 50 4e 59 52 54 56 52 5b 57 4b 5c 56 55 4c 50 53 4a 4b 4c 4e 49 52 50 54 54 4d 55 54 4f 5a 54 57 5f 60 59 5a 5a 5d 57 64 5f 62 65 66 5f 61 5b 61 5f 66 5a 5e 46 15 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 09 11 49 76 87 8b 84 83 78 75 78 75 6f 73 77 69 72 6f 71 69 70 72 75 6b 6a 6e 6c 78 7d 7a 82 72 78 6d 6e 67 60 5e 58 5a 57 5b 5b 4e 57 52 54 58 57 54 57 62 54 57 5b 52 55 57 4f 4d 52 5a 5b 53 4d 4b 4a 50 50 4b 52 4b 50 4d 4d 52 4f 58 54 4e 50 55 58 59 4e 5a 54 4d 5b 5a 53 5c 59 5b 56 57 59 5a 4e 62 56 5d 5e 59 60 5a 61 5b 5b 65 4e 54 44 39 38 2f 1d 17 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 09 00 06 10 11 28 46 63 79 7f 87 71 62 58 5a 5a 63 68 63 68 60 67 5f 5e 65 74 6a 65 5b 57 59 54 50 53 55 54 52 54 56 5b 56 5d 57 4e 52 53 59 54 4c 55 43 51 50 50 5a 56 55 54 57 53 4c 51 56 51 4f 51 51 4e 49 4d 52 57 5b 57 51 52 4f 4f 59 56 53 58 59 5b 5e 5b 50 5d 5f 53 5f 5f 64 5d 59 5e 60 61 62 67 61 68 53 45 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0f 45 76 89 89 86 75 7f 79 75 73 70 70 69 67 75 75 6c 69 62 70 6b 68 6e 63 68 6a 70 75 75 70 6e 6c 73 5f 61 5a 62 56 58 54 64 5b 58 5c 4c 57 5a 58 5d 5d 5b 55 59 5b 57 58 56 4e 52 4d 54 4f 52 55 4f 50 4a 4e 53 4b 53 4d 4d 53 4a 53 4a 51 51 5e 54 54 55 59 50 5d 5e 58 59 4d 56 52 56 59 57 59 57 5a 56 63 5e 5b 56 5a 5a 65 5f 61 55 4a 4a 39 3d 20 16 16 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 06 05 06 06 15 0f 12 20 34 4c 6e 7f 8b 76 6c 62 5b 5c 65 68 66 6f 73 6b 67 6b 63 5f 62 5b 58 52 58 50 53 56 56 50 56 54 5a 59
 5d 52 55 51 5d 50 49 54 4d 52 56 54 50 58 50 48 55 53 55 54 57 53 56 4c 56 55 5a 4d 4f 53 4d 58 4e 50 51 52 4d 55 55 51 54 52 5a 5b 5d 5c 5e 5c 5b 5c 5f 5b 69 5f 62 62 5e 60 64 5d 5b 60 5d 48 0f 01 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 10 44 7b 85 8e 89 77 7f 77 6b 78 7c 6e 6b 6b 6e 6d 66 6c 6a 72 70 6f 6d 70 6e 70 6d 6a 70 6d 69 6a 66 63 65 62 5a 60 5e 59 5c 5e 53 4f 5c 56 5c 5a 54 56 56 55 59 5b 5d 5d 54 4e 52 56 56 55 5b 4f 51 5b 58 55 48 49 4e 4f 4d 50 4e 53 50 54 64 54 4f 51 58 58 5e 4f 5f 55 50 5c 51 5d 52 59 4f 5a 58 56 5c 5e 64 5e 5d 5b 62 65 59 5a 4c 48 42 39 35 22 14 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0c 06 10 11 1e 2a 3f 5f 74 85 79 66 6e 65 5d 69 6a 71 75 71 75 65 61 62 63 59 54 52 52 56 55 52 54 51 54 4b 50 51 5d 53 53 55 4f 53 53 4d 58 50 53 57 53 4f 43 56 4e 4c 4e 4f 54 54 4c 52 52 4f 55 4e 4e 47 52 5e 56 59 55 4c 4c 60 57 5b 50 54 5b 61 61 5c 56 5d 5c 5f 5d 5b 63 62 5d 62 61 5c 5c 5f 57 5a 5c 5e 4c 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 01 0d 36 72 85 8b 84 7a 7f 77 7a 73 79 70 6d 6d 72 73 68 72 6a 6b 74 6c 6d 6d 64 61 6d 69 6a 5d 70 60 69 5c 5f 5b 59 51 5a 5d 57 59 5b 56 53 4f 5c 4e 4e 5e 50 53 5b 55 58 56 59 5d 50 55 4e 55 57 58 51 4f 55 52 51 4a 4b 4c 4e 50 55 51 4f 54 4a 57 4f 52 5c 58 54 57 58 5e 53 53 5a 58 5b 57 59 62 56 55 5e 5f 66 5e 5d 5b 57 5d 5f 5b 4f 51 42 42 26 21 0e 11 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 08 05 0c 14 19 29 40 62 74 81 6e 64 6d 5c 68 65 6e 76 77 72 64 63 60 4f 54 50 50 57 4e 54 51 4e 52 54 52 56 56 59 52 59 52 4a 52 4c 4d 50 4c 55 4e 4c 50 4b 4f 4f 51 55 53 56 48 56 4c 4e 55 52 50 50 4a 56 4f 55 52 49 58 57 54 52 59 4e 50 52 57 5c 63 53 58 55 59 54 56 5a 5c 5f 5b 62 5c 51 5b 5a 59 5d 55 45 17 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 30 72 81 8d 83 7b 7d 72 73 75 74 6a 6d 72 72 6d 6c 68 74 6c 6e 68 6b 69 65 67 6a 6b 65 69 67 63 5f 60 5d 56 59 50 60 55 56 56 52 52 52 55 4b 4e 54 56 59 4f 54 51 59 55 50 5d 4c 56 5b 4d 54 4f 54 4f 50 4c 4a 4e 52 4b 4c 4c 54 4f 55 4d 4d 4d 53 56 58 58 5c 4d 52 4d 50 57 53 5c 53 57 5a 5c 5a 5e 5b 5e 5e 60 5f 5c 57 5b 56 4f 46 41 3e 2f 25 1f 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 07 10 0b 14 1d 25 43 60 75 7d 6c 5c 56 52 56 58 65 65 61 60 67 5f 4e 54 51 48 4e 50 50 58 4c 4e 50 50 45 4d 4c 4c
 47 4e 4c 53 4f 4d 49 49 4a 4a 45 4a 4c 44 45 46 4d 4f 47 4a 46 49 50 43 51 46 49 47 3f 45 45 4c 4c 42 47 4b 4b 50 49 49 50 4e 4b 55 53 4b 4f 52 56 54 5a 56 57 53 5c 53 52 53 58 55 55 50 4f 3b 1e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 20 5d 6a 76 6e 73 6f 72 6c 6e 63 66 64 64 64 63 55 64 5e 67 66 5c 60 64 5f 63 63 5d 66 62 5f 66 63 65 63 62 64 58 59 56 57 52 55 52 51 4a 42 51 45 4d 52 4e 4b 4b 53 4f 53 4b 4f 4d 46 4c 50 46 4d 47 46 4b 49 4e 47 47 4d 47 4b 49 4a 4b 52 46 52 56 50 59 53 4e 55 56 59 57 50 5b 54 50 5a 52 56 59 4f 54 52 4b 51 52 53 59 4c 50 55 4b 4e 39 2a 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0e 10 0b 18 21 3d 57 71 73 65 5e 57 53 5c 60 65 63 5e 64 57 4c 4f 4d 50 51 4c 49 4b 4c 4b 50 4d 53 4b 51 4f 4d 4d 50 42 4b 49 4b 46 47 46 43 41 3f 43 4d 46 4b 47 46 47 46 49 48 48 47 49 4a 52 4a 3e 3c 47 49 42 48 4b 48 4d 49 52 4b 52 52 4f 51 4d 54 54 53 57 51 55 57 56 5b 55 50 4e 56 57 54 4c 58 50 47 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 56 72 74 78 73 6e 6e 64 6d 66 69 6a 63 68 67 64 64 60 5d 5a 5b 64 58 5b 65 63 61 5f 5b 65 5e 66 67 61 67 5d 57 58 56 4f 50 4e 4c 50 4f 50 49 4a 50 50 4b 4b 50 4e 50 53 4a 50 44 46 47 4d 45 52 43 49 4a 45 47 48 4e 50 4c 49 49 4f 4e 4b 53 57 51 53 57 5b 54 51 54 52 5d 58 53 54 4f 50 57 53 54 50 4f 4b 50 56 53 4e 54 5a 54 48 50 42 39 29 0f 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0b 05 03 10 0f 1b 2b 3f 69 6d 66 56 4f 52 5d 63 6d 76 63 5a 5b 49 46 50 4c 4d 47 4a 43 44 52 50 47 54 4a 4d 4a 4d 4d 49 41 48 49 4b 3b 49 42 56 41 42 4b 52 44 44 41 47 42 49 4a 42 46 44 49 49 51 38 47 43 4b 4d 43 44 45 54 47 47 49 4e 57 50 4d 54 52 58 4b 57 57 51 54 5b 4f 5a 52 54 56 52 51 55 53 4d 50 44 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 51 6a 73 75 67 72 6c 6d 68 67 68 65 55 69 60 5b 62 62 5f 5f 54 59 5d 5e 61 5d 62 66 62 5a 56 62 60 6d 73 6b 62 58 58 50 5e 4e 52 52 4e 4f 4c 4c 4b 4b 52 51 43 45 49 44 4e 44 51 4c 49 4f 50 4e 45 41 3d 47 44 49 4c 48 4b 4a 4b 4f 47 4a 4c 4b 53 56 55 5c 4e 54 52 54 58 51 5b 5c 50 5a 51 55 55 52 4d 54 5b 53 57 51 55 4d 4d 46 45 46 33 18 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 06 10 13 12 13 1f 2b 43 53 65 61 5e 55 56 5b 60 6c 72 6a 65 58 4e 48 4f 48 4e 51 4a 4e 4d 4c 4b 4d 51 43 43 43 4e
 49 4e 4b 4a 49 4b 46 53 45 43 4f 4c 41 46 49 4c 48 4b 42 50 48 4e 46 40 4a 47 47 4b 48 4a 4d 4e 4e 49 41 4c 43 4c 52 4c 50 4c 51 52 4d 54 50 54 52 55 58 5f 54 5f 55 4f 50 4c 57 4e 52 49 4e 40 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 49 64 71 71 6f 6e 69 6c 72 74 62 61 5f 65 63 5d 5e 5e 5d 63 59 5a 5a 5e 60 5a 56 61 5e 64 58 5c 60 63 6c 73 63 5b 56 52 52 51 4e 50 4a 4a 4c 50 4a 4c 4f 51 4c 4e 52 4a 48 41 4f 47 41 44 44 4e 4e 4a 4c 4c 47 49 4c 46 49 50 50 52 4a 4d 4e 53 4c 52 57 56 54 58 4e 55 5a 53 51 57 54 5a 4d 50 58 4f 50 58 5b 52 56 58 50 52 53 4a 49 42 2a 1a 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 09 0c 0a 14 16 17 28 37 41 60 63 5b 50 57 63 60 60 6c 68 59 4f 52 53 49 51 50 48 49 46 4f 4b 52 49 4b 47 45 4d 46 49 51 4c 49 48 41 40 4e 45 4a 45 4b 44 47 4d 45 4c 46 41 45 43 4b 49 48 4a 44 42 4f 4e 4b 4f 48 4f 4f 4d 4d 50 45 49 4c 55 51 54 55 4a 53 4e 4e 58 52 55 58 4b 59 57 58 47 50 55 4f 50 4c 48 43 19 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 44 69 6b 71 6b 6c 6d 67 6d 64 5f 63 5e 65 61 5c 59 60 57 60 5d 5f 5c 5d 64 5e 5c 61 61 5d 55 5c 5d 66 6d 6c 64 5e 56 4e 4d 4f 50 50 4c 4a 4a 49 4a 4e 4b 4d 49 47 52 4e 4d 4a 4d 45 44 49 48 45 4f 46 47 46 48 4c 43 4c 4d 49 4d 48 50 4d 52 50 51 5d 57 5c 4f 4f 57 58 52 58 59 5b 4c 5c 5e 54 54 53 54 50 4e 52 5d 5d 56 54 52 4c 43 36 2b 12 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 06 07 0f 11 14 29 2f 47 54 5f 5f 57 5f 58 55 5b 5b 5b 5d 4a 50 40 42 4e 45 56 4e 4d 45 47 45 46 4b 44 48 45 4e 42 51 43 4d 42 3f 43 43 42 46 4a 42 46 43 3c 50 46 47 4a 4d 43 4a 46 4a 49 49 41 4f 42 46 48 4d 49 49 53 4f 56 47 4b 51 4f 51 4c 49 4a 4d 53 4f 58 4f 54 51 52 59 52 4e 4e 4f 54 51 4c 45 46 45 28 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 38 61 65 6c 6e 6f 6d 65 65 6b 5a 6b 59 61 5b 57 5d 59 5d 5f 5f 56 5d 55 57 59 53 63 5e 5e 5c 57 5f 56 61 64 60 5b 56 4d 4e 4d 4d 57 51 4a 51 54 45 49 50 50 4c 4c 4e 49 49 47 50 4a 44 46 43 4a 47 4a 50 4d 46 48 56 4a 50 4e 4e 4d 42 4d 4c 4b 54 51 4a 5a 48 50 5c 58 59 55 54 5b 57 5b 59 4e 5d 4b 4f 57 53 56 59 54 55 53 52 4e 43 3c 20 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0d 15 14 14 23 36 41 54 5d 60 56 5d 5f 53 58 50 50 55 4d 56 43 4c 4b 49 50 50 46 44 52 47 43 49 44 52 4c 52
 40 47 47 48 4d 4b 3f 48 4e 48 4f 46 46 4a 4c 49 4a 45 45 47 4b 49 47 52 50 48 4a 45 4d 4d 51 46 4f 51 4c 53 47 4c 50 54 56 4c 4d 48 52 50 4f 53 59 55 56 54 53 5f 5e 52 50 57 51 4c 4b 52 51 48 24 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 3e 57 65 70 66 6e 63 6b 6b 6b 63 60 5d 61 64 62 5d 5d 63 60 62 5d 55 60 54 58 57 5a 58 5b 5a 61 56 57 56 56 61 5a 4e 54 50 4a 52 52 4e 46 4e 50 58 53 50 4f 4c 4b 55 57 4e 4a 44 4b 49 48 45 4d 49 47 4d 44 42 4f 50 45 49 52 44 52 52 56 52 54 55 5b 50 5b 53 53 5d 55 5b 5d 5a 5e 57 55 5f 56 5d 56 5a 57 50 51 56 59 51 5a 53 4d 44 30 20 10 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 02 10 1f 21 26 2e 4e 54 5f 60 5a 5b 53 50 4d 50 4d 3f 44 4b 4e 4b 4b 42 49 48 4e 45 51 48 4f 4c 4e 4c 44 4a 4b 46 48 4d 46 41 48 42 43 43 49 49 41 49 4b 49 46 4e 42 46 4c 4d 4d 4b 4c 4a 49 48 46 50 4f 55 50 4b 48 4d 50 57 51 52 4f 56 52 50 52 50 4f 56 4c 53 5c 57 59 5a 56 51 51 54 56 4b 4f 4b 40 30 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 36 5f 5c 62 60 6b 65 60 62 64 60 60 60 5f 67 58 5c 5e 55 64 5d 56 53 5f 58 59 55 57 5a 5c 55 55 56 5b 55 51 59 56 52 55 4e 51 50 58 4e 4f 48 53 52 48 4b 52 4c 43 49 4b 46 47 53 4f 4c 45 46 4c 46 46 51 47 3e 3f 4e 4c 50 48 4e 54 44 51 4e 4f 52 5d 58 5f 50 58 4d 52 5f 51 54 55 59 59 55 55 5c 52 56 55 54 53 56 53 5b 4a 56 44 40 2f 17 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 09 0b 0e 0f 17 1d 23 37 44 44 54 58 5f 57 4e 4d 4f 4c 45 51 4d 4f 46 51 4d 47 47 4e 52 48 48 50 53 45 48 47 42 47 45 47 48 42 42 4c 43 4d 4a 45 45 49 48 43 49 4b 4d 4a 47 3f 4f 51 4b 56 52 48 48 4c 4f 51 56 56 45 4c 51 52 47 4b 4c 4b 54 56 4f 52 51 48 53 57 53 53 51 58 5b 59 5c 4e 56 4a 4d 4a 4b 45 44 29 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 30 55 5a 63 61 60 66 61 66 60 5d 55 5c 5d 5d 5d 5c 56 60 53 5b 5c 57 55 57 54 56 51 5b 53 58 5e 5a 5d 54 57 55 49 55 50 46 4b 4c 48 44 4b 49 48 4b 4a 4b 49 4c 51 4d 41 4d 4f 4e 44 48 4f 41 54 4f 4c 4b 51 4b 47 4b 47 4e 49 4e 4c 47 50 53 54 50 50 52 52 59 51 5a 55 55 56 57 5c 56 55 59 58 62 5a 52 57 57 52 4e 52 50 52 4b 43 2f 26 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 09 13 10 13 21 2e 38 44 58 55 5d 5c 4c 47 4b 47 4e 4a 4a 50 49 49 40 46 47 49 4f 51 4b 4d 4d 52 48 50 4f
 44 4b 51 3d 47 43 47 49 4a 43 4c 4b 4e 49 45 49 49 4b 4b 4e 47 4a 4f 47 4f 49 4b 48 4c 4c 58 40 29 3b 58 55 4f 4c 4a 4f 53 56 53 4d 49 4d 4c 51 58 51 57 51 4d 53 58 53 5c 54 53 4f 51 53 41 40 36 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 34 56 65 66 5d 61 5d 5f 65 5e 62 5f 5c 58 60 58 58 5b 55 5b 52 58 5c 58 4b 5b 5e 53 54 5a 58 58 51 57 5d 53 51 51 4a 49 50 49 54 48 45 41 41 4d 52 46 46 51 49 4c 50 50 4e 50 4e 4a 49 49 49 53 46 4c 4d 4d 50 48 4b 47 46 47 51 4e 50 50 54 5b 51 4b 55 53 53 56 57 56 59 56 5a 5f 5f 58 5e 5c 5a 53 54 51 51 5b 52 51 52 4d 50 37 2e 23 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 07 10 11 13 1c 1d 28 3d 3c 4a 52 55 57 54 49 4d 43 49 4d 4a 4c 4f 47 4c 49 4e 4e 4c 4c 4e 49 4a 4d 49 4c 47 45 47 49 4a 4a 49 49 4a 48 4a 4f 46 53 4a 42 4c 4f 44 4f 48 50 50 4d 46 54 4a 49 54 4a 51 4e 4c 51 54 57 4f 4c 50 51 51 57 50 50 52 4d 4f 50 4b 4b 4d 4c 55 5b 5d 5b 60 58 5e 60 58 4a 50 48 44 33 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 26 49 5a 5a 57 5a 5a 5a 5b 60 59 5b 55 5e 5e 4e 5b 59 54 5a 55 5f 5b 52 55 50 50 4c 52 57 5b 54 58 5d 59 50 50 55 59 50 45 4d 50 4b 4b 4d 53 54 4e 4d 4f 47 43 51 51 4d 48 4d 42 56 45 45 4e 57 45 4d 4e 4d 51 4c 50 4d 45 4a 47 57 46 51 43 55 4f 54 5e 56 55 58 5d 51 58 58 5e 58 55 62 58 54 5a 5b 5a 4f 54 57 4b 57 58 51 51 40 2f 1d 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 03 0b 0f 17 20 24 32 38 4a 4d 4e 59 54 49 4d 4a 3f 48 46 4c 4c 4f 4c 4c 45 4e 47 4c 3f 4c 4c 47 4e 45 46 45 44 48 44 48 50 44 48 4a 45 44 43 4b 53 46 49 4e 4a 4b 45 4b 4e 48 4e 51 54 49 51 4d 49 58 50 4c 49 4b 53 46 4e 52 48 56 56 53 52 4b 53 51 54 59 54 51 4e 55 56 53 59 52 5b 61 59 56 53 3f 46 37 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2a 4a 54 59 54 5e 5e 51 60 56 58 61 53 5b 54 57 54 59 54 5b 51 58 52 52 52 54 56 53 51 5b 4d 59 58 5a 5b 53 46 4d 4a 4c 4b 48 4e 45 4b 47 47 45 4c 52 45 4a 3e 4d 51 4f 4a 4d 4d 4b 46 45 47 4f 42 49 44 4a 45 50 44 50 41 4c 4f 4a 4d 50 4d 50 50 55 59 57 50 55 55 54 56 50 59 5b 54 5c 53 57 58 50 4d 57 4c 4d 4f 50 53 43 42 33 29 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 14 1c 2f 21 2b 33 48 47 4c 52 4d 4e 47 45 42 49 44 4a 45 4a 43 40 4b 4c 51 4a 4f 4a 47 48 41 50 4b
 42 48 52 43 4c 44 4b 46 46 4d 49 48 45 4f 4f 4e 45 47 47 51 40 45 41 47 4f 53 4a 45 4f 48 4d 4e 51 4b 4d 54 4d 4b 4b 4f 4a 52 59 59 51 4f 47 52 56 5b 58 58 51 58 51 57 59 5a 65 6b 60 52 50 42 34 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1b 47 51 5d 50 54 53 55 57 5d 57 56 50 5b 59 5b 57 57 50 50 57 57 55 51 55 57 56 51 4e 50 4c 51 53 56 51 53 51 52 4d 4c 4a 4d 4d 48 44 47 4a 47 41 4e 4d 4c 47 4c 47 48 4b 51 46 49 52 4f 53 47 4b 4d 4c 4a 44 40 4c 4f 48 4a 51 50 45 52 4d 50 52 57 59 5c 5c 51 55 50 5b 59 5c 5b 5a 58 53 56 52 53 56 4e 52 58 4a 4b 49 4b 44 3a 1d 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0d 15 0d 13 23 29 33 3d 46 48 47 50 4b 4e 44 47 4c 42 41 49 45 46 46 42 4f 4a 4f 44 4d 49 48 4b 45 4c 4c 4a 45 51 4c 4c 47 4b 4f 4d 4a 4c 53 4c 4e 4b 4c 47 4f 45 48 49 46 49 4b 4c 42 4d 52 4d 4e 50 4e 51 50 5b 54 4c 56 51 5a 5e 50 55 53 4f 4e 59 4f 4c 4d 5a 5a 5b 59 5c 56 58 57 62 6a 58 54 4f 46 38 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 1f 43 47 57 59 59 4e 58 5b 58 4e 57 55 5e 51 60 54 57 55 65 55 50 55 56 4e 51 4e 52 55 58 55 59 4e 5a 5f 53 52 4b 4a 49 4c 4d 48 46 49 3f 4b 47 47 51 49 45 47 4f 43 4c 50 4b 57 4a 46 4f 4a 4b 43 49 4a 4c 47 4b 50 48 52 50 56 54 4b 56 4b 54 50 58 53 55 56 5b 5b 5d 5e 5a 59 58 58 5a 54 53 52 4b 4f 54 55 56 4f 4c 5a 51 40 35 1e 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 10 1d 19 2a 3c 3f 45 4b 4b 46 3d 46 3c 46 4e 45 4a 44 4c 42 4c 44 49 45 4a 47 4c 4c 49 49 43 4f 4a 44 4d 59 55 52 4e 4b 43 4e 50 4c 4a 4c 45 43 4b 42 4e 49 46 4a 49 47 49 50 51 57 46 40 4a 47 52 50 4f 4e 4d 50 51 51 5e 4f 48 4d 4f 56 54 54 4e 56 58 51 4c 4b 4e 4a 50 55 63 6e 65 5e 4a 48 3b 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 37 4f 54 4e 47 51 51 56 53 4a 52 55 5e 54 54 52 50 52 54 54 53 4e 58 4d 50 54 56 52 56 52 50 49 57 4b 54 55 4f 52 4d 43 51 49 44 4a 4a 4c 4c 4c 4b 48 4e 4e 4a 53 4d 46 49 4b 51 43 45 43 4d 46 45 4a 47 45 4b 47 4b 4b 4b 4b 58 4e 50 54 4e 5a 56 52 5e 53 5a 56 5b 5f 5a 54 61 56 54 4f 48 50 52 4b 47 45 54 53 53 52 44 3f 2b 0b 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 13 13 1a 2b 34 3f 48 4c 49 45 4a 4e 43 4a 41 43 46 45 45 48 48 3e 4c 46 52 44 47 48 49 44 41 41
 42 4a 56 55 60 51 48 45 4b 4b 4a 4b 43 46 42 44 53 45 43 4c 44 49 4f 47 54 44 43 47 48 47 48 46 53 49 4c 52 53 4b 50 56 54 4b 56 49 48 51 48 52 4c 4a 52 55 59 4e 51 52 57 4f 54 5f 60 5c 4a 4b 3d 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 40 49 51 49 4b 49 48 49 4e 4e 57 4c 5e 5c 58 50 53 55 54 5c 53 56 52 50 5b 4d 54 4f 4f 50 51 50 50 53 49 50 47 41 47 47 4f 50 4b 3d 47 53 45 4a 4a 3f 4d 4a 42 50 45 4d 4a 4b 4f 42 4e 49 49 48 4b 51 48 47 47 45 47 4c 55 45 4e 4c 4f 4e 4e 4c 52 62 59 5a 53 59 56 58 59 5b 54 50 50 51 54 4c 42 4f 4f 4d 4f 51 48 4d 3d 36 1c 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 0d 12 20 23 23 2e 46 3c 44 4c 50 42 44 47 4f 42 47 44 50 3e 41 48 40 49 4b 51 4f 4e 4b 48 47 44 3e 47 4d 4f 5b 59 52 4a 48 45 46 4c 47 46 4b 43 44 42 41 48 4b 45 4f 53 49 4b 46 49 47 4c 45 48 45 4c 49 49 4c 4c 4e 4d 53 51 4d 52 56 51 4e 4d 55 4d 51 4b 51 4a 59 4d 4e 4b 51 55 5d 5e 5a 4f 4d 3a 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 36 42 4d 49 4b 51 4d 57 54 4f 52 4e 4f 50 51 57 57 57 4e 53 59 54 57 4d 5c 58 5e 4a 4b 55 52 4c 53 50 54 4e 45 4d 4a 49 4e 49 51 45 50 45 4e 50 4b 4c 47 53 4b 49 4a 51 4a 4f 47 46 4c 3e 4f 49 46 56 4b 3e 44 48 55 55 54 4d 4c 47 51 4f 52 56 52 57 5c 57 58 62 5b 56 53 55 58 57 50 54 54 54 46 50 4e 4b 4d 4f 4b 4c 41 2c 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 16 13 20 28 2f 41 44 44 4d 45 43 4a 48 47 45 3f 4a 4a 45 47 41 4c 48 4a 4d 46 50 48 46 46 4d 40 3e 4f 49 51 53 50 4a 4a 4c 49 48 4f 4c 49 42 48 42 3e 41 41 3d 47 46 4a 46 45 4b 49 44 47 43 49 50 4e 50 4f 55 4a 49 4b 4d 4a 56 4c 50 49 4c 4b 48 4e 4f 4c 49 4f 43 4e 4b 48 4c 51 52 50 4e 4b 40 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 30 49 45 4b 50 4e 4e 4e 4d 4d 56 51 52 54 51 57 4f 53 54 50 58 56 59 4e 58 53 57 51 48 54 4e 4c 4a 49 51 43 50 4a 51 4b 4f 4e 49 4b 4a 40 49 49 4c 4b 4d 44 40 4f 4c 4e 50 4d 45 49 4b 4a 47 4a 41 3e 49 48 56 47 50 4e 4f 49 54 4c 47 4a 4f 60 53 5a 62 57 53 55 4f 52 4e 4e 53 52 51 55 5c 4e 4b 51 49 4b 4d 4d 51 45 3b 28 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0a 15 19 20 2b 3a 4a 44 4a 4a 3e 46 45 4a 49 48 3f 4d 41 45 44 4b 49 45 4d 47 4d 4b 4a 46 40 45
 4c 47 43 47 46 4f 48 4a 45 42 48 4b 3d 3e 45 4c 40 44 43 49 3d 48 45 44 47 42 43 49 46 43 42 46 45 48 48 4b 46 47 4b 4c 49 4b 50 4b 48 48 49 4e 4c 45 4a 46 45 48 51 46 46 46 4c 4f 4a 50 3e 45 38 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 30 4a 3a 47 41 4a 52 48 4e 4c 4e 4f 4e 4f 51 4c 58 4d 5d 49 53 53 53 52 4e 4f 4b 4b 55 4d 49 4c 4e 45 44 42 43 50 45 46 46 47 43 4b 43 44 49 44 44 44 45 48 44 4a 4a 4a 45 41 42 3f 4c 48 48 51 4b 4b 4e 44 45 40 48 4b 50 4d 4e 50 4e 4b 58 59 53 59 51 55 5a 53 54 55 56 56 50 52 53 52 45 4e 49 4f 51 4d 4c 49 43 48 32 23 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 0f 1e 1c 2d 3a 45 47 4d 4a 44 44 4b 49 49 4a 48 4a 41 45 4a 4a 49 4a 45 43 49 49 45 47 48 50 42 40 42 41 40 48 45 44 48 4c 45 3d 39 47 4a 47 48 3c 43 4d 42 3d 49 42 41 46 45 4a 45 45 42 4f 49 48 41 42 48 49 49 4e 4e 48 4e 49 46 50 40 4c 49 44 43 4a 49 4b 4c 43 3e 47 40 4a 45 4a 48 42 3e 2a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 28 47 44 4a 41 4b 49 47 4c 4d 54 4b 4b 4f 4b 51 53 51 50 4c 52 4d 52 53 51 57 49 4d 53 51 54 4c 5a 42 47 48 4a 4f 4d 48 44 4a 43 45 4a 4c 4b 4c 4e 3e 4b 47 4b 52 4c 4a 50 4e 52 48 48 47 51 50 43 48 48 45 4e 48 4d 50 53 4d 58 4e 4f 55 4c 4b 5a 56 5d 51 5b 5c 54 59 5a 4b 57 4b 56 4f 51 52 4a 46 46 43 50 4a 46 46 26 1a 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 13 25 2b 3c 3b 3e 4e 47 43 48 3d 49 43 4a 42 41 49 49 42 44 49 4c 43 4b 49 46 47 41 43 4c 4e 4e 3d 40 45 45 41 43 43 48 3e 47 45 47 4b 49 4a 45 43 47 3d 46 46 41 44 42 41 4a 47 4e 4c 49 46 48 47 41 44 43 47 4c 4a 45 4b 50 49 50 41 4a 48 44 42 45 3a 4c 42 48 41 47 45 44 49 41 3a 35 36 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 20 3f 4a 44 48 45 44 4b 4b 4b 4d 4b 4c 53 54 4b 4e 49 52 4d 52 56 52 51 4e 53 56 4b 4e 55 4e 4a 52 49 4b 47 4e 47 4f 41 4b 4b 44 46 44 41 4c 47 4e 51 4a 4b 4a 50 4f 44 4b 4c 4b 4a 4c 48 45 4e 4b 4a 48 44 53 50 48 51 4f 47 52 4e 53 51 59 54 52 59 5a 51 58 4e 50 5b 52 56 4d 4a 4d 4c 48 4b 4c 4f 4b 4e 4f 44 4e 39 1e 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 02 19 1d 21 2c 3e 4b 47 44 4b 49 45 42 48 46 45 48 43 47 3b 3e 41 47 43 42 43 49 49 46 47 44
 3d 47 3b 3e 3c 3e 3f 42 43 4b 42 40 44 45 45 45 40 3d 4a 48 40 44 45 3d 3c 3f 38 40 3c 46 3f 43 42 41 41 44 41 4a 44 4c 45 43 46 4a 43 48 44 46 44 3d 43 3e 43 41 3d 3f 41 41 47 3f 40 44 42 35 37 1f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 44 4e 3f 43 49 49 4f 46 40 4d 44 4f 4c 54 52 4e 53 53 58 55 50 57 55 51 4e 4e 4a 4e 4c 48 4d 4e 40 50 47 46 43 47 46 46 47 47 43 44 4d 45 48 48 4d 4c 49 49 41 57 48 45 49 4d 44 49 49 4e 51 4d 48 44 46 44 4f 4b 4c 4d 4a 4c 46 4e 52 53 52 4f 52 5b 52 52 4e 4b 4b 51 46 4e 50 47 50 4b 4c 44 45 48 3d 4c 4d 35 29 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 12 14 22 2f 37 41 49 48 48 3f 45 41 49 3f 42 48 48 44 4b 41 43 47 45 45 4a 4b 3f 44 47 40 44 43 39 3c 3a 3b 41 3a 44 3b 3f 3d 3d 41 44 3f 44 41 47 44 45 40 42 3e 41 3f 44 40 3f 43 45 3c 45 46 45 49 39 43 46 46 48 47 4c 47 40 45 4d 45 4d 41 45 44 46 3f 3b 36 3d 4a 46 46 45 3e 3a 3b 2f 1f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 43 41 45 3f 46 49 4b 4d 4e 4c 49 4f 62 58 59 5b 59 54 56 4e 50 58 50 4f 4f 4d 49 4d 43 47 44 45 4c 3f 49 44 4f 4b 3f 46 42 4d 3f 40 4a 46 4a 46 50 50 52 4f 4b 4b 4a 4a 47 49 49 53 4d 51 4a 43 4d 44 44 4d 4a 46 52 56 4f 4f 4a 4f 56 54 52 57 51 5b 51 4e 4d 4e 4a 56 45 58 4c 46 46 45 51 47 4e 50 43 43 45 35 2a 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 12 14 1b 32 38 3d 47 49 44 3f 45 45 44 54 49 4d 4b 41 3f 45 44 4c 41 41 4e 44 4a 4d 43 47 41 46 39 44 3f 3e 3c 41 43 4c 37 40 3d 3f 43 48 45 41 42 3f 3c 46 3d 3e 41 41 47 3e 3f 39 3f 48 40 42 4b 40 46 41 3e 40 43 4f 43 4c 3f 41 47 41 44 4a 41 42 43 49 40 41 3d 37 43 3b 3a 3e 39 3f 35 28 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 3c 40 3f 43 43 49 4c 51 4d 49 4e 5e 5b 63 62 5f 58 50 45 55 4b 54 50 56 53 53 4b 4e 48 4a 42 4d 46 47 4a 48 49 43 48 4d 42 48 47 4a 52 47 45 4e 48 49 48 46 4a 4b 4a 46 45 4b 40 49 4e 48 45 43 4a 47 4b 53 4c 48 49 5b 54 52 4f 4f 4c 4f 4e 51 4c 50 53 50 4d 4e 54 53 4c 4e 43 51 4d 4c 47 47 44 4c 40 42 3a 2b 21 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 08 14 15 2b 2f 3c 4b 4f 4b 4e 4c 53 4a 41 42 43 49 3e 44 3e 42 48 41 45 3d 44 3d 3d 45 44
 47 3e 45 40 42 42 3b 3f 39 35 40 44 3e 3d 3c 3f 4c 3a 48 42 43 39 3c 44 3e 43 44 3e 3a 3b 3c 3d 41 39 3f 42 3e 3e 3e 3f 43 4a 4c 44 42 3d 3d 3f 3d 3a 40 3e 40 47 3a 3a 37 3b 33 46 3f 3b 33 34 33 2b 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 3e 43 42 43 44 45 48 4a 50 54 60 66 66 6a 66 5c 4d 55 52 48 53 4e 52 52 49 48 42 4d 4e 46 4c 4c 45 42 45 48 47 4c 40 3c 47 48 48 43 4c 4d 4e 40 4d 48 43 4a 4b 46 48 4f 42 48 48 49 41 4f 44 4f 4a 47 4f 50 48 4c 40 4b 51 4b 4c 52 56 55 51 54 45 54 51 44 52 4f 4f 4b 51 4f 4a 4a 46 4a 4c 4d 44 40 3e 41 2f 25 19 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 11 14 12 1f 30 34 49 47 4a 49 47 46 48 42 49 50 49 46 3e 47 46 47 41 43 4a 44 4a 47 41 3e 43 3b 44 41 39 3c 3e 3b 37 45 3d 36 40 44 40 40 42 43 46 40 39 48 43 43 44 3c 43 47 39 3e 47 3f 44 3e 42 42 42 3f 4a 48 3d 40 44 3f 44 44 40 47 3e 45 44 3e 41 46 3d 3f 41 3f 3c 43 3c 3d 3e 35 38 2b 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 36 43 48 3e 3d 44 45 4d 49 4e 57 6b 6b 64 61 58 54 53 54 58 4b 54 51 4d 4f 4b 4c 51 48 4c 49 4e 48 47 47 4f 4b 46 3e 4a 47 42 4d 49 55 51 4f 50 44 47 4b 45 4b 4f 4a 4b 4b 45 4a 51 4b 52 47 43 53 53 4f 4b 48 4b 5b 4f 4e 4c 50 53 53 55 4f 54 53 53 4c 47 49 55 4e 4a 4e 44 4a 4b 46 4e 4a 42 40 4c 39 3a 38 21 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 0a 10 11 28 28 38 4c 47 47 4d 49 47 44 40 44 4a 3f 40 3e 42 41 3f 47 46 3f 40 3f 42 42 40 42 43 3d 44 3b 40 39 40 37 41 41 3b 40 42 3b 49 3c 3b 3e 4a 37 38 49 41 43 4d 39 47 40 3c 39 3e 47 3c 49 43 3a 3d 3c 41 45 41 44 40 3b 3e 3c 47 3e 41 43 37 40 42 3d 38 3c 3c 3d 45 37 47 3c 35 31 26 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 2f 45 44 48 40 4e 45 4f 4a 55 5e 64 6d 65 60 54 52 4e 4b 51 52 54 4e 4b 48 4e 44 50 49 4d 4a 4b 4b 47 51 51 4b 4f 44 45 4d 48 45 40 4b 45 47 49 45 43 52 4d 4c 4e 47 44 4c 4a 3b 52 4a 4b 4f 46 49 4f 4a 4a 4d 4e 51 4e 4f 49 51 4d 4f 4e 4d 51 56 50 50 4f 51 48 4e 4a 46 45 47 46 47 46 45 46 48 42 3b 31 2d 1c 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0b 11 16 25 34 3d 45 49 4b 40 41 3e 46 4e 3e 4c 45 48 41 3e 45 3e 42 3a 39 38 3f 42 41
 45 3a 3b 3a 41 40 3d 36 3b 3b 3b 3d 3d 40 44 43 40 3e 3e 40 34 48 3e 3f 3c 40 44 3f 3e 3b 44 3f 36 3f 3e 3e 46 3e 3d 43 40 44 41 45 3e 3a 42 43 42 39 3b 3f 39 3b 3c 3d 3c 38 39 3a 3a 3e 35 34 31 25 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 36 3e 3d 3f 47 47 47 4c 4f 5b 5b 61 6d 59 52 55 4a 4c 53 50 58 50 4b 4f 4e 4d 3e 46 4d 51 42 4f 48 45 4a 45 47 47 44 44 46 48 4c 46 48 4e 46 54 4d 4b 46 4f 51 4f 50 48 47 4c 47 47 50 50 4f 46 4f 47 46 4f 4d 49 4c 4b 56 4e 4b 4e 4f 46 50 51 4d 58 4d 42 47 4c 41 46 51 50 3d 4a 49 4b 49 39 41 42 36 2b 17 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 04 00 0a 07 11 18 21 33 3f 4d 51 4a 48 41 40 45 46 4c 45 49 3f 44 42 43 41 45 43 44 41 3e 39 3e 44 45 3f 34 37 3a 3b 3d 3a 38 3d 34 3d 3a 42 43 3e 3e 36 45 39 48 3c 38 38 39 37 3d 3a 3d 35 41 3e 39 3f 3d 42 41 41 42 3f 35 47 38 43 44 41 40 41 3f 38 3d 3c 32 3a 37 40 3c 3c 3c 37 35 38 31 2f 24 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 32 42 40 49 43 46 4b 52 4f 58 4e 58 57 55 51 4e 4b 56 50 50 48 4e 4f 4f 44 4b 4a 50 48 4c 46 4a 48 4e 4a 4e 48 4e 45 45 50 4b 4c 45 4d 46 46 49 49 4c 46 46 4c 49 51 49 48 4d 49 45 49 4b 4b 48 50 48 49 4e 4b 4a 57 54 50 4e 50 4f 54 47 4a 50 48 52 4b 50 4a 52 4b 4a 44 44 45 43 47 44 48 42 42 3a 31 2d 13 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0b 08 12 17 1f 2c 3c 3f 3e 3f 46 46 48 49 46 44 48 46 42 44 44 42 43 43 47 41 3d 3f 47 42 3f 3c 47 43 3a 38 39 3b 3b 3d 3a 3d 43 38 3b 41 45 3c 3e 3c 3f 3d 40 3d 39 40 39 43 3b 3a 3d 3e 43 39 3b 40 40 3a 3c 3e 43 44 3e 3b 45 39 35 41 3f 42 3a 3d 3c 3a 34 37 3e 3a 3d 3c 34 3b 34 2f 31 2c 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 35 41 42 46 42 47 47 50 44 53 49 4f 49 47 4c 51 4a 51 4a 4c 52 53 58 4c 53 51 48 47 46 52 50 4f 4c 48 48 4a 4d 4c 47 47 51 4c 43 4b 45 4b 4e 4c 50 48 44 4f 47 54 4d 4c 44 49 46 4d 53 52 52 54 49 4c 4a 51 4f 54 48 52 4e 51 50 59 4e 51 50 51 4a 4f 4d 4c 4b 4a 4b 4a 4b 4a 4c 49 47 45 44 47 3e 3b 33 23 14 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 18 20 31 41 42 3e 43 4a 49 46 4c 3d 42 47 40 45 41 40 41 4d 47 40 47 3d 3d 44
 46 3c 41 43 38 3b 3e 3a 3f 3f 3f 3c 3d 38 37 41 45 3e 39 40 3e 40 36 35 46 3d 3e 3b 35 40 3c 3b 3e 3f 39 3d 37 3d 38 3e 44 34 34 35 35 35 37 40 34 3f 3c 35 41 33 3d 44 3c 3c 36 38 3d 3c 35 32 31 31 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 2a 45 41 40 4c 3c 43 42 44 46 4d 4c 52 4d 46 50 4a 51 49 4e 4e 50 52 4d 54 48 4c 51 49 4b 4a 51 4d 46 4e 48 49 49 44 42 41 44 4d 50 46 4c 4a 47 4a 49 4d 4d 4c 4f 47 4f 48 46 46 4e 44 4e 49 47 4a 44 4a 4b 4e 4a 4b 4a 48 45 4a 47 54 4a 4b 51 4e 4c 4c 41 4e 46 3f 46 49 49 47 46 49 4a 46 42 41 3a 23 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 12 2a 33 3d 3d 41 48 40 45 49 40 46 49 42 3f 3e 3f 44 49 44 3e 4b 37 36 43 35 41 3d 39 39 3e 33 3c 3d 37 3b 39 41 34 3f 40 42 39 3e 43 3b 3c 3c 3f 3a 3e 3c 31 39 35 3b 3b 3c 3b 38 3c 3d 3a 39 39 39 3b 34 40 3c 39 42 37 3b 34 36 32 35 3a 39 37 39 3c 34 3c 3d 34 34 37 30 36 27 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 2a 44 43 43 44 42 41 44 3c 3e 42 45 4b 49 45 49 50 4a 51 4f 58 4e 4a 4d 47 4b 52 51 46 47 4a 4b 47 47 49 50 47 43 47 45 4e 48 47 43 49 4f 4a 4c 53 51 4d 43 47 45 43 4f 4f 4d 4e 4d 4a 55 48 4d 48 45 49 4f 4c 49 4e 51 4a 4f 42 51 45 46 43 52 51 4f 48 50 41 47 4c 47 45 41 4c 4c 4e 47 44 46 3a 36 1f 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 05 09 12 17 1f 2b 3e 41 46 44 48 45 44 4a 42 47 43 43 41 47 44 41 46 45 48 44 45 3d 42 3d 43 42 40 3d 3e 3e 3c 39 3c 40 41 35 45 3c 45 40 39 46 41 37 41 3c 3a 43 36 3c 45 31 3b 40 3a 3f 41 3c 37 37 31 40 39 39 39 3a 35 2f 3e 3d 38 3e 3c 35 3c 2e 39 3b 34 36 3d 41 38 37 3e 39 35 36 35 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 28 44 3e 45 4d 44 49 4d 49 45 3c 48 47 45 4c 46 57 54 51 4d 45 46 51 48 51 50 47 4a 43 48 4a 4f 52 4a 48 49 49 48 4a 46 47 43 46 49 54 4e 52 4a 49 4b 4a 4b 50 49 48 4e 4f 46 4d 4a 4b 4d 48 49 4c 4f 4b 51 4e 4b 4c 53 4f 4f 48 50 4d 47 4d 49 4a 4a 49 4a 47 4e 49 44 4c 44 44 44 52 42 49 3e 30 2d 25 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0a 19 26 30 44 44 3f 48 3d 3e 47 4a 47 43 41 3d 40 3e 4e 3f 3e 45 3d 36 3b 45
 3d 43 33 3a 39 3e 33 3e 3e 38 3e 3b 3f 42 40 39 39 3f 37 39 3f 3d 3f 3b 3a 38 35 3b 3a 3d 3f 40 35 3e 3d 3d 34 39 3c 35 39 31 3b 30 35 3a 36 35 38 34 35 3a 36 39 38 34 3a 32 3c 34 30 39 36 39 37 2e 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 25 39 41 45 41 4c 41 41 41 4a 42 4b 45 46 4f 4a 4d 44 4d 49 45 4c 4d 53 47 46 46 4c 49 4e 54 41 4a 48 52 4a 46 4d 40 4b 48 41 45 51 49 51 4a 4a 4b 54 4a 4a 4b 50 4d 4f 49 50 4a 45 4c 4a 52 4d 51 46 4b 52 4d 46 52 48 49 45 52 4b 45 54 47 4b 4a 51 4e 4c 45 40 46 42 4e 44 46 49 47 43 48 44 32 32 12 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0c 1c 1e 2f 41 3c 3c 44 45 48 42 48 44 43 3c 43 39 40 4a 42 3e 41 3c 46 3f 37 41 40 40 40 39 42 37 3b 3c 38 37 38 3b 3e 37 35 33 33 34 3e 3d 3b 3f 2f 3a 39 39 39 38 39 36 3d 3c 3a 40 3c 35 38 3f 35 39 3c 42 3a 36 34 39 38 30 34 35 38 38 3c 3a 33 3a 35 37 3a 3c 30 36 34 33 2e 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 45 49 43 44 43 44 4b 41 44 44 4c 4c 47 41 49 51 48 4d 45 42 4c 44 52 46 4d 49 48 51 4d 4a 50 3e 46 46 43 3d 4b 4b 47 45 46 4d 4b 4a 46 49 4d 48 50 4c 48 4c 49 4e 4c 51 50 49 49 44 4e 50 51 50 4d 49 44 51 47 48 50 46 48 48 4b 52 45 51 52 4b 52 48 46 47 41 4a 4e 3c 45 4a 43 4b 42 4a 2e 31 23 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0b 0e 23 2b 36 45 43 44 43 45 41 4c 48 43 37 3f 44 3c 3f 4a 41 46 3e 3d 42 3d 49 44 3f 3d 3b 43 41 40 39 3b 36 3a 38 3f 3a 35 3c 33 3d 3a 36 3b 3a 39 3d 45 34 3d 3e 36 3c 39 37 35 38 3f 34 33 36 39 3a 38 31 30 3f 33 39 3d 3d 33 35 34 38 3b 39 31 36 30 44 3b 3b 33 30 34 2d 31 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 15 46 35 50 4e 3e 45 40 40 41 3f 45 45 3d 42 48 43 48 44 49 50 45 48 4c 43 4a 4a 49 52 4a 51 4e 47 4b 4f 4e 54 51 4e 43 50 4f 4b 45 49 46 4d 4e 49 4d 4e 4b 55 4b 4e 4b 51 4c 4d 47 49 4f 52 4a 4e 4b 4c 4f 4c 49 50 51 4e 42 46 49 3f 46 48 46 51 4d 50 47 45 40 40 3f 44 47 43 4e 53 46 42 39 26 1b 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0b 0f 18 23 28 38 3c 3d 4a 44 4f 4c 45 40 48 40 44 45 44 46 44 44 3e 45 47 3d 4a
 44 49 39 3b 37 49 3d 44 3a 41 30 39 32 3c 3e 33 39 3b 36 44 3e 34 39 3b 3d 36 3c 3d 35 3d 39 44 47 3a 40 3e 35 46 3b 3b 3d 3a 32 3c 40 39 2e 30 37 33 38 37 34 35 35 2a 3d 2e 33 36 38 3d 37 33 28 2f 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1e 39 3d 49 47 4b 49 3d 40 46 3d 48 47 49 4a 42 49 4b 44 45 42 44 47 4c 4a 55 48 51 48 47 44 50 42 42 49 46 4c 46 4b 4b 51 4e 4b 4a 49 4d 43 49 4f 35 56 51 49 52 47 49 49 51 4c 4f 4e 50 4b 4f 52 4f 45 4b 48 49 50 50 45 4b 50 4a 4c 45 46 50 51 50 52 4c 49 44 45 4d 4b 47 45 4c 4a 50 40 33 23 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 0c 1e 1d 2c 39 3c 44 4a 3e 43 4b 43 43 41 3f 3e 3f 37 42 41 45 42 3d 3d 3e 45 3b 36 3f 3a 41 3b 38 3b 3a 3a 40 37 34 39 35 40 3d 39 3e 41 39 3b 2e 38 37 3c 3e 36 37 3a 37 3b 38 39 41 3d 36 32 38 3a 3b 34 36 38 32 30 3a 3b 36 2b 36 2f 34 32 29 33 3b 39 3c 35 2f 31 30 30 29 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 3d 42 3e 42 48 42 3e 44 39 39 3f 43 38 40 3e 44 47 43 44 46 48 4a 46 48 3f 42 4a 4a 46 49 4c 4a 4e 41 4d 4b 51 45 4a 51 45 49 53 47 49 51 4a 4f 52 43 48 4a 49 41 4d 43 4d 52 51 4f 57 54 51 56 58 4e 4f 4e 4a 48 4f 44 56 4c 4c 4e 48 4d 4b 4c 4d 4b 4a 48 4a 4d 42 43 43 4a 51 51 40 3a 2b 15 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0b 12 27 2d 32 42 4a 4d 48 40 4b 42 40 42 38 40 3e 48 47 40 41 44 3e 43 41 3b 3d 41 3b 3a 48 3d 43 39 3e 3c 3b 32 39 34 3c 3e 40 37 36 3a 3e 3b 39 34 37 3a 33 3b 3c 42 37 39 39 3b 3e 39 39 3f 39 37 3a 2e 3e 3b 31 31 34 3a 32 35 36 37 36 32 39 2f 34 32 31 2d 36 33 31 2b 26 1d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 32 39 3e 44 44 40 40 3f 3f 3c 37 42 38 48 3e 38 45 3f 43 45 43 44 3f 47 46 41 4a 41 4c 42 4d 40 47 48 4f 4b 50 53 50 52 4b 48 4e 4f 46 4a 43 4d 49 44 4d 49 53 50 47 54 4f 52 60 59 5f 5a 52 52 54 55 4e 4c 4f 59 53 55 57 55 4e 53 4c 48 4b 47 4f 48 49 52 42 4a 4b 47 44 4b 49 45 43 37 20 18 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0f 14 1f 2b 32 41 40 48 44 4a 44 49 47 44 44 45 4b 45 4a 45 4a 4c 44 46 3f
 3d 42 40 3c 3b 43 3a 3c 3a 3d 39 3f 3c 35 34 37 3a 38 35 3b 33 38 3d 37 41 34 37 38 3a 3e 43 41 3b 3c 3b 45 38 37 33 3c 36 33 37 3c 3d 3f 31 36 36 36 2f 39 3b 31 37 39 33 30 3f 31 36 37 36 2e 2e 2f 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0d 2e 44 3d 42 3f 3b 3a 38 45 3d 3a 40 38 3c 41 3b 3e 43 43 3d 40 3f 40 42 46 42 45 42 48 45 46 4b 3d 4c 56 53 51 4e 50 4e 49 52 4e 4a 48 44 4b 47 54 4c 50 4c 45 4d 51 50 53 5c 68 6a 65 69 55 53 54 51 59 59 55 53 56 58 59 55 58 53 4c 4c 52 4e 43 48 53 50 4a 55 47 43 48 41 4c 42 37 2c 21 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 11 16 20 2a 40 46 46 41 4a 46 43 46 46 3e 36 3f 44 3e 4a 41 41 42 3e 3a 41 3c 43 3b 40 3c 37 41 43 3d 36 42 32 31 38 37 33 33 36 43 32 37 3b 2d 37 34 36 32 36 31 35 3d 43 35 34 3c 36 32 3a 38 3a 30 3d 35 35 3c 30 3b 36 37 2d 2f 35 37 35 35 3b 33 35 35 35 33 32 3d 31 2f 1d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 2a 37 36 2f 38 49 3e 3c 3c 36 3d 3f 3c 34 3d 39 3d 3e 3d 3c 37 43 3e 3c 44 47 45 43 44 44 44 3d 48 44 48 4e 49 52 50 4b 4e 45 47 4e 4e 4d 48 47 49 4c 46 4a 47 52 4e 55 5d 69 6c 65 64 5c 56 5c 59 52 57 4c 53 5b 5b 52 5d 59 53 48 57 51 50 50 48 4f 4a 45 49 47 49 4d 46 43 41 3b 35 1f 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 13 1b 26 2b 39 3b 3b 45 3b 4a 47 46 4a 45 47 40 4a 45 4b 4f 3c 49 41 45 42 43 40 3f 47 3c 41 36 35 4c 42 40 3c 38 3a 39 37 34 3c 38 3c 2b 37 36 3b 31 3e 41 3e 30 38 37 39 34 39 40 2e 36 33 2f 32 39 35 3e 33 3c 33 3d 32 33 3e 35 33 3a 3a 36 34 30 3a 35 39 33 2e 32 2b 27 26 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 30 31 3b 3d 3c 41 39 37 3b 36 3f 3a 42 38 3d 40 45 39 45 36 3e 45 3d 44 3c 43 3c 3b 48 47 4e 42 4a 4c 46 4e 54 4c 53 47 52 4b 4a 4f 4f 4f 3e 4b 45 4d 4d 51 4b 4e 5c 5e 6e 6c 6d 62 62 53 4e 4b 52 4e 4b 4c 58 4e 56 5b 58 5a 50 52 48 52 51 56 4f 44 47 4e 4e 52 4c 47 46 38 40 37 29 18 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 13 12 26 30 3b 44 3c 43 34 4e 49 42 41 42 42 42 48 46 40 47 44 3e 3f 43
 41 3d 43 3d 40 43 3b 43 39 36 3d 3d 33 3e 3a 3b 38 37 3b 3d 34 3a 39 3b 33 3d 34 35 34 2f 3a 35 38 38 3c 3a 38 39 35 3b 42 3e 3e 39 3b 40 2f 39 3b 39 35 3d 36 38 3b 34 37 35 2c 36 32 32 35 38 36 2b 2a 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 32 3a 3e 43 3a 37 3b 38 3d 38 43 35 41 3f 3b 3d 3f 3a 40 45 41 49 3b 43 47 3f 47 43 41 45 49 3e 4b 4c 45 4f 49 4a 4d 4f 54 4e 4c 49 45 47 41 49 46 4a 51 49 4b 56 51 60 6b 66 5a 61 56 4d 46 48 4c 47 4d 53 51 52 50 4a 4a 4f 4d 5d 50 56 60 53 5c 4d 50 4a 4b 52 50 42 4b 45 38 3b 1c 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 18 17 25 30 39 40 40 41 40 3f 41 4f 3e 45 48 40 4b 44 43 3e 42 44 3f 3c 3e 38 42 41 3b 3b 38 3e 38 36 32 37 3d 3d 34 3a 3a 35 35 3a 2b 39 3e 40 3d 3c 3f 35 39 39 37 37 3f 3c 36 34 38 38 3d 3f 34 35 38 3a 3b 3c 3b 35 34 34 3b 3c 39 3b 35 30 3a 28 35 2f 31 30 31 32 2d 2d 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 35 34 3d 3a 3b 34 3a 35 2a 40 3c 36 35 3b 3f 43 39 36 38 41 45 43 3e 46 47 49 47 4c 40 41 46 43 45 3e 49 53 47 4a 4b 4c 4b 4c 43 4a 4d 50 4f 49 4c 4b 52 4d 4c 55 60 65 5b 55 55 53 4d 50 42 48 48 4d 50 4b 4c 4d 41 41 45 4d 45 49 52 5f 64 5a 4c 49 44 41 48 3f 48 43 38 3b 26 1a 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0c 0a 10 1a 2c 3e 3d 3f 45 47 45 46 40 4a 3e 42 3f 42 44 46 3e 3c 43 3d 3f 42 39 42 3c 42 3a 46 40 43 3d 44 38 39 39 38 36 37 41 30 35 35 29 39 36 36 36 36 37 3b 3c 3f 37 3d 36 37 39 40 37 3c 3e 35 3b 42 36 38 3f 37 3a 32 33 39 37 39 35 36 38 38 3a 3c 2b 37 2b 31 33 2c 26 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 3d 3d 42 38 34 39 3a 35 41 3e 3c 36 33 38 47 43 42 3f 46 3e 40 43 41 42 42 4b 47 4e 4b 47 49 3b 42 46 4f 49 4a 4e 48 47 48 4e 54 50 55 47 4c 52 49 4a 48 54 4a 55 66 5f 5b 56 4c 4a 47 3b 42 41 44 44 47 45 49 4b 44 36 41 4b 4a 50 55 5e 56 55 52 44 4a 47 4b 47 49 4b 3f 33 25 09 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 10 16 32 2c 33 37 3c 3d 43 41 4a 48 40 52 4f 40 46 4a 43 3e 45 44
 3f 42 3e 3c 3c 3a 42 45 42 43 36 3c 38 3e 3c 39 40 3b 36 3a 3e 33 35 39 34 36 3f 3a 38 3a 36 32 38 39 3b 3f 39 3a 37 35 40 3c 3a 3e 32 3f 32 3a 42 39 3b 42 41 38 34 3b 32 38 34 30 2d 2f 36 35 3e 35 34 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1c 34 35 37 37 37 41 39 41 47 44 40 3b 44 47 4b 45 44 49 4a 4b 48 50 43 49 43 3e 3c 44 49 45 4b 44 43 51 47 45 51 46 4d 4a 45 50 48 48 52 53 52 5b 50 4e 47 4d 52 5f 63 54 52 4a 4c 51 4a 45 44 46 40 46 43 45 43 43 3f 4c 4a 4a 4e 49 51 56 59 4c 49 43 4a 4a 47 4e 4b 4c 43 2f 12 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0d 14 1f 2e 34 33 3c 48 44 42 41 40 4d 47 4a 4b 42 45 40 46 45 47 3a 3f 41 3d 44 42 3c 41 44 3e 3b 3a 33 40 3a 34 3b 37 3b 3a 30 35 34 36 31 3a 32 36 3c 40 3b 35 34 3b 37 32 34 34 3a 39 3f 36 3a 36 36 3f 33 36 3d 36 35 3f 30 38 41 35 37 36 36 38 2e 39 34 31 36 32 2c 1e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 2c 32 39 30 3c 34 35 41 40 41 49 48 49 48 47 34 4a 48 49 4f 46 4d 46 43 4c 50 46 55 4b 4c 48 46 4c 4a 4b 4a 49 46 3f 45 4d 50 52 46 4a 4d 58 55 4e 4a 4e 47 52 56 58 50 4a 4e 46 45 46 3f 34 44 39 48 49 43 47 3c 42 44 47 4f 47 4a 4d 4b 4a 4b 48 51 53 54 55 4a 51 4a 36 21 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 15 19 2b 31 3e 36 43 48 43 41 46 46 3f 43 41 45 48 43 43 44 41 41 47 40 3b 40 3e 3f 40 4b 3a 3c 44 3c 39 37 3b 3d 38 3c 3c 37 31 3b 39 37 2d 32 37 35 37 36 33 37 34 34 3b 36 34 34 37 3c 36 39 3a 3a 3e 33 37 34 32 32 32 37 36 36 37 3b 31 3a 40 36 39 3b 2f 30 30 33 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 26 35 37 37 3b 3d 3a 45 45 4e 45 48 3a 3d 3b 4a 47 46 4d 48 4d 49 43 4c 4e 4b 4e 4c 45 4a 4d 44 44 4f 4a 40 48 4a 4c 46 4b 50 47 51 53 51 4f 4b 4f 4f 4e 4c 4b 4b 4d 45 45 44 40 48 44 43 49 42 3d 40 3c 40 46 3f 46 40 33 41 48 41 44 4f 4c 56 51 49 52 55 4f 60 58 45 35 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 08 14 14 22 32 30 33 3c 42 43 40 41 49 49 47 47 41 47 45 42 40 47
 3f 44 42 3b 3c 40 42 3d 42 42 45 47 3b 42 38 36 44 3b 3e 3c 37 3a 36 32 3d 39 3d 38 38 33 39 40 41 3e 43 37 3d 38 35 3e 35 37 3f 37 3e 39 32 39 3f 3e 3d 3d 39 37 33 3b 32 3c 40 40 38 41 3f 3b 32 33 38 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 2b 32 40 3c 40 3d 39 42 3b 43 4a 41 43 43 48 4c 47 48 48 4a 45 4b 4c 4a 48 4a 46 56 4e 46 44 41 4d 43 48 4e 50 4d 47 47 57 4f 56 53 4a 41 4d 52 4e 50 48 45 50 47 44 45 43 3e 4a 40 3b 41 43 41 42 40 42 44 4c 3c 3f 44 3d 42 43 4b 46 51 57 59 56 56 62 66 6c 58 54 4a 31 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 21 26 31 3c 38 45 44 45 41 41 44 47 44 4a 4c 3f 4e 43 41 40 41 3e 41 3d 45 45 45 43 42 3d 42 3c 40 3d 40 34 34 36 3b 34 31 41 33 3c 36 36 33 32 3b 38 39 3e 35 32 3d 33 35 37 37 39 34 40 3b 3a 3a 3d 40 39 40 3e 36 3e 3b 41 37 3e 40 3e 45 3d 46 3a 36 34 30 2e 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 2d 39 42 3a 40 3a 40 43 3a 3d 3c 39 41 42 3b 45 47 43 46 4d 38 43 47 45 4b 41 4c 4f 4c 4f 4e 45 4f 49 4c 4f 4c 4a 4b 54 4f 43 56 4d 53 47 41 49 4e 42 52 44 4b 4d 41 47 44 45 3e 44 4b 3c 44 45 39 3c 3f 3a 42 42 4d 44 44 49 46 50 5a 5e 65 68 66 78 69 6a 66 53 54 37 20 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 19 1b 28 38 32 37 3c 42 3e 43 47 3e 41 44 42 49 45 45 42 42 42 3f 3b 42 3f 39 37 44 3a 45 41 3c 39 3e 45 3c 37 30 39 3c 3a 3a 32 33 2f 30 37 38 31 37 36 38 39 39 38 33 30 38 3b 37 3b 3e 3d 41 3a 36 35 3e 35 36 33 31 35 3e 43 43 3d 3f 3d 3b 40 38 3e 33 2a 24 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 2b 35 41 3a 38 3d 3e 40 3a 42 38 33 3d 3c 34 42 42 4a 4a 49 44 41 44 43 3d 44 45 4c 4f 4c 40 4c 3f 4b 48 45 50 46 4c 42 49 47 48 44 44 49 4a 49 3a 43 41 3c 44 41 45 41 3d 46 44 46 45 43 3a 3c 38 42 4b 4d 46 46 38 54 45 4b 60 53 6c 6d 76 79 75 79 6b 69 60 54 46 2b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0b 19 29 2b 3e 3b 3a 40 3e 44 45 40 4c 4d 45 41 45 3e 3e
 40 45 3e 40 3c 46 3e 45 3d 41 43 42 3e 3d 38 42 3b 3b 3a 39 3a 3b 32 38 34 32 38 36 32 38 35 3a 3a 34 3b 40 34 38 3b 36 42 33 42 3d 38 3a 33 3c 41 3c 3d 37 3a 3f 3e 46 42 3c 41 3f 37 42 33 33 29 23 2b 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 2e 40 3d 37 40 3a 39 42 31 32 3e 3c 38 39 3d 3c 43 3f 3d 43 3d 49 41 43 41 41 4a 45 47 4a 42 45 46 4a 49 4c 4c 4a 45 45 45 45 46 41 49 45 49 46 46 45 41 46 3d 3a 42 43 3d 42 46 40 42 44 3d 41 41 3f 40 47 4f 4f 4d 53 55 62 68 73 7c 76 77 6f 42 5e 68 69 59 49 35 15 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 1d 25 38 33 39 43 3f 40 44 41 46 47 36 47 44 3c 4c 41 44 42 48 3e 39 43 44 44 40 4a 41 40 43 3c 4d 40 39 40 33 38 34 3e 39 35 31 36 36 39 30 36 35 36 3e 3c 33 3c 3d 39 3a 3f 39 39 3b 32 38 3d 3a 39 39 39 3d 40 38 42 3b 3e 45 49 39 36 39 36 29 2d 2e 2c 26 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 36 39 37 38 3b 3a 3e 3c 30 30 3c 37 3b 41 38 3f 32 3d 3c 40 41 41 42 36 3d 3f 40 41 3e 45 44 42 44 3c 43 42 48 41 45 45 4a 4c 49 3e 45 43 40 45 3c 3c 44 44 3d 3f 40 3d 3c 4b 3f 50 42 4b 40 49 47 50 55 57 67 59 5b 6e 6e 75 7a 7c 76 7f 78 78 70 69 55 5e 4a 34 27 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 11 18 25 31 36 34 37 41 40 3c 41 40 44 4a 45 44 49 46 49 44 46 41 44 45 44 40 44 3e 3e 45 44 4f 50 41 40 39 41 3b 3a 33 27 36 36 3b 32 2c 37 31 35 35 38 38 37 34 3d 37 32 39 3a 3d 3b 42 3d 33 38 37 3d 36 3a 3a 38 39 41 3d 34 3b 3d 3c 2b 35 36 2a 2b 2c 28 23 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 22 30 3f 3a 37 30 35 35 33 3c 38 36 2b 38 39 37 38 35 3b 37 33 3b 3a 3c 3a 3b 3f 44 3f 42 3f 41 3c 46 3f 43 44 43 49 47 4a 3f 3a 3f 43 46 47 48 43 47 3c 42 4b 44 44 3c 3f 44 44 4b 4a 4d 59 54 54 5d 63 70 71 76 77 7c 78 7b 7e 7c 81 72 79 72 65 69 54 48 3d 2d 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 15 22 2f 37 3d 40 35 36 42 39 47 41 3e 3f 40 47 46
 4b 48 3b 42 45 48 3f 3f 45 4a 4b 4a 4f 54 52 4f 47 44 45 3a 35 35 35 37 3e 33 35 30 29 35 35 39 3d 34 38 3b 3b 37 36 42 31 36 3a 38 34 33 31 36 40 3d 44 3c 41 3e 3e 44 3a 36 3a 32 31 35 2e 32 2d 2f 29 1c 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 27 31 34 33 34 31 2a 3e 36 3c 39 38 38 34 3e 36 3b 35 36 3c 3e 3e 39 35 3c 3c 36 43 41 40 3e 42 3e 43 42 45 48 40 42 3b 3d 41 41 45 46 42 49 3e 46 3d 40 44 4c 46 4c 55 4c 5b 54 55 58 59 60 67 6c 6f 73 74 74 7f 83 7d 7b 82 7b 7e 7e 6e 76 6e 63 5c 4c 41 2d 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 1c 28 30 2f 34 3f 3b 43 3e 3c 3e 44 3d 42 45 40 40 3e 3d 44 47 41 44 47 3d 46 44 49 4b 55 58 57 4b 52 40 40 36 39 39 3a 39 32 3a 33 39 36 39 3b 39 36 3b 40 2f 3a 39 32 32 3b 3b 3d 37 43 35 3c 39 38 42 42 38 44 39 3c 3c 34 35 32 31 2b 28 35 25 2e 2a 29 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 33 35 3b 35 30 2f 33 32 32 38 32 36 3a 32 39 34 3a 3b 3d 3c 3c 3a 40 3f 38 37 39 3c 47 40 3e 3d 3f 40 4a 43 3e 3f 42 47 45 48 46 43 49 44 45 45 47 4a 4e 4c 51 51 51 4f 5e 65 71 6d 6c 76 75 75 7e 7c 7e 7c 7b 73 7f 76 81 75 77 6f 71 73 61 59 57 3e 2b 21 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0e 15 23 32 36 39 3a 3f 39 37 38 3b 40 3b 44 4b 41 4d 48 44 42 46 41 41 41 43 49 3c 46 50 55 65 5a 54 5b 52 4c 42 47 3e 36 42 3b 3e 39 39 39 31 3d 36 3e 36 38 3e 30 30 38 32 35 38 38 3c 3b 39 41 3c 3a 3e 3b 41 3b 3d 38 33 2e 36 33 2d 30 2b 2b 2b 29 2d 24 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 31 31 39 31 2e 32 38 32 37 34 35 3b 3b 36 37 33 37 36 36 3b 35 36 3c 38 3e 39 3b 40 3d 40 37 3e 3f 3a 46 44 3f 3f 42 46 47 47 4c 4f 4c 4d 4e 49 4c 56 55 5e 51 61 66 6d 6e 72 70 77 75 7c 7e 79 75 80 7b 78 7a 70 79 72 77 7e 6d 6e 66 64 5b 52 40 32 1c 0e 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1a 26 2b 3a 3c 41 3b 3c 3f 3a 3e 4a 47 43 43
 4b 46 49 4d 39 4a 43 48 47 51 45 49 4f 56 58 63 5f 5d 5c 56 46 46 3e 40 42 44 40 3e 3a 3f 3b 40 34 36 3c 40 33 36 38 37 3e 33 39 37 33 3f 3b 40 43 39 43 3d 39 3b 39 3a 33 2c 34 37 3c 2e 2c 2b 2a 2f 28 25 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1c 2d 30 3b 3b 32 31 36 2b 33 39 37 32 37 31 34 33 3a 3b 40 36 3e 36 36 3f 42 34 3c 34 40 3c 3f 3f 3c 42 47 47 4b 4c 4b 4d 55 4f 4f 59 57 57 59 5a 61 64 62 6e 6c 74 76 78 7b 79 83 85 7e 7e 72 77 80 80 74 7b 7a 72 78 6e 6b 71 69 63 61 5e 53 3d 34 1e 0c 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0e 16 2d 36 3b 41 3a 3f 3c 3a 43 3d 42 3b 41 41 4b 47 43 45 44 44 45 46 4b 48 48 50 52 51 62 5a 5c 5e 57 4d 4d 4f 48 4d 43 4b 45 45 46 3d 44 43 43 42 39 3a 38 37 31 37 32 36 3a 3c 3c 38 37 3f 40 38 3f 41 34 37 2f 35 31 2f 36 34 35 2d 2a 2e 2b 26 24 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 2e 30 3a 34 34 27 36 2d 2c 2e 32 34 2f 3f 38 2b 32 3d 35 39 3c 39 41 41 38 3a 3e 3a 39 41 39 40 4c 40 44 49 54 4c 57 5a 5a 62 6b 68 68 60 6c 6e 70 76 75 7f 7d 78 7e 7c 79 7b 7d 80 7d 7e 76 7c 7c 73 75 73 76 76 6d 5f 6c 64 58 5f 5a 52 45 2e 26 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 12 24 22 35 3e 3c 3c 3d 3c 38 3c 3b 36 3c 44 4f 3e 46 3e 48 47 3d 44 48 43 46 44 50 49 4e 49 56 50 55 50 4b 50 4d 48 4d 42 4d 4b 40 3f 43 3e 3f 3e 3e 3c 38 30 37 35 2d 2b 39 35 38 3d 40 3a 36 34 39 37 3f 30 2c 36 2a 2a 26 30 30 2d 2c 29 26 23 24 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 32 2a 29 31 36 30 35 2b 2f 2d 2e 30 35 36 36 2f 2b 33 38 37 3a 30 39 39 39 35 39 3c 40 39 39 3d 4c 4e 54 56 5e 59 6b 61 65 6b 6e 74 6f 77 7b 7b 7a 7b 7b 7c 7a 79 7e 7b 76 77 76 75 6d 74 79 6e 6d 74 68 6e 7a 6e 66 5f 5f 60 5a 52 4e 44 37 28 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 1d 26 2f 36 3e 3f 46 41 41 40 39 44 3f
 3f 42 44 46 41 46 40 45 41 46 40 3f 41 49 4c 4c 48 4c 57 4c 51 4e 44 47 4c 46 43 43 40 46 47 41 3c 3a 3a 3d 3f 3e 32 31 35 34 35 3d 38 37 2a 38 3d 3b 3f 42 31 39 2e 30 33 32 29 28 2b 2b 2f 2e 2c 29 26 2f 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 2b 36 2b 2e 31 2c 38 32 30 35 32 33 2b 31 2b 34 36 35 32 38 30 2a 2f 3d 3d 36 39 33 45 43 45 4c 57 5d 64 6a 6f 77 76 70 71 7c 80 79 76 87 79 72 7a 7f 7f 78 79 7c 7e 77 75 76 70 74 6e 75 66 6b 69 5e 63 5f 65 67 60 56 5b 57 55 4e 3e 38 30 14 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 15 1b 23 3a 30 42 3b 38 47 40 3f 45 3f 42 48 44 43 41 44 3a 47 43 4b 43 3b 42 45 3d 3f 49 42 44 4d 44 49 40 46 43 3d 3f 41 46 45 40 3a 37 41 3a 3f 34 3c 38 39 43 39 3c 35 35 3e 3f 37 3f 34 34 36 32 31 33 30 2d 33 34 35 32 32 2f 22 2e 27 28 24 16 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 23 30 2e 33 33 2d 33 2e 2d 35 36 2c 3a 30 34 33 2f 32 37 32 35 36 34 34 35 40 42 3d 41 4a 58 5c 65 70 71 6d 73 74 6f 83 7e 7c 7f 7d 79 84 79 79 7d 78 79 75 7c 77 75 77 6f 76 69 73 6e 6e 4f 62 61 62 62 68 5d 5e 5f 57 50 4b 4d 45 3a 2a 17 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 24 28 34 38 3f 3f 3d 3f 37 3b 36 46 42 3e 44 42 44 42 39 3c 42 3d 47 41 45 3f 47 3d 4c 44 44 40 3e 42 39 3c 44 3c 40 37 38 38 3e 35 38 36 2f 22 38 30 39 38 34 36 39 3a 35 3a 31 33 31 32 3a 30 33 35 27 2e 2a 27 2f 30 2c 1f 24 2c 29 31 23 1b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 29 21 2c 2a 2c 25 34 23 3b 36 28 2d 2e 2f 38 3a 34 30 33 33 31 32 39 3e 39 3c 4a 46 53 63 61 73 75 76 79 78 73 81 76 7a 78 77 78 77 70 76 7c 7b 73 76 73 6e 73 67 68 69 66 65 6c 60 61 69 60 68 62 58 59 5b 58 51 59 49 46 3f 3b 33 27 17 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 17 22 38 34 36 3a 46 3d 42 3f 40
 3d 44 42 3e 3d 3b 3d 3c 3e 3d 44 41 44 3f 41 3b 36 42 40 47 4e 4b 45 3a 33 34 38 3b 38 3a 36 3d 37 39 39 38 2e 27 2b 34 35 3d 31 2d 2e 29 36 34 2e 2c 32 2e 32 33 32 27 2d 30 33 38 2c 29 2d 27 26 29 28 25 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 2b 2f 2f 2a 23 26 30 2b 24 2f 28 2a 31 28 2d 37 2b 2d 35 2f 3a 41 3c 41 41 50 52 68 6a 6e 73 7a 78 75 7f 76 7e 80 7a 79 6e 7a 7d 79 7a 70 6e 6d 6f 6f 69 70 6a 6a 62 62 66 61 60 58 65 57 5b 5e 55 4e 55 51 4e 46 45 44 3e 3e 2a 20 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0c 19 2d 31 40 38 42 40 41 40 3a 42 38 3f 39 3c 42 3e 3e 48 43 3d 3e 43 3e 44 47 3b 3c 41 4a 45 4d 48 42 3f 3d 3e 37 2f 34 35 42 3c 36 37 34 31 2e 32 32 33 28 32 2f 2e 33 34 2c 2d 2a 2d 2d 30 31 2e 22 2e 2f 36 32 2a 2d 27 2b 27 2a 27 26 1d 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 27 29 2f 34 2c 28 2b 2f 2a 2a 2d 2f 2f 2e 2f 2b 35 33 35 26 3a 3d 43 4f 5c 5f 75 70 66 7c 75 7f 76 76 78 78 77 76 74 78 6a 71 76 6a 7a 6e 66 6f 6c 6b 6b 65 69 67 6b 65 5b 64 5b 5e 5a 56 53 5b 57 51 55 50 4e 48 43 3e 3b 2c 1b 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 14 22 28 35 37 38 3f 3f 3e 3c 3f 41 44 3d 3c 46 3d 44 3d 3a 3f 3e 40 41 44 46 41 43 45 49 40 4b 3e 43 44 39 3b 32 33 2f 35 37 3c 3a 3f 36 27 2c 2a 2f 34 2a 27 32 2c 26 28 2c 2d 2f 29 2b 2e 2f 34 2f 2d 2a 33 2f 28 34 29 25 2d 25 21 24 11 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 24 27 2e 27 29 2d 27 2a 2b 24 2a 30 2a 2e 2c 2c 2a 31 34 37 3c 45 48 5a 6b 6a 72 70 75 76 74 76 76 78 72 6e 6d 67 68 6a 68 6a 6c 66 6b 68 65 66 6b 63 5a 61 5e 5a 5a 5b 55 5c 59 54 50 5a 47 46 4c 48 5a 49 4b 44 3d 37 2b 1b 0b 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0d 1e 2f 34 3b 36 36 3b 3a
 3f 3d 35 3f 39 38 37 3c 45 45 3d 3d 3e 3a 37 43 3d 48 3e 43 44 48 49 3c 3f 36 34 36 37 27 2a 3f 35 38 39 3a 34 2f 27 2a 2d 29 26 2b 2b 30 21 28 22 27 24 21 28 2b 2b 2a 2f 2d 27 2f 2e 31 26 2f 24 21 25 24 1f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 21 28 22 2a 2a 28 20 2b 25 1a 2a 2e 24 30 2c 23 27 2d 35 36 47 5e 52 64 6f 6e 66 6f 66 64 69 64 6c 6c 62 62 66 69 66 5e 6a 65 66 5e 5f 69 5b 60 5f 5b 59 58 52 50 55 52 4f 56 55 46 48 46 50 51 4f 48 45 41 39 3d 24 1f 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 1a 21 2f 3a 3e 41 3e 41 3b 3c 3f 3f 3b 46 3d 3d 42 40 40 3c 39 44 3e 37 41 3f 3b 43 37 44 48 42 3d 3a 35 39 3f 39 3a 2c 30 30 3b 36 2c 26 2e 32 2c 2a 2d 27 1f 28 22 2a 25 21 20 23 27 2b 2a 26 31 25 31 2c 24 2c 26 2c 23 25 22 24 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 17 22 23 21 2f 29 25 25 26 25 23 2c 2c 31 27 2f 25 32 3d 4b 59 5a 60 65 63 63 67 68 62 63 61 64 64 5e 5b 5e 56 51 64 59 60 54 5c 5e 59 52 53 5b 5d 59 52 52 50 53 49 4f 4d 4d 42 45 43 4a 43 4d 4d 3b 40 3b 2e 28 1a 1b 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 1d 29 32 37 32 36 39 3d 41 39 3f 43 3f 34 36 3e 47 39 38 3e 43 40 3e 3d 3c 42 44 3b 46 40 3e 3d 36 32 39 37 2e 34 38 3b 2f 2f 33 32 32 2d 25 26 20 27 27 24 20 15 18 22 1f 1a 25 22 2c 28 2a 2e 2e 1f 2c 25 27 29 23 23 20 28 23 13 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 12 1a 22 1b 18 1e 1d 1e 1a 16 1f 1d 2a 20 21 2c 37 36 3a 46 53 58 57 5c 55 5b 56 56 52 4b 4b 50 58 4d 4c 4c 4e 50 52 4a 4d 4b 4c 4a 49 49 44 44 45 44 43 47 4b 41 3f 4a 48 43 45 43 42 48 3a 36 3a 37 37 2d 26 16 08 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 1a 26 28 38 35 35
 40 40 36 36 37 3c 3d 38 36 3a 37 38 34 39 3c 3a 38 3a 3e 43 43 47 41 34 37 39 33 31 37 29 2d 33 39 2a 2c 32 24 25 25 24 29 22 22 22 16 14 07 13 11 13 17 1c 1f 24 27 24 25 1c 21 25 16 21 24 23 1f 18 18 1d 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 12 14 10 0d 16 13 16 14 15 19 15 18 1e 21 2a 29 43 40 3c 44 41 40 36 43 41 38 36 2e 3b 36 35 37 35 36 32 31 31 32 35 3a 36 3b 35 41 32 34 35 33 37 33 31 35 30 31 30 3b 32 35 36 32 30 34 30 25 1d 12 0f 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0d 23 1c 33 36 36 37 38 37 39 41 41 36 39 38 38 3d 37 2f 38 3b 43 3d 37 44 40 46 46 4a 40 3d 3d 31 2f 2f 2b 2b 35 30 27 33 2c 37 2d 23 27 25 1f 1e 1c 0e 0a 06 0d 0e 0f 12 1b 21 1a 20 24 1a 22 1b 1f 19 1d 20 1b 13 12 11 0d 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0b 06 07 05 06 0e 0c 0b 08 0f 1a 15 24 21 29 25 29 28 24 2e 28 2a 29 1d 23 2b 20 25 24 29 24 26 26 26 26 1f 23 25 24 26 25 27 26 2d 23 1d 2b 22 29 22 22 2c 23 21 1d 24 29 1f 1d 20 18 1b 13 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0f 1c 23 24 2d 3c 3b 36 35 37 3b 33 34 39 3a 38 39 3c 39 3d 3d 39 3b 41 44 3d 41 4a 43 49 3f 31 2b 2d 29 2a 27 28 20 2a 2b 2b 27 29 24 21 1f 1a 15 11 02 06 05 07 01 0e 06 12 16 19 1a 11 11 14 0e 06 10 09 05 11 0c 09 07 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 0c 0b 05 03 0a 0c 0e 0f 0d 1d 18 13 16 1b 18 1d 1c 15 23 19 16 0d 14 12 10 10 16 16 13 15 17 10 10 15 18 1c 1f 11 15 1a 10 0d 19 16 18 15 19 1b 1a 12 14 1c 0e 17 10 07 10 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1f 1e 33
 32 34 33 36 33 2c 34 36 37 31 2c 35 37 39 36 40 44 3f 47 42 3e 47 3b 40 38 31 2a 28 2a 19 2a 1f 1e 19 1f 26 1d 1c 12 11 17 16 0b 05 03 00 06 05 03 00 06 05 05 06 06 08 06 00 06 08 03 0a 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 10 05 05 06 11 0a 01 06 06 03 05 06 05 08 01 06 05 0c 01 06 05 03 0b 06 09 0a 09 06 07 03 05 06 0c 05 06 06 05 03 00 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 16 27 28 34 32 2e 32 2f 39 37 35 35 34 38 36 3c 43 40 3e 3c 40 40 3e 41 37 31 35 26 19 19 1e 1e 19 19 1c 22 19 1a 12 16 10 10 09 0a 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 11 26 26 2a 2a 2f 28 2c 31 32 2e 2d 25 39 31 3b 36 36 37 3a 40 37 30 33 2f 25 1f 1b 12 09 0f 0c 0e 0b 0f 0d 0d 06 00 08 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 0d 0d 16 20 20 24 25 28 21 2b 1b 27 27 2a 29 2d 25 23 28 1f 1e 20 27 16 1a 10 10 0c 03 02 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 11 0f 20 1a 12 1d 18 1b 1a 10 16 12 11 12 10 0f 14 0c 0d 10 09 08 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 07 12 06 05 07 08 06 08 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
