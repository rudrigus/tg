((X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"03", X"04", X"06", X"05", X"08", X"00", X"0a", X"06", X"05", X"0c", X"10", X"0a", X"08", X"0b", X"06", X"05", X"08", X"0f", X"0c", X"05", X"11", X"0e", X"16", X"21", X"1e", X"17", X"21", X"24", X"2d", X"36", X"36", X"45", X"49", X"4b", X"44", X"4b", X"4b", X"44", X"44", X"3f", X"40", X"44", X"3f", X"37", X"35", X"3d", X"3f", X"38", X"31", X"2f", X"34", X"24", X"2a", X"2b", X"32", X"37", X"2a", X"23", X"21", X"15", X"16", X"13", X"0f", X"10", X"0a", X"13", X"06", X"0e", X"14", X"0b", X"06", X"0b", X"0f", X"19", X"15", X"0e", X"13", X"0b", X"0b", X"10", X"03", X"05", X"0d", X"0c", X"0b", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"09", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"01", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0b", X"06", X"0a", X"0c", X"03", X"08", X"07", X"0a", X"0c", X"0d", X"07", X"15", X"0c", X"16", X"1b", X"11", X"1a", X"16", X"14", X"11", X"17", X"15", X"0f", X"16", X"15", X"15", X"14", X"1c", X"1c", X"2d", X"33", X"3a", X"3a", X"36", X"3a", X"53", X"59", X"72", X"7b", X"77", X"84", X"80", X"83", X"7b", X"78", X"71", X"76", X"74", X"75", X"7e", X"71", X"71", X"70", X"5e", X"60", X"5b", X"5f", X"50", X"4e", X"4f", X"4d", X"56", X"5b", X"50", X"4e", X"47", X"44", X"31", X"34", X"32", X"25", X"28", X"30", X"31", X"25", X"24", X"2d", X"30", X"2d", X"26", X"31", X"38", X"2d", X"1e", X"20", X"0c", X"11", X"0d", X"09", X"0f", X"14", X"12", X"15", X"0a", X"0a", X"0c", X"10", X"0d", X"05", X"04", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"0c", X"04", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"0f", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"03", X"06", X"07", X"0a", X"0a", X"11", X"10", X"08", X"0d", X"0e", X"10", X"12", X"13", X"15", X"17", X"1e", X"10", X"12", X"23", X"20", X"25", X"32", X"2f", X"32", X"25", X"2b", X"26", X"1c", X"25", X"24", X"1f", X"1f", X"26", X"30", X"42", X"4a", X"58", X"63", X"70", X"83", X"96", X"9d", X"ac", X"b6", X"be", X"c6", X"c7", X"c5", X"c1", X"ba", X"ad", X"a7", X"bc", X"c0", X"b8", X"ab", X"a2", X"91", X"94", X"97", X"94", X"86", X"7c", X"89", X"81", X"78", X"7f", X"71", X"65", X"6f", X"70", X"5e", X"53", X"3f", X"44", X"3e", X"3d", X"36", X"33", X"33", X"3b", X"3a", X"49", X"4d", X"52", X"49", X"54", X"49", X"39", X"34", X"21", X"1a", X"11", X"12", X"1b", X"11", X"13", X"06", X"05", X"06", X"0b", X"06", X"0a", X"04", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"0a", X"03", X"06", X"0b", X"03", X"00", X"06", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0d", X"0d", X"15", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"01", X"0a", X"05", X"03", X"07", X"06", X"05", X"0c", X"08", X"06", X"05", X"03", X"0f", X"18", X"14", X"10", X"16", X"10", X"1b", X"16", X"1f", X"1f", X"1d", X"2e", X"2d", X"27", X"2c", X"27", X"46", X"69", X"65", X"44", X"40", X"56", X"4b", X"41", X"3d", X"33", X"3b", X"4a", X"55", X"62", X"7a", X"87", X"96", X"a6", X"b5", X"ca", X"cc", X"dc", X"de", X"e5", X"f0", X"f9", X"fb", X"f7", X"f1", X"ea", X"e1", X"e3", X"e6", X"e0", X"da", X"d0", X"c4", X"c0", X"bf", X"c2", X"b9", X"ba", X"be", X"be", X"c7", X"c9", X"c1", X"b2", X"a2", X"9c", X"8d", X"83", X"79", X"68", X"66", X"59", X"4f", X"51", X"4e", X"40", X"42", X"41", X"4e", X"54", X"50", X"5a", X"68", X"77", X"79", X"5c", X"43", X"31", X"2a", X"1d", X"23", X"14", X"1d", X"18", X"0c", X"16", X"0f", X"06", X"0c", X"08", X"09", X"0d", X"05", X"06", X"00", X"06", X"06", X"04", X"09", X"06", X"0b", X"03", X"0f", X"07", X"0a", X"17", X"12", X"0d", X"05", X"03", X"02", X"06", X"06", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"09", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"04", X"00", X"06", X"05", X"03", X"00", X"09", X"08", X"03", X"00", X"06", X"11", X"0d", X"09", X"09", X"09", X"05", X"1d", X"1b", X"16", X"22", X"20", X"25", X"2d", X"33", X"32", X"37", X"29", X"28", X"30", X"39", X"3c", X"3e", X"55", X"6f", X"74", X"6b", X"69", X"6c", X"74", X"7f", X"80", X"76", X"77", X"91", X"92", X"95", X"a5", X"b8", X"be", X"c3", X"dd", X"e9", X"e0", X"f3", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"ee", X"f5", X"f2", X"fc", X"fa", X"fa", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"e6", X"d5", X"b4", X"a9", X"a1", X"92", X"7c", X"7d", X"77", X"7c", X"74", X"68", X"63", X"5d", X"59", X"66", X"66", X"69", X"77", X"8a", X"96", X"7d", X"74", X"54", X"4a", X"38", X"31", X"25", X"1f", X"15", X"14", X"14", X"10", X"0f", X"15", X"07", X"0e", X"09", X"05", X"03", X"04", X"06", X"07", X"05", X"05", X"06", X"09", X"0b", X"09", X"0d", X"1e", X"25", X"19", X"0d", X"05", X"03", X"03", X"06", X"06", X"05", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"0f", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"0e", X"05", X"03", X"06", X"0e", X"08", X"15", X"10", X"0c", X"14", X"1c", X"1d", X"1b", X"1b", X"19", X"1b", X"37", X"4c", X"60", X"54", X"42", X"3a", X"4a", X"44", X"53", X"55", X"68", X"76", X"7f", X"86", X"8f", X"91", X"95", X"94", X"9b", X"9e", X"96", X"a0", X"9d", X"ab", X"ba", X"c3", X"ca", X"ce", X"d5", X"d4", X"ea", X"e5", X"f4", X"fd", X"fd", X"fe", X"ff", X"ff", X"f7", X"fa", X"f3", X"ee", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"de", X"c5", X"cf", X"af", X"a1", X"9e", X"98", X"96", X"8e", X"8d", X"87", X"85", X"85", X"86", X"81", X"8c", X"9a", X"ac", X"ae", X"a3", X"9b", X"81", X"7b", X"63", X"4a", X"2c", X"2d", X"17", X"19", X"12", X"13", X"06", X"12", X"10", X"0d", X"0f", X"0a", X"0d", X"0e", X"0f", X"07", X"0b", X"04", X"0c", X"0a", X"12", X"18", X"16", X"25", X"21", X"0c", X"0f", X"06", X"09", X"02", X"07", X"08", X"08", X"0f", X"06", X"09", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0d", X"22", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"0e", X"15", X"06", X"06", X"07", X"03", X"06", X"0b", X"05", X"0e", X"0b", X"08", X"0c", X"13", X"12", X"13", X"15", X"26", X"39", X"2a", X"29", X"35", X"30", X"36", X"59", X"6c", X"65", X"5b", X"5d", X"6f", X"79", X"92", X"99", X"9c", X"95", X"93", X"8a", X"8d", X"9e", X"a1", X"9a", X"a6", X"9c", X"ab", X"a4", X"a1", X"a9", X"af", X"c1", X"c0", X"cb", X"cc", X"c2", X"d2", X"e2", X"e9", X"ec", X"e3", X"f0", X"f2", X"f7", X"f2", X"f3", X"ed", X"f2", X"ee", X"ee", X"e7", X"eb", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"ef", X"d7", X"c2", X"b6", X"ad", X"a4", X"a9", X"ac", X"9c", X"a6", X"a1", X"99", X"97", X"9d", X"ae", X"b2", X"bf", X"c2", X"c0", X"b2", X"a4", X"8d", X"73", X"53", X"36", X"29", X"1a", X"22", X"1d", X"24", X"1d", X"10", X"07", X"13", X"0f", X"0a", X"0e", X"11", X"0f", X"0a", X"0b", X"13", X"15", X"25", X"30", X"35", X"28", X"23", X"1a", X"07", X"0c", X"0d", X"0b", X"0d", X"05", X"06", X"0a", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"15", X"24", X"20", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"0d", X"03", X"09", X"06", X"0a", X"0e", X"09", X"07", X"0d", X"0d", X"0c", X"19", X"17", X"1c", X"1d", X"17", X"2c", X"30", X"32", X"2f", X"3f", X"48", X"49", X"5e", X"80", X"88", X"93", X"a6", X"ae", X"c6", X"cb", X"c3", X"b1", X"a2", X"90", X"82", X"7e", X"87", X"9d", X"a0", X"a9", X"ae", X"b5", X"b2", X"b4", X"b9", X"ac", X"bf", X"c9", X"cf", X"d7", X"dc", X"d0", X"df", X"ee", X"f2", X"fb", X"f3", X"f7", X"f2", X"f7", X"f6", X"f4", X"f5", X"ef", X"e4", X"d9", X"d1", X"c5", X"c1", X"cd", X"cf", X"e4", X"f3", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"d8", X"cc", X"be", X"b4", X"b6", X"b8", X"ad", X"ab", X"a8", X"a7", X"a1", X"a6", X"b2", X"b6", X"bb", X"be", X"c2", X"bb", X"bf", X"b7", X"aa", X"87", X"62", X"3e", X"2d", X"28", X"2a", X"25", X"25", X"28", X"1e", X"1d", X"1e", X"18", X"16", X"18", X"14", X"12", X"11", X"1b", X"1b", X"29", X"30", X"36", X"3d", X"3e", X"2a", X"27", X"1c", X"15", X"0f", X"06", X"05", X"10", X"07", X"07", X"0d", X"03", X"04", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"0e", X"2a", X"29", X"18", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"05", X"06", X"06", X"05", X"0a", X"04", X"09", X"0e", X"0b", X"0f", X"0e", X"0c", X"16", X"16", X"17", X"19", X"21", X"25", X"2e", X"32", X"2b", X"3c", X"44", X"4c", X"5d", X"7e", X"98", X"af", X"c9", X"de", X"eb", X"f1", X"e5", X"cd", X"b8", X"9b", X"8e", X"7b", X"76", X"89", X"7f", X"93", X"a2", X"b4", X"b5", X"c6", X"ca", X"c3", X"c0", X"bd", X"cf", X"dc", X"de", X"dd", X"ea", X"e3", X"f4", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"f0", X"e1", X"da", X"d4", X"c5", X"b5", X"b7", X"b4", X"b0", X"bb", X"c6", X"c1", X"be", X"c5", X"c4", X"bc", X"c6", X"c4", X"cb", X"d6", X"db", X"e2", X"f5", X"f0", X"e0", X"ca", X"c7", X"b9", X"b1", X"c6", X"b7", X"b0", X"b4", X"aa", X"af", X"bf", X"c4", X"c2", X"bc", X"c6", X"c7", X"d2", X"c9", X"c1", X"c3", X"ae", X"94", X"77", X"5d", X"4c", X"46", X"3b", X"38", X"32", X"2f", X"26", X"24", X"20", X"19", X"24", X"19", X"16", X"1f", X"20", X"34", X"40", X"48", X"65", X"5d", X"54", X"4f", X"55", X"53", X"3b", X"16", X"0d", X"12", X"0a", X"0b", X"0b", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0d", X"2a", X"37", X"25", X"0b", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"04", X"0c", X"06", X"0a", X"07", X"08", X"07", X"05", X"0a", X"04", X"06", X"05", X"0a", X"1b", X"11", X"0b", X"12", X"1b", X"16", X"15", X"23", X"1f", X"2c", X"2b", X"36", X"3c", X"3b", X"41", X"45", X"55", X"63", X"88", X"a5", X"c2", X"d1", X"e0", X"e4", X"fe", X"ff", X"eb", X"d9", X"bd", X"9c", X"87", X"7e", X"81", X"7d", X"87", X"94", X"9b", X"ae", X"c5", X"cb", X"cf", X"d4", X"d5", X"d8", X"dc", X"e2", X"f4", X"fa", X"f2", X"fe", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f3", X"e3", X"dd", X"c6", X"be", X"b5", X"b1", X"b7", X"ae", X"b8", X"b1", X"ae", X"b4", X"aa", X"ab", X"aa", X"b0", X"ae", X"b3", X"b4", X"b9", X"cf", X"d6", X"ce", X"c3", X"bd", X"b9", X"af", X"b8", X"b1", X"ad", X"b4", X"ac", X"a7", X"be", X"ca", X"c2", X"bf", X"bb", X"ca", X"d5", X"d9", X"dc", X"cf", X"c9", X"c2", X"b6", X"96", X"7d", X"7e", X"64", X"5f", X"51", X"51", X"49", X"32", X"37", X"34", X"2b", X"31", X"32", X"34", X"3b", X"62", X"6a", X"87", X"98", X"a3", X"a2", X"95", X"a1", X"8b", X"5e", X"3c", X"1b", X"1b", X"1c", X"1d", X"22", X"0d", X"03", X"06", X"07", X"0a", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"16", X"30", X"2d", X"21", X"0a", X"01", X"06", X"05", X"05", X"00", X"06", X"08", X"09", X"06", X"06", X"0d", X"0c", X"16", X"20", X"0d", X"0f", X"11", X"12", X"14", X"17", X"18", X"1d", X"1d", X"1e", X"21", X"28", X"25", X"26", X"33", X"2f", X"42", X"42", X"4d", X"53", X"54", X"67", X"7f", X"9d", X"b5", X"cf", X"dc", X"e4", X"e5", X"f1", X"fd", X"e6", X"de", X"c7", X"ab", X"93", X"96", X"93", X"8d", X"8f", X"8e", X"9c", X"a4", X"ad", X"c4", X"cb", X"d5", X"da", X"da", X"e8", X"e6", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"ee", X"df", X"ca", X"c4", X"c3", X"b8", X"b9", X"bb", X"b4", X"af", X"b3", X"b6", X"b3", X"af", X"a9", X"b2", X"a9", X"a6", X"b3", X"b5", X"b9", X"bc", X"b8", X"ac", X"b3", X"b7", X"af", X"ac", X"ad", X"a4", X"ae", X"ae", X"af", X"b4", X"bf", X"bf", X"b6", X"ba", X"c1", X"d7", X"e0", X"e6", X"e4", X"dc", X"db", X"d5", X"c0", X"b1", X"b0", X"a0", X"9d", X"88", X"79", X"6a", X"5f", X"58", X"5d", X"5d", X"5b", X"61", X"59", X"7d", X"87", X"a0", X"b0", X"c7", X"c5", X"ce", X"c6", X"ac", X"91", X"73", X"55", X"4b", X"46", X"37", X"35", X"29", X"13", X"11", X"0d", X"0d", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"11", X"17", X"23", X"21", X"08", X"03", X"00", X"06", X"05", X"03", X"08", X"0a", X"05", X"0d", X"0d", X"0b", X"1c", X"25", X"25", X"2f", X"2c", X"1d", X"1f", X"20", X"24", X"28", X"25", X"24", X"25", X"33", X"36", X"38", X"3d", X"3f", X"46", X"47", X"52", X"53", X"5e", X"78", X"85", X"97", X"a4", X"c6", X"d6", X"e2", X"eb", X"e7", X"f2", X"fc", X"f1", X"e7", X"d2", X"b7", X"aa", X"a1", X"9c", X"a7", X"a0", X"9d", X"92", X"a7", X"b3", X"b5", X"c7", X"d9", X"d8", X"dd", X"e3", X"e7", X"ee", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ea", X"d4", X"dd", X"d2", X"d0", X"ce", X"c4", X"c4", X"bc", X"b8", X"b8", X"b9", X"ae", X"af", X"b0", X"ad", X"a8", X"b6", X"b5", X"b7", X"be", X"b3", X"b9", X"ab", X"b0", X"af", X"a9", X"a3", X"a0", X"a4", X"aa", X"a6", X"a9", X"ab", X"a8", X"af", X"b0", X"b9", X"c4", X"ca", X"d9", X"e7", X"ea", X"ef", X"ed", X"e0", X"e4", X"da", X"d6", X"ca", X"b7", X"af", X"96", X"8d", X"8c", X"91", X"8f", X"87", X"86", X"8b", X"8c", X"8c", X"99", X"a0", X"ac", X"bb", X"bc", X"b3", X"b6", X"a3", X"89", X"71", X"61", X"59", X"51", X"46", X"3b", X"29", X"31", X"1f", X"1a", X"0d", X"11", X"09", X"09", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"07", X"12", X"18", X"14", X"05", X"03", X"04", X"06", X"11", X"0e", X"18", X"1b", X"1e", X"1f", X"25", X"2a", X"2e", X"34", X"3b", X"3d", X"37", X"2f", X"2e", X"25", X"34", X"37", X"39", X"3f", X"38", X"3c", X"38", X"40", X"46", X"51", X"5f", X"6d", X"74", X"7c", X"86", X"9c", X"a3", X"ac", X"bf", X"d3", X"e9", X"f3", X"f1", X"fa", X"ff", X"ff", X"f5", X"e5", X"c8", X"b7", X"b7", X"b3", X"bc", X"b0", X"b1", X"b0", X"a8", X"b5", X"be", X"c7", X"d3", X"dd", X"e4", X"ea", X"e6", X"f5", X"f2", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f0", X"e6", X"e0", X"d5", X"d6", X"d4", X"d2", X"c9", X"cd", X"c7", X"c2", X"b9", X"ba", X"b4", X"b9", X"b7", X"b3", X"b2", X"c1", X"bb", X"bf", X"b6", X"b9", X"a7", X"b1", X"ae", X"ae", X"af", X"a5", X"ae", X"a6", X"ad", X"9f", X"a9", X"a8", X"a8", X"b0", X"bb", X"cb", X"c8", X"db", X"e8", X"eb", X"f6", X"fc", X"f6", X"ff", X"f3", X"f7", X"e5", X"d5", X"c1", X"b1", X"a1", X"93", X"92", X"92", X"90", X"91", X"99", X"94", X"95", X"a2", X"a1", X"aa", X"ad", X"ac", X"ac", X"a6", X"94", X"86", X"77", X"77", X"5e", X"4c", X"4a", X"4d", X"47", X"43", X"3a", X"24", X"21", X"13", X"11", X"08", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0f", X"0d", X"11", X"06", X"08", X"05", X"0c", X"0c", X"17", X"20", X"25", X"29", X"2d", X"28", X"32", X"3f", X"35", X"41", X"44", X"41", X"37", X"32", X"3c", X"37", X"45", X"4c", X"4f", X"50", X"50", X"51", X"4d", X"58", X"5f", X"6b", X"77", X"85", X"8c", X"94", X"99", X"a7", X"ad", X"bc", X"d2", X"e0", X"ef", X"fb", X"fe", X"ff", X"ff", X"ff", X"fb", X"e5", X"d8", X"c9", X"ce", X"ca", X"c2", X"c4", X"b5", X"bd", X"bf", X"c9", X"ce", X"db", X"e5", X"ef", X"f8", X"f6", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f1", X"e3", X"e4", X"e4", X"e6", X"da", X"d3", X"d3", X"d8", X"c0", X"c9", X"be", X"c1", X"c6", X"b5", X"b8", X"be", X"c1", X"c0", X"c4", X"c3", X"b6", X"ba", X"b1", X"b4", X"bb", X"b0", X"b3", X"b2", X"b1", X"b1", X"af", X"a9", X"ae", X"ab", X"b1", X"bf", X"c1", X"cb", X"cd", X"d1", X"e4", X"ec", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f0", X"d7", X"c7", X"b7", X"9f", X"a1", X"9b", X"97", X"99", X"a3", X"9d", X"99", X"a9", X"b5", X"b7", X"bb", X"b3", X"a7", X"9b", X"97", X"83", X"74", X"7d", X"66", X"5f", X"61", X"5c", X"62", X"56", X"55", X"4d", X"2c", X"26", X"12", X"06", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"14", X"11", X"04", X"06", X"05", X"12", X"18", X"12", X"1b", X"1c", X"25", X"2b", X"39", X"38", X"43", X"44", X"45", X"43", X"4a", X"42", X"43", X"45", X"4c", X"49", X"4d", X"52", X"52", X"59", X"5b", X"6b", X"6c", X"65", X"71", X"77", X"85", X"99", X"a0", X"a9", X"af", X"b6", X"c3", X"cc", X"d3", X"e4", X"f2", X"ff", X"ff", X"ff", X"ff", X"fd", X"f2", X"eb", X"e2", X"e1", X"dd", X"db", X"d8", X"cd", X"cd", X"ca", X"d4", X"df", X"e3", X"e5", X"ea", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"f3", X"f8", X"ef", X"eb", X"e2", X"db", X"d9", X"d2", X"d5", X"c4", X"ca", X"ca", X"c4", X"ca", X"bd", X"c4", X"c4", X"c3", X"cc", X"cb", X"c6", X"c4", X"c1", X"c3", X"ba", X"bc", X"bb", X"bb", X"b3", X"b8", X"b1", X"b9", X"c1", X"b9", X"bc", X"c1", X"c3", X"cc", X"d3", X"ca", X"d4", X"e5", X"e7", X"f3", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"f1", X"ea", X"d5", X"c2", X"b8", X"b1", X"a5", X"ae", X"b1", X"a7", X"ae", X"c3", X"b7", X"be", X"b6", X"aa", X"9f", X"94", X"91", X"89", X"83", X"80", X"7d", X"70", X"6f", X"6f", X"61", X"64", X"60", X"52", X"3c", X"2c", X"19", X"09", X"09", X"05", X"03", X"0b", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"0a", X"17", X"07", X"0b", X"0e", X"0c", X"10", X"20", X"1b", X"24", X"25", X"2c", X"2d", X"34", X"3f", X"40", X"45", X"53", X"55", X"54", X"49", X"50", X"5a", X"58", X"59", X"53", X"56", X"5c", X"6c", X"64", X"6b", X"6c", X"6d", X"78", X"88", X"a0", X"ae", X"bb", X"d2", X"d2", X"db", X"e4", X"e6", X"e0", X"f3", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"ff", X"ff", X"ff", X"fb", X"e8", X"e7", X"e8", X"ef", X"ef", X"fa", X"ef", X"ef", X"fa", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f7", X"f7", X"f6", X"f3", X"e5", X"eb", X"e4", X"da", X"d6", X"d1", X"d1", X"d2", X"cd", X"d1", X"be", X"cc", X"ce", X"cf", X"d8", X"d4", X"ca", X"c9", X"c7", X"cc", X"c6", X"bd", X"cb", X"c7", X"c4", X"c5", X"c4", X"bd", X"c2", X"c7", X"c5", X"ca", X"c1", X"c7", X"ce", X"d4", X"c8", X"cd", X"d0", X"d3", X"e1", X"df", X"fb", X"ff", X"fd", X"ff", X"fc", X"f8", X"f1", X"dc", X"d4", X"c0", X"b6", X"c1", X"c9", X"bd", X"c7", X"c6", X"d0", X"c4", X"b6", X"9e", X"98", X"94", X"95", X"90", X"90", X"91", X"8b", X"7e", X"82", X"71", X"69", X"62", X"51", X"3d", X"38", X"2d", X"1a", X"18", X"0f", X"0b", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"17", X"1b", X"12", X"14", X"10", X"0f", X"1b", X"1d", X"1b", X"18", X"24", X"2d", X"30", X"3e", X"41", X"3e", X"51", X"55", X"65", X"5a", X"5e", X"5d", X"54", X"57", X"5e", X"51", X"54", X"55", X"59", X"64", X"67", X"6a", X"60", X"71", X"84", X"9d", X"c5", X"cc", X"e5", X"ef", X"f9", X"f4", X"ff", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f1", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"fc", X"f3", X"fa", X"ee", X"ec", X"ed", X"e3", X"db", X"dc", X"de", X"d1", X"d4", X"d2", X"ce", X"d6", X"d2", X"d7", X"d6", X"d3", X"d3", X"df", X"d3", X"d3", X"d1", X"d1", X"ca", X"cd", X"cf", X"c7", X"cf", X"c9", X"cd", X"c6", X"d1", X"cc", X"c9", X"cf", X"cf", X"c6", X"cc", X"c5", X"c6", X"cd", X"c8", X"d0", X"db", X"e6", X"f4", X"ff", X"f9", X"f8", X"ec", X"ea", X"dc", X"d2", X"d7", X"d5", X"de", X"dd", X"dd", X"cf", X"c8", X"c3", X"aa", X"99", X"92", X"9b", X"9a", X"96", X"9b", X"92", X"84", X"92", X"87", X"74", X"69", X"50", X"35", X"34", X"29", X"25", X"23", X"21", X"14", X"0c", X"0e", X"10", X"06", X"07", X"03", X"00", X"06", X"09", X"05", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"0d", X"0a", X"17", X"10", X"09", X"10", X"11", X"08", X"0f", X"1c", X"20", X"2a", X"25", X"2f", X"35", X"32", X"48", X"48", X"54", X"67", X"63", X"66", X"60", X"60", X"5e", X"54", X"52", X"51", X"55", X"50", X"4e", X"50", X"67", X"67", X"64", X"76", X"84", X"9f", X"ba", X"d1", X"ee", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f5", X"fd", X"fb", X"f3", X"f4", X"ed", X"ee", X"e2", X"e4", X"d9", X"d7", X"d8", X"d5", X"d6", X"d6", X"da", X"d9", X"d9", X"da", X"d9", X"e3", X"e1", X"de", X"d6", X"da", X"d3", X"d5", X"d4", X"d1", X"ce", X"d7", X"d1", X"d6", X"d2", X"d2", X"c9", X"ce", X"c9", X"cb", X"cf", X"c9", X"c4", X"c9", X"cb", X"cc", X"d2", X"cf", X"e5", X"f1", X"fa", X"f1", X"f1", X"e8", X"d8", X"df", X"da", X"e3", X"ec", X"e7", X"dc", X"d9", X"c0", X"a9", X"9d", X"a0", X"a2", X"9e", X"9e", X"a1", X"a4", X"a7", X"9b", X"9f", X"94", X"8c", X"7b", X"57", X"48", X"35", X"2b", X"31", X"28", X"29", X"20", X"1b", X"16", X"14", X"09", X"09", X"03", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"0f", X"10", X"13", X"14", X"0d", X"1c", X"17", X"1e", X"20", X"2b", X"2d", X"32", X"36", X"3b", X"3e", X"48", X"55", X"5e", X"64", X"68", X"69", X"6e", X"63", X"65", X"60", X"61", X"5b", X"50", X"54", X"51", X"5c", X"5f", X"65", X"5d", X"69", X"80", X"9e", X"c2", X"d7", X"ed", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"f7", X"f3", X"e9", X"ef", X"ec", X"e2", X"e5", X"e0", X"df", X"da", X"de", X"d6", X"e0", X"e1", X"e0", X"e0", X"ea", X"e3", X"e4", X"e5", X"e1", X"e6", X"da", X"e6", X"d8", X"e2", X"dc", X"d2", X"d9", X"d1", X"d7", X"db", X"d6", X"d0", X"ce", X"d5", X"d5", X"ce", X"cc", X"cf", X"c6", X"ca", X"d0", X"d5", X"d6", X"ea", X"e8", X"e1", X"ea", X"d5", X"e1", X"db", X"e6", X"e4", X"ef", X"de", X"da", X"cc", X"bc", X"a8", X"9e", X"99", X"a3", X"a6", X"ab", X"af", X"b1", X"b2", X"ae", X"b0", X"a5", X"98", X"8b", X"7c", X"5d", X"4c", X"49", X"41", X"35", X"2f", X"23", X"18", X"12", X"15", X"16", X"14", X"12", X"0d", X"07", X"07", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"08", X"06", X"07", X"07", X"10", X"0f", X"0d", X"15", X"12", X"13", X"19", X"20", X"1f", X"2e", X"31", X"3c", X"46", X"4b", X"4a", X"53", X"4d", X"5d", X"5b", X"64", X"66", X"6a", X"69", X"65", X"66", X"6b", X"70", X"6d", X"67", X"63", X"62", X"62", X"64", X"64", X"6d", X"71", X"7f", X"94", X"b1", X"c6", X"e1", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"fe", X"f5", X"f7", X"ed", X"f3", X"f5", X"ed", X"ec", X"e7", X"e3", X"e5", X"e6", X"e6", X"e7", X"e9", X"ef", X"e5", X"ee", X"ea", X"e9", X"e7", X"ec", X"f2", X"ea", X"e8", X"e4", X"de", X"dd", X"d8", X"dd", X"de", X"da", X"d5", X"d5", X"d5", X"cf", X"d5", X"dc", X"d3", X"d3", X"cd", X"d0", X"d6", X"dc", X"dd", X"da", X"e4", X"d4", X"de", X"d5", X"d1", X"d4", X"d7", X"db", X"d9", X"dd", X"d3", X"c6", X"aa", X"9b", X"a2", X"a5", X"a6", X"b1", X"b7", X"be", X"c2", X"cd", X"bd", X"c0", X"c5", X"b2", X"a9", X"93", X"7e", X"70", X"63", X"52", X"46", X"2e", X"35", X"25", X"1c", X"1f", X"1d", X"15", X"1d", X"10", X"07", X"0c", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"01", X"06", X"0c", X"05", X"0e", X"0b", X"0c", X"16", X"21", X"22", X"2e", X"36", X"32", X"41", X"3f", X"4b", X"4a", X"4f", X"4f", X"5a", X"59", X"60", X"65", X"6e", X"6f", X"6d", X"62", X"66", X"6b", X"7c", X"76", X"74", X"62", X"62", X"66", X"64", X"6b", X"71", X"7f", X"8a", X"9c", X"ab", X"c9", X"e6", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"fe", X"fd", X"fa", X"fb", X"f5", X"f4", X"f1", X"e7", X"e9", X"e5", X"e8", X"ed", X"e7", X"e7", X"f0", X"eb", X"ef", X"f4", X"ee", X"f6", X"f5", X"f8", X"f9", X"ef", X"eb", X"e7", X"e6", X"e3", X"d7", X"e1", X"d7", X"d8", X"d8", X"d2", X"d8", X"d1", X"de", X"d4", X"d5", X"d3", X"de", X"e1", X"d6", X"e2", X"e0", X"e1", X"dc", X"db", X"cf", X"ce", X"cc", X"d3", X"cd", X"d0", X"c9", X"b9", X"b7", X"a3", X"9f", X"a6", X"a4", X"aa", X"b8", X"c1", X"cc", X"d3", X"d1", X"d3", X"cf", X"d1", X"c7", X"b1", X"a3", X"94", X"85", X"74", X"6c", X"63", X"5d", X"45", X"35", X"36", X"27", X"19", X"1b", X"11", X"17", X"06", X"08", X"06", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"09", X"03", X"04", X"0a", X"0f", X"11", X"0f", X"11", X"14", X"16", X"28", X"33", X"45", X"42", X"49", X"4b", X"4b", X"4c", X"50", X"4e", X"4e", X"52", X"63", X"64", X"66", X"65", X"70", X"73", X"73", X"75", X"77", X"78", X"7e", X"7e", X"71", X"76", X"79", X"77", X"7a", X"82", X"8d", X"9e", X"a9", X"a5", X"bc", X"ce", X"e0", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"f8", X"fd", X"fb", X"fd", X"f9", X"f4", X"f2", X"ef", X"eb", X"e8", X"ef", X"ed", X"ee", X"ec", X"f3", X"f5", X"f7", X"f5", X"fc", X"ff", X"fe", X"ff", X"ff", X"fb", X"ee", X"ec", X"e5", X"eb", X"e5", X"e6", X"e2", X"e1", X"e4", X"e2", X"e2", X"e0", X"e3", X"e4", X"e2", X"e6", X"e4", X"ed", X"ef", X"e7", X"e4", X"dd", X"e0", X"d8", X"d3", X"d4", X"ce", X"cb", X"c8", X"c6", X"c0", X"ae", X"a6", X"9a", X"9a", X"a2", X"ab", X"b0", X"b8", X"cb", X"d7", X"cf", X"de", X"e1", X"e0", X"e2", X"de", X"ca", X"b6", X"a0", X"9c", X"85", X"81", X"72", X"71", X"68", X"5c", X"4d", X"40", X"2b", X"1d", X"20", X"1e", X"15", X"10", X"0b", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"0a", X"06", X"05", X"0c", X"0d", X"16", X"17", X"1d", X"15", X"12", X"17", X"20", X"2f", X"41", X"43", X"45", X"42", X"49", X"4b", X"4c", X"51", X"50", X"55", X"55", X"5c", X"62", X"72", X"74", X"7b", X"79", X"74", X"78", X"77", X"81", X"8e", X"88", X"81", X"7f", X"7d", X"7d", X"8a", X"93", X"a5", X"bb", X"bc", X"b8", X"b7", X"c8", X"d8", X"e6", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fc", X"f9", X"f5", X"f9", X"f9", X"f3", X"f1", X"fa", X"f5", X"f5", X"fc", X"fd", X"f7", X"fe", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f7", X"f1", X"fa", X"f2", X"ea", X"f0", X"e9", X"e5", X"e9", X"ef", X"f6", X"f0", X"f1", X"f5", X"f0", X"f7", X"ff", X"fb", X"fd", X"f4", X"f1", X"ea", X"e3", X"d7", X"d0", X"d3", X"cd", X"ca", X"c5", X"bd", X"a7", X"9d", X"9e", X"a9", X"a7", X"b3", X"c1", X"d3", X"dd", X"de", X"dc", X"e4", X"e4", X"ee", X"ec", X"dd", X"d3", X"b5", X"b4", X"a6", X"99", X"94", X"8f", X"7f", X"74", X"6e", X"59", X"61", X"42", X"27", X"1a", X"20", X"12", X"07", X"0a", X"09", X"10", X"05", X"0a", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"0a", X"05", X"06", X"06", X"0d", X"16", X"1a", X"1e", X"1a", X"16", X"19", X"15", X"1e", X"28", X"3a", X"40", X"4a", X"42", X"41", X"4d", X"40", X"51", X"54", X"4f", X"60", X"5e", X"5e", X"67", X"6e", X"71", X"79", X"75", X"72", X"7e", X"7e", X"8e", X"91", X"8d", X"92", X"89", X"90", X"88", X"9a", X"ad", X"c1", X"c3", X"bb", X"b4", X"bb", X"c0", X"cf", X"e2", X"e4", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fd", X"ff", X"fd", X"ff", X"ff", X"fe", X"fe", X"ff", X"f8", X"f5", X"f2", X"f1", X"fe", X"fc", X"ff", X"fd", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"f2", X"f4", X"f9", X"f9", X"f1", X"ee", X"f3", X"f8", X"fb", X"fc", X"ff", X"f7", X"fc", X"ff", X"ff", X"ff", X"fd", X"fc", X"e9", X"ec", X"e5", X"de", X"d5", X"dd", X"c9", X"cf", X"be", X"b5", X"ae", X"a8", X"af", X"a7", X"bc", X"c7", X"da", X"e5", X"e8", X"ec", X"e0", X"e7", X"ee", X"eb", X"e5", X"dd", X"d5", X"bc", X"b7", X"a7", X"97", X"9b", X"8f", X"87", X"77", X"6d", X"6d", X"5c", X"4f", X"37", X"2a", X"0b", X"13", X"09", X"06", X"0a", X"0f", X"1a", X"0b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"02", X"09", X"05", X"07", X"0c", X"0d", X"13", X"15", X"1f", X"29", X"17", X"22", X"28", X"29", X"3f", X"49", X"4c", X"45", X"4a", X"4b", X"4a", X"3f", X"4f", X"50", X"58", X"61", X"63", X"62", X"66", X"6c", X"6a", X"6c", X"7a", X"77", X"81", X"85", X"86", X"8d", X"8f", X"91", X"95", X"95", X"a2", X"a8", X"b1", X"bd", X"cb", X"ca", X"c6", X"c0", X"c0", X"c7", X"cd", X"cb", X"de", X"ee", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"ff", X"fc", X"ff", X"ff", X"ff", X"ff", X"f9", X"ff", X"fb", X"ff", X"fb", X"f3", X"fa", X"fb", X"ff", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"ff", X"fb", X"f9", X"f1", X"ed", X"f8", X"f6", X"fc", X"fe", X"fa", X"ff", X"fe", X"fd", X"ff", X"ff", X"ff", X"f6", X"ed", X"f0", X"f1", X"e9", X"e7", X"e9", X"e8", X"db", X"db", X"cd", X"b4", X"b9", X"b5", X"b5", X"c4", X"ca", X"dc", X"e8", X"e6", X"e5", X"e6", X"ea", X"ee", X"ea", X"e2", X"e5", X"dc", X"db", X"ca", X"b7", X"a1", X"96", X"99", X"98", X"90", X"80", X"7f", X"7b", X"6c", X"6e", X"52", X"3a", X"21", X"10", X"06", X"04", X"09", X"0e", X"0e", X"10", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"06", X"0a", X"05", X"05", X"19", X"15", X"15", X"19", X"1c", X"30", X"3c", X"41", X"43", X"5a", X"63", X"6d", X"6b", X"5e", X"59", X"57", X"44", X"4e", X"53", X"54", X"5e", X"64", X"64", X"73", X"73", X"70", X"80", X"83", X"8b", X"8b", X"89", X"94", X"9d", X"97", X"9f", X"aa", X"a9", X"b4", X"c3", X"bf", X"ce", X"d4", X"d6", X"d4", X"cf", X"c9", X"ce", X"cf", X"c9", X"cf", X"d5", X"dd", X"e1", X"ee", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"fb", X"fe", X"fe", X"ff", X"fe", X"f9", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f4", X"f5", X"ef", X"ed", X"ed", X"eb", X"e6", X"e1", X"ba", X"d4", X"ca", X"cf", X"d1", X"d2", X"dd", X"e5", X"f3", X"f8", X"ec", X"e6", X"ec", X"eb", X"e1", X"e1", X"e5", X"dc", X"e4", X"d5", X"c8", X"bf", X"ae", X"9c", X"9f", X"9f", X"9a", X"93", X"7c", X"77", X"77", X"77", X"69", X"59", X"3c", X"1a", X"0e", X"0d", X"11", X"0b", X"14", X"1b", X"17", X"08", X"04", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"0b", X"05", X"09", X"01", X"06", X"11", X"15", X"1d", X"17", X"0d", X"18", X"27", X"3d", X"4a", X"50", X"58", X"72", X"85", X"8a", X"87", X"7d", X"72", X"55", X"50", X"57", X"5b", X"65", X"6e", X"72", X"78", X"7c", X"84", X"8e", X"94", X"9b", X"9c", X"a3", X"a3", X"aa", X"a6", X"ad", X"b0", X"ba", X"c4", X"d2", X"e8", X"da", X"d4", X"cd", X"ca", X"db", X"cc", X"d5", X"cc", X"cd", X"d6", X"d1", X"d5", X"d6", X"e0", X"df", X"ec", X"f1", X"eb", X"f2", X"f5", X"f7", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fe", X"f9", X"ff", X"fd", X"fd", X"f9", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f8", X"fa", X"fa", X"f5", X"f4", X"fd", X"ed", X"e7", X"f1", X"e1", X"e8", X"e5", X"e4", X"e7", X"f4", X"f8", X"ff", X"ff", X"f4", X"f1", X"eb", X"dd", X"d6", X"df", X"d4", X"d4", X"d7", X"cd", X"c8", X"b5", X"b0", X"a0", X"9c", X"9f", X"9f", X"95", X"88", X"7e", X"76", X"70", X"69", X"5a", X"4b", X"26", X"1b", X"12", X"07", X"0c", X"0e", X"0e", X"0f", X"11", X"03", X"00", X"06", X"05", X"09", X"00", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"06", X"06", X"10", X"0c", X"12", X"13", X"06", X"17", X"23", X"2f", X"46", X"63", X"6f", X"71", X"7e", X"83", X"91", X"8d", X"7b", X"72", X"6e", X"6a", X"6d", X"72", X"7f", X"82", X"86", X"99", X"99", X"a0", X"ad", X"b6", X"c5", X"c9", X"bc", X"ce", X"c0", X"ca", X"ce", X"d4", X"d2", X"d7", X"e9", X"e7", X"dd", X"cf", X"d6", X"d5", X"d3", X"cf", X"d6", X"d6", X"d9", X"d6", X"db", X"d9", X"dc", X"dd", X"e3", X"e3", X"e0", X"e6", X"e0", X"ea", X"f0", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"ff", X"ff", X"fc", X"fd", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"fb", X"fd", X"ff", X"fe", X"ff", X"ff", X"f6", X"fe", X"f7", X"f5", X"f7", X"f6", X"fc", X"fb", X"ff", X"fa", X"f4", X"ef", X"ec", X"e0", X"db", X"da", X"de", X"d1", X"ce", X"c7", X"bf", X"bd", X"c5", X"b2", X"a6", X"9c", X"9b", X"99", X"8e", X"73", X"6f", X"6b", X"6f", X"64", X"5b", X"53", X"42", X"2f", X"20", X"11", X"0e", X"0c", X"0a", X"14", X"0c", X"0e", X"00", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"0b", X"0c", X"0c", X"06", X"0c", X"0f", X"13", X"10", X"1b", X"2f", X"46", X"59", X"6d", X"7c", X"85", X"87", X"8e", X"93", X"8a", X"7d", X"7b", X"77", X"78", X"83", X"83", X"86", X"97", X"9a", X"9b", X"a5", X"b0", X"ba", X"cd", X"d5", X"e0", X"db", X"de", X"dd", X"e3", X"e9", X"e8", X"ea", X"e3", X"df", X"e5", X"d8", X"d8", X"d5", X"da", X"db", X"d6", X"da", X"de", X"e1", X"e9", X"e4", X"dd", X"e5", X"e4", X"e6", X"e8", X"e2", X"e5", X"ed", X"ec", X"f9", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f4", X"ec", X"e6", X"e0", X"dc", X"cf", X"d3", X"cd", X"c6", X"cd", X"c0", X"bd", X"bd", X"a8", X"a2", X"99", X"8c", X"87", X"7d", X"65", X"66", X"5e", X"54", X"48", X"51", X"4b", X"3f", X"3d", X"29", X"23", X"12", X"10", X"0d", X"0c", X"09", X"0a", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"0a", X"06", X"05", X"09", X"03", X"0a", X"0d", X"18", X"19", X"20", X"28", X"38", X"5f", X"81", X"72", X"7b", X"88", X"80", X"8a", X"8d", X"86", X"81", X"7e", X"7e", X"77", X"82", X"8e", X"95", X"9c", X"9e", X"a8", X"b0", X"ba", X"bd", X"da", X"db", X"e5", X"ea", X"ec", X"ec", X"ed", X"f1", X"e5", X"e6", X"dc", X"e1", X"d4", X"db", X"de", X"e0", X"d4", X"e6", X"de", X"e3", X"ed", X"e8", X"e7", X"ed", X"f1", X"ed", X"e7", X"f0", X"eb", X"f1", X"f4", X"f5", X"f4", X"f1", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"fd", X"f6", X"e6", X"de", X"da", X"d6", X"da", X"cd", X"c2", X"be", X"ba", X"b9", X"ae", X"b2", X"ac", X"a1", X"92", X"8d", X"7b", X"72", X"6d", X"5b", X"58", X"56", X"4f", X"44", X"43", X"48", X"49", X"37", X"33", X"1c", X"12", X"06", X"0b", X"0d", X"0c", X"0c", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"04", X"0a", X"0d", X"15", X"0f", X"1a", X"17", X"31", X"5a", X"85", X"9e", X"8c", X"84", X"87", X"7d", X"84", X"80", X"7b", X"75", X"82", X"86", X"87", X"8b", X"8d", X"98", X"9b", X"a3", X"a8", X"af", X"b8", X"c8", X"cc", X"cf", X"e0", X"e9", X"e9", X"ed", X"eb", X"e6", X"e4", X"d7", X"df", X"d4", X"d6", X"e0", X"d3", X"e0", X"db", X"de", X"e1", X"e3", X"e5", X"ea", X"ea", X"ef", X"f5", X"f3", X"f3", X"f1", X"f7", X"f0", X"f5", X"fa", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f6", X"fb", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f8", X"ea", X"e5", X"db", X"e1", X"d1", X"d1", X"c6", X"c1", X"b5", X"b2", X"b1", X"ad", X"a3", X"a5", X"9f", X"94", X"89", X"7d", X"6a", X"6a", X"5a", X"5e", X"53", X"4c", X"51", X"4b", X"44", X"48", X"41", X"36", X"25", X"17", X"14", X"06", X"07", X"10", X"12", X"0f", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"0a", X"07", X"05", X"0c", X"10", X"09", X"06", X"14", X"17", X"1d", X"3e", X"64", X"97", X"b5", X"91", X"79", X"7f", X"7f", X"84", X"85", X"81", X"85", X"84", X"7c", X"8b", X"87", X"8c", X"90", X"92", X"a5", X"b1", X"b5", X"ba", X"c2", X"c9", X"ce", X"d6", X"e2", X"de", X"e9", X"d9", X"da", X"d3", X"df", X"da", X"df", X"d4", X"dd", X"dd", X"e4", X"e4", X"e7", X"e8", X"e3", X"f0", X"ec", X"f1", X"f7", X"fc", X"ff", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"fc", X"ff", X"fb", X"ff", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f3", X"f0", X"e8", X"e3", X"e6", X"d5", X"cb", X"c9", X"b6", X"b6", X"bd", X"b4", X"af", X"a2", X"9f", X"a3", X"94", X"84", X"78", X"6a", X"6e", X"5f", X"61", X"57", X"4d", X"51", X"53", X"46", X"50", X"44", X"4c", X"3d", X"29", X"1b", X"0d", X"06", X"04", X"12", X"06", X"09", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"12", X"06", X"09", X"16", X"0e", X"12", X"0f", X"17", X"16", X"32", X"58", X"82", X"b4", X"c9", X"94", X"83", X"7e", X"84", X"87", X"92", X"8d", X"8d", X"8b", X"91", X"8c", X"8b", X"89", X"99", X"a0", X"a3", X"ab", X"b3", X"bc", X"cc", X"c8", X"d0", X"d7", X"d5", X"d2", X"d5", X"dc", X"d6", X"da", X"d5", X"d6", X"d5", X"d9", X"e4", X"e1", X"e8", X"e7", X"e5", X"e7", X"ed", X"ed", X"ec", X"f5", X"f8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f8", X"ff", X"ff", X"ff", X"fe", X"f9", X"ff", X"f5", X"fa", X"f9", X"f7", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f7", X"ec", X"ea", X"e0", X"d9", X"d6", X"cf", X"bf", X"b7", X"b8", X"b5", X"ab", X"a9", X"a5", X"94", X"99", X"96", X"89", X"7c", X"72", X"6d", X"69", X"65", X"55", X"5c", X"53", X"55", X"4e", X"50", X"54", X"54", X"55", X"38", X"24", X"11", X"0e", X"0b", X"09", X"0b", X"0c", X"01", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"07", X"13", X"14", X"11", X"11", X"18", X"1c", X"2a", X"3e", X"6e", X"9d", X"c5", X"bd", X"9a", X"8c", X"89", X"93", X"95", X"95", X"99", X"97", X"97", X"94", X"91", X"95", X"99", X"9e", X"9f", X"aa", X"b2", X"b4", X"b8", X"c0", X"c3", X"ca", X"d3", X"d1", X"d6", X"d3", X"cb", X"d7", X"d2", X"ce", X"d5", X"de", X"db", X"e0", X"e2", X"e7", X"eb", X"ec", X"e2", X"f1", X"e7", X"f4", X"f6", X"fd", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f9", X"fc", X"f4", X"f7", X"ff", X"fd", X"f5", X"f5", X"ef", X"ee", X"f0", X"f4", X"f5", X"f4", X"f4", X"ff", X"ff", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"ff", X"fe", X"fb", X"fb", X"e9", X"e4", X"dc", X"da", X"cb", X"ca", X"c2", X"b8", X"b7", X"b6", X"aa", X"a8", X"a4", X"98", X"9f", X"94", X"8e", X"7f", X"7a", X"74", X"62", X"61", X"59", X"5a", X"5e", X"59", X"56", X"5e", X"5b", X"66", X"62", X"49", X"3a", X"24", X"10", X"0e", X"06", X"07", X"10", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"0e", X"12", X"1b", X"15", X"14", X"1b", X"20", X"37", X"4d", X"84", X"b2", X"c7", X"a5", X"a2", X"9e", X"91", X"95", X"9b", X"9b", X"9d", X"9a", X"a5", X"a4", X"9e", X"a5", X"a3", X"a5", X"a6", X"ab", X"ae", X"b7", X"bf", X"c5", X"c5", X"c6", X"d1", X"cf", X"d5", X"d0", X"c9", X"c8", X"cb", X"d3", X"d6", X"d7", X"e0", X"dd", X"e8", X"e9", X"e2", X"e8", X"e7", X"e9", X"f3", X"f5", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"fe", X"f4", X"f4", X"fd", X"fe", X"f9", X"f0", X"f2", X"ec", X"eb", X"e7", X"e9", X"f2", X"fc", X"f4", X"fc", X"fd", X"fa", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"ff", X"fc", X"f9", X"f0", X"e7", X"df", X"dd", X"d9", X"d0", X"ca", X"c2", X"ba", X"bd", X"b6", X"ad", X"a5", X"9d", X"9c", X"94", X"92", X"8d", X"81", X"7a", X"6f", X"5e", X"6f", X"64", X"67", X"5e", X"5d", X"59", X"69", X"6f", X"7c", X"73", X"65", X"43", X"25", X"1c", X"18", X"0d", X"15", X"12", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"0a", X"0a", X"06", X"11", X"14", X"1c", X"17", X"19", X"22", X"29", X"3e", X"68", X"a0", X"c0", X"be", X"ab", X"a8", X"a3", X"a0", X"a6", X"ae", X"a7", X"b0", X"af", X"ae", X"aa", X"b2", X"aa", X"af", X"b8", X"b5", X"b3", X"ba", X"c0", X"bd", X"c7", X"ce", X"c7", X"d1", X"d7", X"d3", X"d6", X"c9", X"cc", X"d2", X"cf", X"d2", X"dd", X"e1", X"e2", X"e0", X"e9", X"e3", X"e7", X"e6", X"f2", X"f5", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fe", X"ff", X"f5", X"f7", X"fe", X"f8", X"f0", X"ed", X"ec", X"ec", X"ed", X"e9", X"e9", X"fa", X"f4", X"f5", X"f8", X"fb", X"ff", X"ff", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"f5", X"ef", X"f0", X"ef", X"e6", X"e0", X"d8", X"d2", X"c7", X"ca", X"c0", X"bd", X"b5", X"ab", X"a8", X"9b", X"9f", X"94", X"91", X"92", X"8a", X"7d", X"7e", X"6e", X"70", X"61", X"6c", X"70", X"67", X"63", X"70", X"79", X"80", X"82", X"6e", X"5e", X"4b", X"2f", X"1a", X"10", X"0a", X"16", X"0e", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"08", X"17", X"18", X"0e", X"14", X"21", X"2f", X"48", X"70", X"94", X"ac", X"b0", X"ba", X"b0", X"b2", X"ad", X"aa", X"ad", X"b0", X"af", X"b6", X"ad", X"b3", X"b3", X"b9", X"b3", X"bc", X"b3", X"bd", X"bf", X"c0", X"be", X"cb", X"cb", X"ce", X"d3", X"d4", X"d7", X"cd", X"d8", X"cb", X"d7", X"d2", X"d2", X"da", X"e1", X"e1", X"e8", X"ec", X"e6", X"f1", X"ed", X"f0", X"f3", X"fd", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"ff", X"fc", X"f2", X"f3", X"f6", X"f7", X"f1", X"eb", X"e3", X"e4", X"e6", X"e3", X"eb", X"e8", X"f1", X"f5", X"f6", X"f9", X"f8", X"f9", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"f0", X"f2", X"e5", X"e6", X"e0", X"e3", X"d7", X"d6", X"cd", X"cf", X"c4", X"be", X"b7", X"af", X"ad", X"a5", X"9b", X"95", X"90", X"8f", X"8d", X"7a", X"7e", X"6f", X"70", X"68", X"70", X"75", X"7f", X"75", X"82", X"80", X"84", X"88", X"8a", X"73", X"5c", X"3c", X"25", X"1f", X"22", X"12", X"07", X"0c", X"05", X"05", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0d", X"09", X"18", X"1a", X"16", X"1e", X"1e", X"40", X"57", X"74", X"84", X"96", X"a5", X"b3", X"c5", X"b8", X"b7", X"b2", X"b8", X"b1", X"b8", X"b9", X"b8", X"ba", X"c0", X"c2", X"bf", X"be", X"c2", X"c8", X"c1", X"c4", X"c3", X"c7", X"c8", X"d1", X"d4", X"cb", X"d0", X"ca", X"c3", X"cd", X"c9", X"d0", X"d5", X"dd", X"e4", X"e9", X"e9", X"ec", X"e7", X"ef", X"ea", X"f5", X"f9", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"f3", X"fb", X"f5", X"f0", X"f5", X"fc", X"f4", X"e4", X"e2", X"de", X"e1", X"e9", X"e2", X"ea", X"e5", X"eb", X"ec", X"f2", X"f0", X"f0", X"fd", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"f1", X"e8", X"e6", X"e4", X"df", X"de", X"d9", X"d6", X"ca", X"c7", X"c7", X"bd", X"af", X"af", X"9b", X"9c", X"99", X"96", X"93", X"86", X"83", X"75", X"6d", X"68", X"77", X"80", X"81", X"90", X"8c", X"90", X"8b", X"89", X"86", X"87", X"81", X"68", X"49", X"2b", X"1d", X"1a", X"15", X"0d", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"09", X"0a", X"06", X"05", X"0a", X"0e", X"06", X"0e", X"20", X"25", X"27", X"35", X"4a", X"67", X"7e", X"84", X"8d", X"98", X"a7", X"bd", X"c5", X"ce", X"ca", X"c8", X"c3", X"c0", X"b8", X"c1", X"c1", X"bc", X"c9", X"cc", X"c7", X"c8", X"c8", X"c3", X"c7", X"cd", X"cd", X"cd", X"cc", X"d0", X"ca", X"cc", X"ce", X"d1", X"c9", X"d4", X"d1", X"d4", X"dc", X"e1", X"e9", X"eb", X"ed", X"ed", X"ec", X"f2", X"f5", X"fc", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"f5", X"fb", X"f8", X"eb", X"f8", X"fb", X"fc", X"ea", X"e5", X"dc", X"df", X"e1", X"e0", X"e7", X"f0", X"e7", X"e5", X"f0", X"ed", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"ff", X"ff", X"fd", X"eb", X"d8", X"dc", X"d9", X"e0", X"cf", X"c9", X"c7", X"c3", X"b6", X"b1", X"ad", X"a5", X"9e", X"98", X"8b", X"87", X"82", X"80", X"80", X"7c", X"8b", X"9b", X"9e", X"9b", X"95", X"99", X"97", X"88", X"7f", X"83", X"99", X"77", X"5a", X"37", X"1b", X"0d", X"11", X"03", X"06", X"05", X"03", X"03", X"06", X"09", X"03", X"00", X"06", X"05", X"07", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"08", X"0a", X"05", X"03", X"03", X"0a", X"11", X"1b", X"2b", X"34", X"44", X"58", X"70", X"73", X"84", X"7a", X"8d", X"a7", X"ba", X"c5", X"d8", X"cc", X"bb", X"cc", X"bd", X"c4", X"d5", X"cc", X"d0", X"cd", X"c6", X"d1", X"cc", X"ca", X"c3", X"cb", X"ce", X"ce", X"d0", X"d1", X"d0", X"cd", X"d0", X"d2", X"d1", X"d1", X"d6", X"d7", X"d4", X"e7", X"ef", X"e3", X"ee", X"ef", X"ef", X"f6", X"f5", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"f8", X"f9", X"f6", X"ed", X"f3", X"f8", X"f8", X"ed", X"e6", X"dc", X"e1", X"e0", X"e5", X"e5", X"e2", X"ea", X"ec", X"ea", X"f3", X"f7", X"fb", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ef", X"e3", X"ea", X"e2", X"e1", X"df", X"d5", X"c5", X"c0", X"bd", X"b0", X"a1", X"9a", X"90", X"89", X"92", X"84", X"89", X"96", X"a4", X"a9", X"a6", X"a9", X"a5", X"ae", X"99", X"87", X"86", X"8d", X"a2", X"8f", X"61", X"3e", X"2b", X"1d", X"14", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"02", X"09", X"05", X"03", X"0a", X"0d", X"20", X"23", X"34", X"3e", X"4b", X"64", X"70", X"71", X"7d", X"8a", X"90", X"95", X"9f", X"c1", X"cb", X"d0", X"ca", X"c3", X"d0", X"d1", X"ce", X"d5", X"dc", X"d6", X"d2", X"cf", X"d9", X"cf", X"d2", X"d2", X"c7", X"ce", X"d0", X"d2", X"ce", X"d4", X"ce", X"d7", X"d4", X"ce", X"d7", X"e2", X"df", X"de", X"ef", X"f3", X"e9", X"f6", X"f6", X"f7", X"fc", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f5", X"f2", X"f3", X"f2", X"eb", X"f4", X"ed", X"ed", X"df", X"e7", X"e0", X"e2", X"db", X"e2", X"e3", X"e0", X"e4", X"ec", X"ef", X"f0", X"f7", X"fa", X"fe", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"e4", X"e4", X"e1", X"e1", X"e1", X"dc", X"d7", X"c7", X"bd", X"b2", X"a7", X"93", X"8a", X"91", X"99", X"a8", X"b5", X"b3", X"b7", X"b4", X"ac", X"b5", X"b6", X"96", X"8f", X"89", X"8e", X"99", X"99", X"63", X"41", X"28", X"16", X"15", X"0b", X"06", X"05", X"0a", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"05", X"06", X"0a", X"14", X"10", X"15", X"1d", X"36", X"44", X"55", X"54", X"6b", X"75", X"86", X"7b", X"8d", X"8e", X"9a", X"a2", X"bd", X"cc", X"d4", X"d5", X"d7", X"d2", X"d6", X"e3", X"db", X"de", X"df", X"d3", X"dc", X"e0", X"da", X"cf", X"cf", X"d9", X"d5", X"da", X"e3", X"d3", X"d9", X"d5", X"dd", X"df", X"df", X"d9", X"e0", X"e5", X"ed", X"e8", X"f1", X"f5", X"f8", X"fb", X"f9", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"fb", X"fc", X"f3", X"f3", X"f8", X"ef", X"f5", X"ee", X"f4", X"ed", X"e4", X"d8", X"dd", X"de", X"db", X"e1", X"de", X"e5", X"e8", X"e7", X"e8", X"e8", X"f1", X"f0", X"f5", X"f9", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"e0", X"df", X"e1", X"de", X"d9", X"d7", X"cc", X"c1", X"b4", X"af", X"a1", X"9a", X"97", X"a6", X"b8", X"ce", X"c4", X"c8", X"bd", X"c6", X"b4", X"af", X"a0", X"96", X"92", X"95", X"aa", X"a5", X"72", X"49", X"20", X"1b", X"16", X"0d", X"06", X"05", X"03", X"06", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"02", X"06", X"09", X"0f", X"10", X"1f", X"26", X"3d", X"55", X"65", X"6e", X"72", X"85", X"82", X"88", X"86", X"97", X"9d", X"a6", X"b3", X"d1", X"dc", X"cf", X"d3", X"d7", X"d9", X"e5", X"e3", X"de", X"e6", X"e6", X"e4", X"e4", X"de", X"db", X"df", X"dd", X"df", X"d8", X"e1", X"e0", X"de", X"e3", X"e0", X"ec", X"db", X"e5", X"ef", X"f0", X"f7", X"f5", X"fc", X"ff", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"ff", X"fc", X"fd", X"f9", X"f4", X"f2", X"f2", X"eb", X"e7", X"ed", X"e5", X"d5", X"da", X"d4", X"de", X"df", X"e0", X"e1", X"e7", X"e7", X"ef", X"e8", X"ee", X"f6", X"f2", X"f8", X"fb", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f4", X"e7", X"e1", X"d6", X"d5", X"cf", X"cd", X"c4", X"bf", X"b2", X"ae", X"ab", X"a2", X"ad", X"c2", X"d9", X"d5", X"d0", X"c6", X"c8", X"c1", X"c0", X"ac", X"a9", X"95", X"a0", X"9c", X"b1", X"a4", X"6f", X"43", X"25", X"13", X"13", X"08", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"07", X"06", X"05", X"03", X"13", X"1c", X"33", X"4a", X"5b", X"75", X"76", X"80", X"82", X"89", X"86", X"94", X"a1", X"a1", X"a5", X"b1", X"d0", X"e9", X"d2", X"d0", X"cd", X"d5", X"e4", X"df", X"e6", X"e8", X"e8", X"ea", X"ea", X"e3", X"e2", X"eb", X"e0", X"e9", X"e3", X"e5", X"e8", X"eb", X"e0", X"ea", X"ec", X"f2", X"eb", X"f4", X"f8", X"f3", X"f7", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"f6", X"fa", X"fa", X"f3", X"f0", X"ed", X"eb", X"e1", X"db", X"dd", X"dd", X"e4", X"db", X"de", X"e1", X"e6", X"e6", X"ea", X"e1", X"e3", X"e1", X"ef", X"f5", X"fd", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"f4", X"ec", X"e8", X"de", X"e4", X"d3", X"d1", X"ca", X"c0", X"bd", X"b6", X"af", X"b4", X"b2", X"bf", X"d7", X"e6", X"db", X"dc", X"ce", X"c4", X"c1", X"b8", X"b6", X"b1", X"b4", X"a9", X"9e", X"b0", X"a2", X"64", X"31", X"1e", X"13", X"07", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"06", X"0a", X"12", X"0d", X"0f", X"14", X"2a", X"3b", X"4d", X"66", X"80", X"75", X"7e", X"8f", X"89", X"93", X"98", X"9c", X"a1", X"ae", X"b4", X"cc", X"f0", X"df", X"d7", X"d0", X"d1", X"e2", X"e4", X"e2", X"f1", X"e6", X"ed", X"ef", X"ea", X"eb", X"e5", X"eb", X"ed", X"f0", X"ed", X"f7", X"f0", X"f0", X"f0", X"f0", X"f6", X"f7", X"fa", X"f8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"f8", X"ec", X"e4", X"e9", X"e2", X"dd", X"d8", X"de", X"da", X"dd", X"dd", X"e7", X"e3", X"dc", X"ee", X"e9", X"e2", X"f1", X"f1", X"f6", X"ee", X"fd", X"ff", X"ff", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ee", X"ed", X"e1", X"dd", X"d7", X"d7", X"ce", X"d0", X"c0", X"b3", X"b3", X"ae", X"af", X"cb", X"d6", X"e9", X"e6", X"e6", X"e0", X"d1", X"c8", X"c4", X"b6", X"bb", X"bb", X"b6", X"a9", X"aa", X"aa", X"9e", X"5f", X"32", X"18", X"10", X"0f", X"02", X"09", X"06", X"03", X"01", X"06", X"05", X"03", X"00", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"10", X"14", X"0d", X"17", X"1f", X"31", X"3e", X"54", X"78", X"89", X"83", X"84", X"91", X"95", X"9d", X"a0", X"ab", X"a6", X"b0", X"ae", X"c2", X"ea", X"e4", X"d7", X"d7", X"d3", X"db", X"e2", X"ea", X"ec", X"ee", X"f0", X"ec", X"ea", X"f0", X"f2", X"f4", X"fa", X"f5", X"f3", X"f0", X"eb", X"f7", X"f9", X"f5", X"ff", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"f3", X"f6", X"e3", X"dc", X"db", X"db", X"e2", X"e5", X"e3", X"df", X"df", X"e3", X"e8", X"e3", X"ea", X"e6", X"eb", X"ef", X"fa", X"ee", X"f4", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"e9", X"e6", X"e1", X"d6", X"d1", X"d1", X"c9", X"bc", X"bf", X"b0", X"b8", X"c9", X"db", X"e5", X"f6", X"ed", X"e5", X"de", X"d3", X"c7", X"c1", X"af", X"be", X"b3", X"ae", X"a7", X"a2", X"ad", X"7f", X"4b", X"29", X"15", X"14", X"0e", X"0a", X"09", X"05", X"0a", X"01", X"06", X"05", X"03", X"00", X"0a", X"05", X"03", X"00", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"16", X"15", X"13", X"22", X"32", X"44", X"67", X"87", X"9d", X"8e", X"89", X"96", X"9b", X"99", X"9e", X"a0", X"ae", X"ae", X"b3", X"c0", X"e4", X"e3", X"d5", X"d4", X"d3", X"d8", X"d9", X"e7", X"e5", X"e6", X"f3", X"f1", X"f0", X"f4", X"ef", X"f3", X"f8", X"f9", X"f3", X"f7", X"f5", X"f9", X"f5", X"f7", X"f7", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"fb", X"fd", X"ff", X"ff", X"ff", X"ff", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"e8", X"e3", X"e5", X"e0", X"e4", X"e0", X"e3", X"e4", X"e0", X"eb", X"e5", X"e1", X"e4", X"e9", X"e6", X"e5", X"ed", X"ec", X"f2", X"f7", X"f6", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"f6", X"f9", X"f2", X"eb", X"e5", X"dd", X"d9", X"ca", X"bf", X"c5", X"b9", X"b8", X"ae", X"c1", X"e6", X"f4", X"ef", X"f0", X"f6", X"e4", X"d0", X"cb", X"bd", X"bb", X"b9", X"ae", X"aa", X"a5", X"a1", X"99", X"9c", X"68", X"37", X"22", X"18", X"0d", X"0b", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"09", X"0d", X"17", X"12", X"12", X"22", X"30", X"43", X"75", X"90", X"a9", X"aa", X"97", X"95", X"9f", X"a3", X"a3", X"af", X"bb", X"c0", X"d2", X"e2", X"ec", X"eb", X"cf", X"d1", X"cf", X"d4", X"d9", X"dc", X"e5", X"e9", X"ec", X"e9", X"ee", X"f3", X"f4", X"ee", X"fa", X"f6", X"f4", X"fa", X"fa", X"f5", X"fc", X"fc", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"fe", X"f9", X"f1", X"f6", X"f7", X"f7", X"f8", X"fb", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f0", X"e6", X"e1", X"d9", X"da", X"de", X"df", X"e1", X"de", X"e1", X"e6", X"ec", X"e9", X"e6", X"e7", X"ef", X"f3", X"ef", X"ed", X"f8", X"e7", X"f4", X"f6", X"fa", X"f9", X"f9", X"f1", X"f4", X"f3", X"f3", X"ec", X"ea", X"e3", X"d5", X"d6", X"cb", X"bd", X"bd", X"bd", X"b5", X"b3", X"c3", X"de", X"f5", X"fb", X"f9", X"e8", X"d8", X"d5", X"c6", X"c4", X"b7", X"b9", X"b0", X"a3", X"a2", X"97", X"91", X"81", X"4d", X"24", X"1e", X"0d", X"16", X"15", X"0e", X"06", X"07", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"02", X"06", X"0a", X"0e", X"11", X"17", X"0d", X"1b", X"1e", X"25", X"4c", X"78", X"91", X"a5", X"b4", X"aa", X"a7", X"9c", X"b0", X"a8", X"b0", X"c3", X"c9", X"db", X"ee", X"f7", X"f5", X"da", X"d4", X"c1", X"db", X"e1", X"de", X"e7", X"ea", X"e1", X"e9", X"f4", X"f0", X"f2", X"f1", X"f7", X"ea", X"f3", X"ff", X"fc", X"fb", X"ff", X"f8", X"fd", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"f7", X"f4", X"f4", X"ec", X"f3", X"e5", X"eb", X"f3", X"ec", X"f0", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"fa", X"f1", X"e3", X"e5", X"e2", X"e3", X"e2", X"e5", X"df", X"df", X"e4", X"ed", X"ed", X"ea", X"eb", X"f1", X"ec", X"e9", X"ee", X"f3", X"f2", X"f4", X"f4", X"f1", X"f0", X"f1", X"ed", X"f1", X"ee", X"ed", X"e8", X"db", X"d9", X"d6", X"c9", X"c2", X"c0", X"bd", X"b4", X"c0", X"c5", X"de", X"f8", X"ff", X"f9", X"eb", X"db", X"d2", X"c6", X"b8", X"b5", X"b0", X"a5", X"a1", X"97", X"84", X"7c", X"5a", X"36", X"1e", X"1a", X"14", X"16", X"11", X"0b", X"06", X"05", X"06", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"04", X"0e", X"0e", X"13", X"1a", X"23", X"2d", X"4b", X"7c", X"90", X"a0", X"b5", X"bf", X"bc", X"b0", X"a9", X"b5", X"b6", X"c2", X"d3", X"d2", X"e0", X"e7", X"ef", X"d4", X"cf", X"c6", X"cb", X"cb", X"d8", X"e0", X"db", X"e7", X"e7", X"e9", X"ed", X"ee", X"f0", X"ef", X"f1", X"f8", X"f0", X"f3", X"f9", X"fa", X"fd", X"fb", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"f0", X"f2", X"ed", X"ec", X"e5", X"e8", X"ec", X"ee", X"ea", X"ec", X"e9", X"e4", X"e2", X"e9", X"e5", X"f5", X"f5", X"f6", X"f5", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ed", X"ea", X"e0", X"df", X"df", X"e4", X"df", X"e2", X"e8", X"ed", X"e9", X"ed", X"e8", X"fa", X"f0", X"ed", X"f0", X"eb", X"f0", X"f6", X"ef", X"f3", X"ed", X"f0", X"ed", X"e7", X"ea", X"f2", X"e7", X"e0", X"d8", X"d4", X"d1", X"c7", X"c1", X"bf", X"c4", X"c8", X"d5", X"f6", X"ff", X"f8", X"e6", X"de", X"d4", X"c6", X"bc", X"b7", X"ac", X"ae", X"a2", X"a0", X"90", X"7d", X"5e", X"36", X"1e", X"1b", X"19", X"11", X"10", X"10", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0d", X"07", X"11", X"12", X"27", X"35", X"4f", X"78", X"8e", X"a7", X"b1", X"c2", X"d8", X"c1", X"ba", X"be", X"c2", X"ca", X"ca", X"cf", X"d3", X"e5", X"e5", X"d5", X"cb", X"c4", X"d0", X"d0", X"d6", X"df", X"dd", X"e4", X"e0", X"ed", X"e7", X"e8", X"f1", X"f2", X"ec", X"eb", X"fe", X"f3", X"f5", X"f8", X"ef", X"f4", X"fb", X"ff", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"ff", X"fa", X"f5", X"f9", X"ff", X"fc", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fa", X"ec", X"e3", X"e3", X"da", X"d4", X"da", X"d3", X"db", X"db", X"d7", X"d2", X"e0", X"dc", X"dc", X"dc", X"de", X"df", X"ed", X"ed", X"ef", X"f5", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f0", X"ea", X"ed", X"e3", X"df", X"da", X"dc", X"de", X"db", X"e2", X"ef", X"ef", X"f7", X"fa", X"f2", X"f1", X"f0", X"ee", X"f7", X"f8", X"f1", X"ef", X"f0", X"ea", X"f3", X"e2", X"e2", X"ea", X"e6", X"e3", X"d7", X"e2", X"e1", X"c9", X"cb", X"c3", X"d5", X"dd", X"dc", X"e8", X"f3", X"e4", X"d6", X"d1", X"c4", X"c3", X"bd", X"b4", X"af", X"a8", X"a0", X"8c", X"84", X"64", X"45", X"31", X"21", X"16", X"16", X"13", X"0c", X"17", X"05", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"06", X"04", X"07", X"05", X"06", X"0d", X"11", X"0f", X"16", X"23", X"31", X"56", X"7a", X"8f", X"a0", X"b1", X"b7", X"dd", X"db", X"d0", X"c5", X"cf", X"d2", X"d0", X"d1", X"d0", X"d8", X"d3", X"c9", X"ce", X"cf", X"cc", X"cf", X"d2", X"d0", X"d6", X"e5", X"df", X"e5", X"ec", X"e7", X"ec", X"ec", X"e8", X"f3", X"ee", X"f3", X"f3", X"f1", X"fc", X"fb", X"f9", X"ff", X"f9", X"f7", X"ff", X"fe", X"fe", X"ff", X"ff", X"f7", X"fb", X"fa", X"ff", X"ff", X"fe", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f2", X"f1", X"dc", X"db", X"cd", X"d0", X"cb", X"cd", X"d1", X"d2", X"d5", X"d3", X"d3", X"d7", X"d7", X"d2", X"d2", X"d4", X"dc", X"d5", X"db", X"e1", X"f5", X"f8", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f9", X"ec", X"e2", X"e4", X"de", X"e2", X"de", X"e0", X"e1", X"e6", X"f1", X"ea", X"f2", X"f6", X"f0", X"f2", X"f7", X"f2", X"f4", X"f5", X"fa", X"f4", X"ea", X"f0", X"e8", X"ed", X"f0", X"f4", X"ea", X"e7", X"f1", X"ea", X"d9", X"da", X"dc", X"d6", X"d9", X"d2", X"df", X"df", X"db", X"dd", X"c4", X"c5", X"c0", X"c0", X"b5", X"b5", X"a9", X"99", X"8f", X"77", X"56", X"34", X"2b", X"19", X"1d", X"1f", X"0e", X"13", X"11", X"10", X"07", X"07", X"08", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"08", X"07", X"12", X"14", X"0c", X"16", X"1b", X"2a", X"35", X"57", X"7b", X"86", X"96", X"a5", X"bb", X"d6", X"e0", X"d4", X"cc", X"c4", X"c8", X"c6", X"c9", X"c8", X"c3", X"c9", X"c9", X"c6", X"c6", X"cd", X"d3", X"d6", X"d6", X"dd", X"e1", X"e1", X"e0", X"e4", X"ed", X"e4", X"e8", X"ef", X"f5", X"f7", X"f1", X"f2", X"f2", X"f3", X"f3", X"f9", X"fd", X"fa", X"f9", X"ff", X"fb", X"ff", X"f7", X"f5", X"f6", X"f6", X"fe", X"f9", X"f7", X"ff", X"fd", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e8", X"e0", X"d1", X"d0", X"d5", X"ce", X"c2", X"ce", X"c7", X"ca", X"d1", X"d3", X"d2", X"db", X"cf", X"d6", X"cc", X"cf", X"d8", X"cd", X"e2", X"d5", X"e3", X"e8", X"ed", X"f4", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"f5", X"eb", X"e8", X"e8", X"e4", X"e1", X"e4", X"e6", X"e0", X"e9", X"ec", X"e8", X"f2", X"ef", X"f4", X"f5", X"f7", X"ee", X"f3", X"f1", X"f0", X"f0", X"f0", X"e3", X"eb", X"ec", X"e9", X"e9", X"e1", X"e6", X"f0", X"e3", X"d8", X"d5", X"d3", X"d2", X"d2", X"d0", X"d1", X"d1", X"ca", X"cd", X"bd", X"c9", X"bb", X"bd", X"b5", X"b6", X"a7", X"94", X"7b", X"5e", X"35", X"25", X"24", X"1b", X"1a", X"12", X"14", X"14", X"0f", X"12", X"07", X"0d", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"03", X"09", X"06", X"08", X"05", X"0c", X"10", X"10", X"1e", X"2d", X"3b", X"52", X"6d", X"80", X"8e", X"99", X"aa", X"c6", X"d0", X"cf", X"c6", X"ba", X"c1", X"c4", X"c3", X"bd", X"c0", X"c0", X"c5", X"c6", X"c6", X"c7", X"c8", X"d3", X"d6", X"d6", X"df", X"d9", X"d9", X"df", X"e1", X"e1", X"e7", X"eb", X"eb", X"ec", X"e7", X"f1", X"f0", X"f4", X"f5", X"f8", X"f9", X"fb", X"fb", X"f7", X"f7", X"fc", X"fa", X"f7", X"fb", X"fa", X"fb", X"f1", X"f7", X"f9", X"fe", X"f9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e0", X"dd", X"ce", X"cd", X"cf", X"cf", X"cf", X"cd", X"d0", X"d2", X"c9", X"d3", X"ca", X"d4", X"d4", X"d4", X"d1", X"d2", X"cb", X"cb", X"d2", X"ce", X"d6", X"dc", X"e2", X"ed", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fb", X"ee", X"e7", X"e0", X"e3", X"dd", X"e2", X"ee", X"e2", X"eb", X"e9", X"e8", X"ea", X"f5", X"f7", X"f7", X"f2", X"f2", X"ef", X"e2", X"e6", X"e9", X"e2", X"e2", X"e6", X"e4", X"e6", X"e3", X"db", X"dd", X"d8", X"d9", X"d2", X"d3", X"d2", X"ca", X"d4", X"d0", X"c8", X"c7", X"c5", X"c7", X"c8", X"bf", X"c0", X"b2", X"a5", X"a5", X"86", X"6d", X"42", X"34", X"20", X"1a", X"15", X"15", X"17", X"18", X"0f", X"0d", X"06", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"01", X"06", X"0c", X"0e", X"16", X"19", X"1a", X"29", X"25", X"39", X"52", X"79", X"83", X"89", X"8f", X"a7", X"b0", X"c2", X"bf", X"bc", X"b8", X"bc", X"bf", X"c0", X"b8", X"bd", X"bd", X"ba", X"c4", X"c8", X"c4", X"cd", X"d0", X"da", X"d0", X"d5", X"db", X"dc", X"df", X"e5", X"e8", X"e5", X"e8", X"eb", X"ef", X"ec", X"f0", X"f5", X"f9", X"f6", X"f2", X"f5", X"ef", X"f5", X"f9", X"f1", X"f3", X"f0", X"f3", X"f5", X"f4", X"f6", X"f9", X"f7", X"f8", X"fb", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"fd", X"f5", X"ef", X"f4", X"fb", X"f5", X"f5", X"fb", X"f6", X"fb", X"fb", X"f3", X"f7", X"f1", X"f8", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e1", X"d9", X"cf", X"ce", X"d0", X"d0", X"c6", X"cf", X"cd", X"d0", X"d1", X"cd", X"d5", X"d6", X"d2", X"d4", X"d0", X"d1", X"ca", X"c5", X"cb", X"cd", X"cf", X"da", X"df", X"eb", X"f2", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f8", X"f3", X"e6", X"e7", X"ea", X"e2", X"db", X"eb", X"ee", X"ee", X"e9", X"ed", X"eb", X"f2", X"f5", X"f6", X"f1", X"ed", X"eb", X"ec", X"e6", X"e7", X"e3", X"de", X"e0", X"e0", X"de", X"de", X"d6", X"d8", X"dc", X"d0", X"d5", X"cf", X"d4", X"c9", X"d1", X"d3", X"c7", X"c9", X"c7", X"ca", X"c2", X"b9", X"ba", X"a5", X"a4", X"94", X"78", X"4c", X"39", X"28", X"1a", X"23", X"16", X"1a", X"15", X"14", X"0d", X"12", X"0e", X"13", X"0e", X"0d", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"05", X"03", X"06", X"05", X"03", X"00", X"06", X"06", X"0a", X"0d", X"21", X"1e", X"2a", X"2f", X"33", X"4f", X"74", X"84", X"87", X"8b", X"96", X"a1", X"aa", X"b0", X"a6", X"ac", X"b8", X"c7", X"b6", X"b8", X"b8", X"c0", X"c4", X"c3", X"c6", X"c9", X"d0", X"d0", X"d6", X"d5", X"d6", X"df", X"db", X"e2", X"e3", X"e3", X"e5", X"e4", X"e6", X"ec", X"e7", X"e3", X"ef", X"f1", X"f2", X"ee", X"e9", X"f0", X"f5", X"f5", X"f7", X"f3", X"f4", X"f5", X"fd", X"f5", X"f8", X"f9", X"f4", X"f6", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fd", X"fd", X"ff", X"ff", X"ff", X"f7", X"fb", X"f3", X"f0", X"eb", X"e8", X"ef", X"e6", X"f2", X"f1", X"ef", X"ef", X"f5", X"f0", X"ef", X"f0", X"f1", X"f8", X"f5", X"f2", X"fd", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ec", X"dc", X"cf", X"cd", X"d2", X"d0", X"c2", X"d2", X"d0", X"cd", X"d6", X"ca", X"d5", X"d7", X"d2", X"ce", X"cd", X"ca", X"ca", X"cc", X"c9", X"c5", X"c7", X"cd", X"cb", X"d6", X"eb", X"e9", X"ff", X"ff", X"ff", X"ff", X"ff", X"ef", X"ea", X"e7", X"e9", X"e4", X"ee", X"e5", X"e4", X"e1", X"e9", X"ee", X"ec", X"eb", X"e6", X"f1", X"f5", X"ed", X"f0", X"e8", X"ee", X"f0", X"e8", X"ea", X"e5", X"e0", X"e3", X"e2", X"e0", X"de", X"dd", X"d4", X"cf", X"d6", X"ce", X"d1", X"d4", X"ce", X"cf", X"c4", X"c5", X"c9", X"ce", X"c6", X"bd", X"b3", X"a6", X"a4", X"85", X"60", X"41", X"2e", X"29", X"23", X"24", X"17", X"1b", X"16", X"15", X"11", X"13", X"11", X"0a", X"07", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"0a", X"05", X"03", X"02", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"03", X"06", X"10", X"0e", X"15", X"11", X"18", X"26", X"24", X"30", X"46", X"73", X"80", X"8b", X"90", X"89", X"93", X"9b", X"9c", X"a1", X"b0", X"b5", X"b0", X"b8", X"b3", X"b5", X"bb", X"bb", X"c9", X"c6", X"cd", X"d0", X"c7", X"d3", X"d1", X"dc", X"d3", X"e3", X"e2", X"e6", X"e0", X"e0", X"dc", X"e7", X"e7", X"e5", X"eb", X"e9", X"ed", X"ef", X"ef", X"ee", X"ee", X"f6", X"ee", X"f2", X"f4", X"f2", X"ee", X"ee", X"ef", X"f6", X"f6", X"f3", X"f9", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fc", X"f9", X"f3", X"fe", X"fc", X"fd", X"f6", X"fc", X"f1", X"ec", X"e2", X"e7", X"da", X"e7", X"e5", X"e6", X"f3", X"f4", X"f1", X"ec", X"e9", X"e7", X"e9", X"f3", X"ea", X"f0", X"f6", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ee", X"de", X"d7", X"cf", X"d3", X"cf", X"ca", X"cb", X"cc", X"d3", X"d4", X"ce", X"ce", X"ce", X"cd", X"d3", X"cc", X"cb", X"c7", X"c8", X"c9", X"c5", X"c1", X"c7", X"ca", X"cf", X"d1", X"df", X"f3", X"ff", X"ff", X"ff", X"fc", X"f7", X"ed", X"ef", X"ed", X"f0", X"f1", X"f0", X"eb", X"ec", X"eb", X"ec", X"ec", X"e8", X"e8", X"e9", X"e4", X"f0", X"eb", X"eb", X"e9", X"e5", X"e8", X"e4", X"e0", X"e3", X"dd", X"e3", X"de", X"db", X"db", X"db", X"d7", X"d0", X"d6", X"d8", X"cd", X"d2", X"d0", X"c6", X"c0", X"c0", X"c7", X"b9", X"ad", X"ae", X"9f", X"89", X"6d", X"4e", X"2f", X"28", X"27", X"27", X"1e", X"1b", X"11", X"12", X"16", X"12", X"11", X"0e", X"06", X"08", X"03", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"0a", X"06", X"0c", X"10", X"15", X"1b", X"2a", X"24", X"25", X"48", X"71", X"8c", X"92", X"8d", X"93", X"8f", X"95", X"97", X"9b", X"9c", X"ae", X"a5", X"a4", X"ad", X"b6", X"bf", X"c0", X"c5", X"c4", X"c9", X"c6", X"cd", X"cf", X"d1", X"da", X"df", X"d7", X"de", X"e4", X"e2", X"de", X"e1", X"e5", X"e9", X"e8", X"e8", X"ee", X"e8", X"f1", X"e7", X"ed", X"e5", X"f0", X"f5", X"f3", X"ee", X"f4", X"f2", X"ea", X"ec", X"f1", X"f6", X"e9", X"ef", X"f4", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"f5", X"f3", X"ed", X"ef", X"ee", X"e7", X"f5", X"f5", X"f0", X"f2", X"e9", X"ec", X"e7", X"ea", X"de", X"d8", X"e0", X"e9", X"ed", X"ea", X"ee", X"ea", X"e5", X"eb", X"e7", X"f1", X"e9", X"f5", X"f8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e5", X"d7", X"db", X"c7", X"d0", X"bd", X"ca", X"c8", X"cc", X"d5", X"d3", X"d4", X"d5", X"d1", X"cd", X"c8", X"cd", X"cd", X"cb", X"c6", X"be", X"b9", X"c4", X"c2", X"c6", X"c7", X"d8", X"e7", X"f0", X"fd", X"f8", X"f9", X"f3", X"e9", X"eb", X"ea", X"f4", X"f7", X"fc", X"f7", X"ef", X"f1", X"f6", X"fb", X"ee", X"f1", X"ee", X"e9", X"f0", X"f4", X"ed", X"ed", X"e0", X"e5", X"e1", X"e2", X"e1", X"e4", X"e8", X"e7", X"e0", X"db", X"de", X"cf", X"cd", X"d4", X"d4", X"d8", X"d5", X"cf", X"c5", X"bc", X"c6", X"be", X"b4", X"b5", X"a4", X"92", X"84", X"65", X"46", X"2d", X"20", X"27", X"2b", X"19", X"18", X"1b", X"0e", X"10", X"14", X"11", X"0e", X"0d", X"07", X"0c", X"09", X"06", X"05", X"03", X"00", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"02", X"06", X"07", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"02", X"08", X"09", X"0d", X"0c", X"16", X"27", X"32", X"24", X"28", X"47", X"6b", X"86", X"8c", X"93", X"90", X"92", X"94", X"94", X"93", X"97", X"9a", X"a2", X"a2", X"a7", X"b5", X"b6", X"c0", X"c4", X"c7", X"c8", X"cd", X"d3", X"cf", X"d3", X"d3", X"dc", X"d3", X"d4", X"de", X"e1", X"e2", X"e2", X"e0", X"e4", X"eb", X"e6", X"e7", X"f0", X"e2", X"f1", X"ec", X"e5", X"ef", X"f2", X"ed", X"f0", X"ed", X"ee", X"e9", X"ea", X"f3", X"f2", X"f6", X"f2", X"fc", X"ff", X"fc", X"f8", X"f8", X"f5", X"f0", X"e9", X"ee", X"e7", X"eb", X"ea", X"f2", X"f7", X"f8", X"f2", X"ee", X"ec", X"ee", X"e5", X"e6", X"e0", X"e1", X"e1", X"e1", X"de", X"ea", X"e7", X"ee", X"f3", X"e9", X"e5", X"f0", X"e9", X"f1", X"f3", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ec", X"db", X"cd", X"d4", X"d7", X"cf", X"c9", X"d0", X"c8", X"d1", X"d8", X"d0", X"d4", X"d9", X"cb", X"d3", X"d0", X"c7", X"cb", X"c7", X"be", X"c2", X"c4", X"bf", X"ba", X"c4", X"c6", X"d8", X"de", X"ee", X"eb", X"f0", X"ef", X"ea", X"e8", X"ef", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"f8", X"fb", X"ea", X"ef", X"f1", X"f3", X"f0", X"ed", X"ed", X"eb", X"e7", X"e0", X"e6", X"eb", X"e5", X"ec", X"e9", X"e2", X"e1", X"d6", X"da", X"d2", X"da", X"d2", X"cf", X"d0", X"cf", X"d1", X"d1", X"c1", X"c3", X"c3", X"ac", X"a0", X"9b", X"84", X"7d", X"57", X"3d", X"36", X"27", X"28", X"1e", X"1e", X"22", X"15", X"19", X"14", X"12", X"11", X"0a", X"09", X"0f", X"0c", X"0d", X"06", X"05", X"04", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"06", X"0a", X"09", X"17", X"1e", X"29", X"2a", X"2a", X"44", X"5f", X"71", X"7f", X"89", X"8f", X"96", X"97", X"90", X"90", X"91", X"92", X"9f", X"a5", X"ab", X"aa", X"b1", X"ba", X"bd", X"c2", X"cc", X"d2", X"c9", X"c6", X"d2", X"d4", X"d4", X"d4", X"d3", X"d4", X"e0", X"d9", X"e3", X"e3", X"db", X"e3", X"df", X"de", X"e3", X"e1", X"e4", X"e8", X"e2", X"ec", X"e4", X"e7", X"e6", X"e7", X"e1", X"e6", X"f0", X"f2", X"f5", X"f3", X"f4", X"fd", X"f5", X"f5", X"f1", X"ed", X"e3", X"e1", X"ea", X"e5", X"ea", X"f3", X"ee", X"ef", X"f4", X"f5", X"f5", X"f2", X"f1", X"ea", X"e7", X"e7", X"e0", X"e1", X"e2", X"e1", X"df", X"e8", X"e0", X"e7", X"e7", X"e5", X"eb", X"ec", X"e6", X"f2", X"ef", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f7", X"d8", X"ca", X"cb", X"cd", X"cb", X"cf", X"c7", X"d0", X"cd", X"d5", X"d0", X"d4", X"cc", X"d7", X"cd", X"c7", X"c1", X"bb", X"c5", X"c1", X"ba", X"bc", X"b9", X"ba", X"bd", X"b8", X"c2", X"ca", X"d8", X"d8", X"e3", X"e5", X"e4", X"e1", X"e7", X"ea", X"f5", X"ff", X"ff", X"ff", X"ff", X"fa", X"fc", X"ed", X"f2", X"ee", X"f3", X"f2", X"ef", X"f2", X"e9", X"ed", X"e9", X"eb", X"eb", X"e9", X"e0", X"ea", X"dc", X"de", X"d3", X"cf", X"d1", X"cf", X"d3", X"cb", X"ce", X"d0", X"cb", X"c8", X"c1", X"b8", X"ad", X"a2", X"95", X"91", X"7c", X"70", X"4e", X"39", X"22", X"2b", X"22", X"24", X"19", X"1e", X"1c", X"14", X"0f", X"10", X"13", X"08", X"06", X"0b", X"05", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"06", X"05", X"09", X"0d", X"13", X"16", X"19", X"2a", X"27", X"3d", X"5f", X"65", X"80", X"8b", X"85", X"90", X"87", X"93", X"9c", X"91", X"a2", X"9b", X"91", X"9f", X"aa", X"b2", X"b6", X"ba", X"c5", X"c5", X"ca", X"cc", X"cd", X"ce", X"d1", X"d1", X"d1", X"cf", X"e1", X"d5", X"da", X"de", X"d8", X"e1", X"e0", X"dc", X"e3", X"e4", X"e1", X"e9", X"e2", X"e1", X"e5", X"de", X"e3", X"e7", X"e4", X"e0", X"f0", X"ed", X"f0", X"f7", X"ef", X"ef", X"f1", X"ef", X"e7", X"e5", X"e1", X"de", X"e2", X"e1", X"e6", X"e8", X"f2", X"f4", X"fa", X"fa", X"f9", X"ef", X"f1", X"e9", X"dd", X"de", X"df", X"e1", X"df", X"db", X"dd", X"e3", X"de", X"e4", X"ec", X"e2", X"e5", X"e0", X"e3", X"ed", X"f7", X"f0", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"d7", X"d0", X"d1", X"cf", X"d8", X"cb", X"cc", X"ca", X"d4", X"d5", X"cf", X"d0", X"d3", X"d4", X"c6", X"c1", X"be", X"c2", X"c0", X"be", X"bf", X"bf", X"b3", X"b4", X"bd", X"b9", X"bc", X"ce", X"d2", X"d1", X"d7", X"d5", X"da", X"da", X"e3", X"e0", X"f1", X"f2", X"fd", X"ff", X"ff", X"fe", X"fc", X"ea", X"f4", X"f0", X"e8", X"eb", X"f5", X"f3", X"ea", X"ec", X"ef", X"eb", X"e6", X"e2", X"eb", X"eb", X"d8", X"df", X"db", X"d8", X"d0", X"d4", X"d3", X"c6", X"c8", X"c9", X"c6", X"bf", X"b7", X"b3", X"a1", X"9d", X"87", X"82", X"6f", X"64", X"47", X"2e", X"23", X"1e", X"1f", X"1e", X"1e", X"20", X"15", X"11", X"1f", X"10", X"13", X"09", X"07", X"06", X"03", X"10", X"0b", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"08", X"0d", X"0b", X"10", X"14", X"1c", X"1f", X"2b", X"38", X"4a", X"5a", X"6b", X"83", X"88", X"97", X"8f", X"9d", X"94", X"9a", X"a1", X"98", X"9f", X"a3", X"ac", X"ac", X"b1", X"b6", X"bb", X"c2", X"c2", X"c9", X"bd", X"d5", X"d3", X"cf", X"cf", X"cf", X"d6", X"d1", X"da", X"d0", X"dc", X"da", X"de", X"d4", X"e0", X"df", X"df", X"e3", X"e1", X"dc", X"dd", X"da", X"e3", X"e7", X"ec", X"e9", X"f3", X"f6", X"f3", X"f7", X"f0", X"e6", X"db", X"e4", X"df", X"db", X"d8", X"e7", X"e8", X"ef", X"ed", X"f9", X"fc", X"f7", X"fb", X"f7", X"f1", X"f7", X"ea", X"e6", X"e8", X"de", X"e2", X"df", X"da", X"e1", X"e4", X"e0", X"e4", X"e4", X"e7", X"e3", X"e4", X"ea", X"ec", X"ee", X"ef", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"d8", X"d7", X"ce", X"d1", X"cb", X"d0", X"ce", X"d7", X"cf", X"d4", X"d5", X"cf", X"cf", X"c6", X"c4", X"c9", X"c7", X"c2", X"bd", X"c2", X"be", X"c4", X"b8", X"af", X"b5", X"b8", X"ba", X"c4", X"cc", X"ca", X"cb", X"c9", X"d0", X"d0", X"cd", X"d8", X"e6", X"f0", X"f6", X"fb", X"f4", X"f2", X"fd", X"ee", X"f3", X"f3", X"e9", X"e6", X"ee", X"e9", X"ed", X"ef", X"e1", X"e3", X"e5", X"dc", X"e3", X"db", X"e2", X"d9", X"d2", X"d3", X"d2", X"cb", X"c8", X"ce", X"c5", X"b6", X"bf", X"b6", X"ae", X"ab", X"99", X"87", X"83", X"83", X"77", X"64", X"3e", X"35", X"29", X"25", X"23", X"24", X"1b", X"1d", X"19", X"15", X"0e", X"12", X"0e", X"12", X"06", X"08", X"08", X"00", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"0f", X"08", X"0e", X"16", X"20", X"23", X"2b", X"3e", X"50", X"62", X"7c", X"82", X"90", X"8d", X"8d", X"98", X"90", X"9a", X"97", X"a2", X"af", X"a8", X"b5", X"b3", X"b1", X"b9", X"b7", X"c8", X"c1", X"c5", X"cc", X"cb", X"c9", X"d2", X"d6", X"d8", X"d2", X"d7", X"d7", X"d4", X"cd", X"d6", X"d7", X"d5", X"d8", X"d5", X"dd", X"d7", X"cf", X"cd", X"d5", X"e0", X"e5", X"e7", X"e8", X"ec", X"f4", X"f7", X"e5", X"e5", X"e0", X"d7", X"d7", X"dc", X"dd", X"e0", X"e5", X"e9", X"eb", X"ee", X"f4", X"fa", X"f8", X"f8", X"fa", X"f2", X"ec", X"e6", X"e1", X"e3", X"e1", X"e2", X"d9", X"da", X"db", X"de", X"dd", X"e3", X"e2", X"e7", X"e5", X"e4", X"ee", X"de", X"e9", X"ec", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e1", X"d4", X"d5", X"cf", X"ca", X"c6", X"d5", X"d0", X"d0", X"d5", X"d8", X"cf", X"cf", X"ce", X"c8", X"cb", X"be", X"bc", X"bf", X"c0", X"bf", X"ba", X"b9", X"ac", X"ac", X"b6", X"b6", X"b8", X"bc", X"bd", X"c5", X"c6", X"c7", X"c7", X"cb", X"d1", X"d8", X"ea", X"eb", X"e7", X"f6", X"f6", X"ee", X"ef", X"ed", X"f4", X"e1", X"ee", X"e6", X"e2", X"e2", X"e5", X"e8", X"e3", X"e0", X"e2", X"dd", X"d9", X"d8", X"d2", X"d7", X"cf", X"c6", X"c2", X"c6", X"c0", X"cc", X"b9", X"b5", X"b1", X"a0", X"9f", X"91", X"8c", X"84", X"81", X"72", X"54", X"3d", X"31", X"2d", X"28", X"2e", X"1e", X"1b", X"1f", X"1a", X"19", X"0f", X"1b", X"12", X"0f", X"06", X"08", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0e", X"0d", X"0b", X"0d", X"0b", X"1a", X"21", X"25", X"3d", X"38", X"57", X"6f", X"79", X"8a", X"93", X"8a", X"8e", X"92", X"9e", X"9e", X"9f", X"a3", X"a1", X"b4", X"b7", X"b9", X"b5", X"ab", X"c2", X"be", X"ca", X"ce", X"d4", X"d1", X"ce", X"d1", X"da", X"d6", X"d8", X"ce", X"d3", X"d3", X"ce", X"e0", X"d6", X"cc", X"d1", X"d1", X"ce", X"cf", X"d4", X"d7", X"e2", X"e6", X"e8", X"ef", X"f8", X"ed", X"ef", X"e7", X"e0", X"dd", X"da", X"da", X"dd", X"df", X"dd", X"e8", X"f1", X"fa", X"ff", X"ff", X"ff", X"f9", X"fb", X"f3", X"f6", X"eb", X"e6", X"dc", X"e3", X"d8", X"d8", X"d9", X"dc", X"de", X"e2", X"d7", X"de", X"e0", X"e7", X"e4", X"e8", X"e4", X"eb", X"ea", X"f0", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ee", X"dc", X"ca", X"d4", X"c8", X"cc", X"d2", X"d2", X"d5", X"d0", X"d1", X"d1", X"ca", X"cc", X"be", X"c8", X"ca", X"c4", X"be", X"be", X"c2", X"ba", X"b5", X"b2", X"aa", X"b5", X"af", X"b0", X"b4", X"bf", X"c1", X"be", X"c8", X"bf", X"c9", X"cc", X"ce", X"d5", X"e6", X"de", X"f0", X"e5", X"ed", X"e8", X"ec", X"ed", X"e2", X"e5", X"e6", X"de", X"da", X"df", X"d7", X"e4", X"da", X"dc", X"d8", X"da", X"df", X"d8", X"d3", X"d5", X"cc", X"cc", X"c3", X"ba", X"be", X"ad", X"b2", X"9c", X"92", X"96", X"8e", X"8c", X"7d", X"83", X"6c", X"5b", X"3b", X"2f", X"2b", X"35", X"28", X"20", X"24", X"1c", X"10", X"12", X"15", X"0d", X"12", X"02", X"0a", X"05", X"0a", X"0a", X"06", X"0d", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"04", X"05", X"0a", X"10", X"0e", X"1d", X"1c", X"1c", X"2b", X"2f", X"3d", X"64", X"72", X"80", X"8d", X"8c", X"8c", X"93", X"96", X"9b", X"a1", X"a2", X"a3", X"ae", X"b4", X"b6", X"c3", X"c5", X"c8", X"c5", X"ce", X"c5", X"cc", X"d2", X"ca", X"c7", X"d7", X"ce", X"ce", X"d5", X"d6", X"c9", X"d9", X"d1", X"ce", X"c3", X"c7", X"c3", X"c8", X"cf", X"cd", X"e4", X"e7", X"eb", X"f2", X"f3", X"ee", X"ee", X"e9", X"df", X"e2", X"db", X"da", X"d5", X"d8", X"e1", X"f0", X"f5", X"fb", X"ff", X"fc", X"fa", X"ff", X"f5", X"fb", X"f1", X"f2", X"eb", X"db", X"e0", X"e1", X"d6", X"dd", X"de", X"d8", X"db", X"db", X"da", X"e0", X"e0", X"e2", X"e9", X"e5", X"e6", X"e9", X"e6", X"fa", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fe", X"d9", X"c9", X"d2", X"c9", X"d1", X"d3", X"cc", X"ca", X"cb", X"d0", X"da", X"d2", X"ce", X"c2", X"c1", X"c0", X"bc", X"be", X"bd", X"b5", X"b5", X"b9", X"aa", X"a6", X"af", X"b3", X"b9", X"b5", X"b9", X"b9", X"be", X"bc", X"b9", X"c3", X"c5", X"ce", X"d2", X"d2", X"da", X"dd", X"df", X"e1", X"db", X"e7", X"e1", X"dc", X"e5", X"da", X"de", X"e0", X"d2", X"dd", X"d4", X"d7", X"d6", X"dd", X"dd", X"cf", X"d7", X"cf", X"cd", X"c9", X"c0", X"c3", X"c4", X"b9", X"b1", X"a4", X"9e", X"89", X"90", X"89", X"8e", X"8f", X"73", X"6b", X"4f", X"34", X"2f", X"2c", X"32", X"2d", X"2a", X"25", X"2c", X"12", X"14", X"14", X"0b", X"07", X"14", X"07", X"10", X"03", X"00", X"0a", X"05", X"04", X"09", X"06", X"05", X"05", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0b", X"09", X"06", X"08", X"05", X"0d", X"0f", X"16", X"18", X"26", X"2c", X"37", X"4d", X"6e", X"71", X"82", X"83", X"8f", X"95", X"92", X"8d", X"98", X"a1", X"a3", X"a5", X"aa", X"af", X"b6", X"c0", X"bf", X"cb", X"cd", X"c7", X"cd", X"c9", X"cb", X"ca", X"d2", X"d0", X"cd", X"d3", X"d5", X"ce", X"c8", X"c6", X"c5", X"c6", X"c4", X"c7", X"c5", X"d6", X"d5", X"df", X"e9", X"ec", X"ea", X"eb", X"e9", X"e1", X"e5", X"e6", X"e1", X"d8", X"cf", X"de", X"e1", X"e9", X"f2", X"f6", X"f8", X"fd", X"f8", X"f4", X"f4", X"f6", X"fb", X"f1", X"f0", X"eb", X"e1", X"e2", X"e5", X"e0", X"e0", X"d6", X"da", X"e2", X"da", X"de", X"d8", X"db", X"e2", X"e1", X"e5", X"e3", X"e1", X"e6", X"ea", X"fe", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"df", X"cd", X"d2", X"d1", X"d4", X"d1", X"d9", X"cc", X"c4", X"cd", X"c2", X"ca", X"c9", X"c0", X"ca", X"bd", X"ba", X"bf", X"b4", X"b2", X"b8", X"af", X"a6", X"aa", X"b1", X"a6", X"ae", X"b8", X"b1", X"b6", X"b3", X"ba", X"ae", X"b9", X"bf", X"bc", X"c3", X"c2", X"cf", X"cb", X"d9", X"df", X"da", X"e4", X"de", X"d6", X"de", X"d4", X"d7", X"d2", X"d0", X"d2", X"d0", X"d4", X"d6", X"d9", X"cf", X"d3", X"d7", X"d2", X"c8", X"c0", X"bd", X"b9", X"af", X"a9", X"a1", X"95", X"99", X"91", X"91", X"8a", X"88", X"79", X"77", X"64", X"43", X"2d", X"26", X"27", X"30", X"28", X"2d", X"1e", X"1c", X"14", X"12", X"17", X"15", X"0f", X"0b", X"09", X"0b", X"03", X"01", X"0c", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"0c", X"11", X"08", X"0d", X"16", X"16", X"1b", X"1b", X"28", X"32", X"3f", X"5b", X"78", X"7b", X"84", X"8e", X"8e", X"92", X"91", X"8e", X"98", X"9b", X"a8", X"aa", X"b1", X"b2", X"b7", X"ba", X"be", X"c9", X"c1", X"ca", X"c5", X"c9", X"cf", X"c8", X"ca", X"c8", X"d0", X"ca", X"ca", X"c2", X"c3", X"c8", X"c7", X"cf", X"c8", X"d9", X"d9", X"d5", X"ec", X"e8", X"ea", X"f2", X"ea", X"ec", X"ea", X"e7", X"db", X"d9", X"d5", X"db", X"e9", X"e6", X"ef", X"fb", X"fc", X"ff", X"fb", X"f6", X"f7", X"f4", X"ec", X"f0", X"ea", X"e7", X"e3", X"e2", X"dc", X"e6", X"e0", X"d5", X"dd", X"d3", X"db", X"de", X"d9", X"dc", X"e4", X"e6", X"da", X"e4", X"df", X"e2", X"ec", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"de", X"d0", X"cf", X"d3", X"d3", X"d0", X"cd", X"d3", X"cd", X"ce", X"c6", X"c1", X"c9", X"c1", X"c7", X"c0", X"c3", X"be", X"c2", X"b0", X"c3", X"b4", X"aa", X"a9", X"a4", X"aa", X"aa", X"a4", X"a8", X"a8", X"aa", X"ba", X"ac", X"ac", X"b0", X"b4", X"bb", X"c0", X"c9", X"c3", X"d3", X"cd", X"d2", X"db", X"d8", X"d4", X"d4", X"d3", X"ce", X"c9", X"c7", X"d0", X"ce", X"cb", X"cf", X"cd", X"c8", X"cb", X"d0", X"c6", X"c7", X"be", X"b7", X"ae", X"aa", X"a2", X"9a", X"96", X"94", X"87", X"8e", X"88", X"7d", X"7d", X"6b", X"52", X"44", X"35", X"2d", X"2d", X"34", X"26", X"2a", X"25", X"24", X"1d", X"19", X"12", X"11", X"0f", X"05", X"06", X"09", X"0a", X"09", X"06", X"0c", X"03", X"0b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"09", X"0a", X"0b", X"0a", X"0d", X"0c", X"1c", X"27", X"26", X"29", X"3b", X"4e", X"70", X"7e", X"84", X"84", X"90", X"8f", X"89", X"8b", X"9c", X"9e", X"a3", X"a4", X"a9", X"a7", X"aa", X"b1", X"ba", X"c3", X"c5", X"c1", X"c2", X"c7", X"cc", X"cf", X"c6", X"c7", X"cb", X"c9", X"c3", X"b9", X"be", X"c4", X"cd", X"d6", X"cf", X"dd", X"e1", X"ea", X"e9", X"e8", X"e7", X"e9", X"e4", X"e6", X"ee", X"df", X"d7", X"d5", X"d9", X"e1", X"e4", X"ee", X"f3", X"fc", X"ff", X"fa", X"f9", X"fa", X"f9", X"f7", X"eb", X"e3", X"e7", X"e7", X"df", X"e9", X"e2", X"dd", X"da", X"d8", X"d3", X"db", X"da", X"dc", X"db", X"e0", X"dc", X"e2", X"e2", X"d9", X"de", X"dc", X"e8", X"f8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e4", X"d4", X"d9", X"ce", X"d6", X"d3", X"d0", X"d2", X"c5", X"c8", X"ca", X"be", X"c4", X"c9", X"c1", X"c7", X"be", X"bd", X"be", X"ad", X"b4", X"b0", X"a6", X"a4", X"a5", X"a4", X"a5", X"ad", X"a3", X"ac", X"a3", X"aa", X"a6", X"a9", X"ab", X"ab", X"b7", X"b6", X"af", X"c2", X"c2", X"cc", X"ca", X"c6", X"cf", X"ca", X"ce", X"c8", X"cb", X"b9", X"c1", X"c4", X"bd", X"b9", X"c3", X"bc", X"c4", X"be", X"bb", X"b8", X"b5", X"b9", X"a9", X"a7", X"98", X"96", X"92", X"94", X"8d", X"8e", X"89", X"81", X"7f", X"77", X"6d", X"51", X"43", X"34", X"35", X"32", X"34", X"2b", X"2a", X"26", X"1c", X"15", X"1d", X"1a", X"17", X"0e", X"0f", X"09", X"12", X"09", X"11", X"06", X"0e", X"12", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"04", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"0d", X"0a", X"09", X"0a", X"07", X"0e", X"0d", X"19", X"1e", X"28", X"29", X"2f", X"46", X"64", X"7f", X"80", X"85", X"90", X"8b", X"93", X"92", X"8d", X"94", X"a3", X"9e", X"a7", X"af", X"b1", X"b4", X"b3", X"b4", X"b8", X"cb", X"c1", X"cc", X"c8", X"ce", X"be", X"c8", X"c5", X"c6", X"ce", X"cc", X"ca", X"ce", X"cf", X"d4", X"e3", X"e3", X"e9", X"ea", X"e8", X"e9", X"e5", X"e6", X"e4", X"f1", X"e8", X"d8", X"de", X"d6", X"d8", X"e2", X"eb", X"f0", X"f8", X"fd", X"ff", X"fb", X"f9", X"f6", X"ea", X"eb", X"e8", X"ee", X"e1", X"d9", X"e1", X"e0", X"df", X"e0", X"d8", X"da", X"d1", X"d6", X"d6", X"da", X"d2", X"dc", X"de", X"e4", X"dd", X"e2", X"e1", X"e4", X"e7", X"f8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f2", X"da", X"db", X"cc", X"c7", X"cb", X"ce", X"c8", X"c5", X"c9", X"cc", X"ba", X"bf", X"c6", X"bd", X"b6", X"b9", X"b3", X"bb", X"b4", X"b2", X"aa", X"aa", X"9f", X"a8", X"9f", X"a6", X"a0", X"a5", X"a5", X"a5", X"a2", X"a4", X"9f", X"a0", X"a0", X"a5", X"a9", X"b1", X"b2", X"b3", X"bc", X"bc", X"bb", X"c0", X"b9", X"be", X"b9", X"b7", X"b0", X"af", X"b3", X"b7", X"b2", X"b9", X"b0", X"bd", X"b5", X"b4", X"b8", X"b4", X"a3", X"9f", X"9a", X"97", X"92", X"96", X"94", X"95", X"8d", X"87", X"80", X"76", X"6e", X"62", X"54", X"40", X"34", X"39", X"34", X"35", X"31", X"22", X"23", X"22", X"1b", X"17", X"08", X"0c", X"11", X"0e", X"09", X"0f", X"03", X"09", X"06", X"10", X"04", X"05", X"06", X"05", X"08", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"09", X"0a", X"09", X"0f", X"15", X"18", X"1b", X"1b", X"22", X"2e", X"36", X"4a", X"5f", X"7b", X"84", X"84", X"88", X"88", X"8a", X"96", X"93", X"a0", X"a2", X"a8", X"a5", X"b4", X"af", X"ae", X"b9", X"bd", X"b9", X"c0", X"c5", X"c9", X"cd", X"c5", X"d0", X"c1", X"c7", X"c8", X"cc", X"c9", X"cf", X"cf", X"d8", X"db", X"e0", X"e0", X"e1", X"e6", X"e6", X"ea", X"e2", X"de", X"e1", X"e5", X"e2", X"d5", X"d8", X"d7", X"d2", X"da", X"ec", X"f1", X"f4", X"f4", X"f6", X"f8", X"f2", X"ee", X"e9", X"e9", X"e5", X"e0", X"e4", X"dd", X"e4", X"e2", X"d5", X"db", X"d8", X"de", X"d5", X"d2", X"d3", X"c9", X"d2", X"df", X"d5", X"de", X"d8", X"dc", X"dc", X"e6", X"e2", X"f1", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ef", X"f8", X"fb", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f6", X"d2", X"c7", X"c2", X"cb", X"c7", X"c8", X"c6", X"c7", X"c0", X"ba", X"c0", X"b9", X"b9", X"bb", X"be", X"b5", X"bb", X"b8", X"a5", X"ab", X"aa", X"a2", X"a1", X"a3", X"9f", X"a8", X"a0", X"a1", X"9b", X"9a", X"9f", X"a6", X"a0", X"a2", X"9c", X"a1", X"a9", X"a5", X"a8", X"a5", X"b1", X"b2", X"ae", X"b5", X"b2", X"ad", X"ac", X"ac", X"ae", X"a9", X"ab", X"a7", X"a9", X"a5", X"ab", X"aa", X"aa", X"ad", X"b1", X"a7", X"9d", X"96", X"9e", X"93", X"98", X"8b", X"85", X"84", X"7d", X"83", X"77", X"73", X"68", X"62", X"54", X"41", X"33", X"3a", X"37", X"37", X"35", X"2b", X"29", X"23", X"1d", X"1a", X"1a", X"0f", X"13", X"0b", X"0d", X"05", X"0e", X"07", X"0c", X"0d", X"07", X"00", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"00", X"06", X"09", X"07", X"09", X"08", X"05", X"08", X"10", X"19", X"1b", X"1f", X"20", X"25", X"2e", X"46", X"59", X"75", X"83", X"88", X"90", X"8d", X"93", X"8c", X"96", X"97", X"a3", X"a5", X"a4", X"ab", X"ae", X"b2", X"b8", X"be", X"bc", X"bd", X"c2", X"cc", X"c3", X"d3", X"c5", X"c6", X"c6", X"cd", X"c7", X"cc", X"d0", X"d5", X"d2", X"d2", X"dd", X"dd", X"e0", X"da", X"db", X"d5", X"da", X"e0", X"e6", X"da", X"d6", X"d5", X"d9", X"db", X"e0", X"de", X"ec", X"ee", X"f0", X"f7", X"fb", X"fa", X"f6", X"e1", X"ed", X"eb", X"e7", X"e7", X"e6", X"e0", X"df", X"d6", X"d9", X"d9", X"da", X"d6", X"d8", X"d6", X"d1", X"d6", X"d7", X"d4", X"dc", X"e0", X"e1", X"dc", X"db", X"e7", X"e3", X"f6", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e3", X"dd", X"cf", X"c7", X"cf", X"e2", X"e3", X"e4", X"f7", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"d0", X"c1", X"c6", X"c2", X"c2", X"cc", X"c2", X"c6", X"c0", X"c7", X"b9", X"be", X"b9", X"b6", X"ba", X"b2", X"b8", X"b4", X"ad", X"af", X"a6", X"a0", X"a3", X"a2", X"9d", X"a7", X"9b", X"a2", X"a0", X"a4", X"a0", X"a1", X"a3", X"9e", X"98", X"a3", X"98", X"a1", X"a6", X"9f", X"af", X"a5", X"a3", X"ab", X"ab", X"a7", X"a6", X"a9", X"a4", X"a5", X"a9", X"9f", X"a8", X"9f", X"9e", X"a3", X"a3", X"a0", X"a3", X"94", X"9b", X"97", X"9c", X"90", X"92", X"89", X"89", X"84", X"81", X"7e", X"7d", X"6b", X"63", X"60", X"48", X"48", X"45", X"4b", X"3c", X"2c", X"35", X"2e", X"2e", X"25", X"1e", X"1c", X"13", X"11", X"18", X"09", X"07", X"10", X"0c", X"07", X"11", X"13", X"08", X"04", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"01", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"0f", X"0e", X"09", X"0e", X"0c", X"13", X"13", X"1c", X"27", X"21", X"27", X"3a", X"52", X"73", X"82", X"88", X"85", X"87", X"94", X"91", X"92", X"9f", X"9b", X"a0", X"9b", X"a5", X"ab", X"a6", X"ae", X"ba", X"c0", X"c3", X"c1", X"c9", X"cd", X"d1", X"c6", X"cc", X"c5", X"c6", X"cf", X"c5", X"c8", X"d0", X"d1", X"d3", X"d3", X"d7", X"d9", X"d4", X"d3", X"ce", X"d5", X"d7", X"dd", X"db", X"d7", X"d3", X"d8", X"df", X"dd", X"e4", X"eb", X"f5", X"f0", X"ef", X"f2", X"f0", X"f0", X"e5", X"e3", X"e1", X"e0", X"e1", X"e3", X"d6", X"da", X"d8", X"d2", X"db", X"d3", X"d3", X"d8", X"d2", X"d8", X"d9", X"d6", X"d3", X"d6", X"dd", X"d5", X"db", X"de", X"dc", X"da", X"f4", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"f5", X"e6", X"e8", X"e0", X"dd", X"e4", X"dc", X"d4", X"c4", X"b5", X"b3", X"ad", X"b5", X"b0", X"b8", X"be", X"d0", X"e8", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ce", X"c5", X"b4", X"bd", X"bc", X"c2", X"c3", X"ba", X"b9", X"b6", X"b3", X"b8", X"b1", X"b2", X"b0", X"b1", X"b3", X"ae", X"aa", X"a5", X"a1", X"ad", X"a2", X"a2", X"a0", X"a2", X"97", X"98", X"9a", X"9d", X"97", X"9a", X"97", X"9f", X"a0", X"9e", X"9c", X"97", X"97", X"9f", X"ab", X"99", X"a4", X"a6", X"a0", X"a2", X"a7", X"a2", X"a1", X"a5", X"9c", X"a5", X"a1", X"9d", X"9a", X"9b", X"a2", X"97", X"a0", X"98", X"8f", X"8c", X"87", X"84", X"88", X"7d", X"7e", X"7d", X"73", X"7c", X"6d", X"65", X"66", X"5d", X"55", X"55", X"46", X"53", X"4d", X"3b", X"35", X"2a", X"26", X"21", X"1d", X"1e", X"14", X"19", X"09", X"18", X"0a", X"09", X"0d", X"10", X"09", X"07", X"0a", X"04", X"06", X"05", X"04", X"05", X"07", X"0b", X"03", X"08", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"05", X"02", X"0a", X"05", X"09", X"11", X"13", X"16", X"1c", X"1f", X"25", X"2d", X"34", X"3f", X"6b", X"8a", X"85", X"8f", X"94", X"8c", X"99", X"8f", X"9a", X"97", X"95", X"9e", X"9a", X"a5", X"ac", X"ad", X"ad", X"bb", X"ba", X"bd", X"c5", X"c5", X"cb", X"c8", X"c1", X"c5", X"c5", X"be", X"c4", X"c6", X"c6", X"cc", X"c8", X"c7", X"c8", X"c4", X"cf", X"ca", X"cd", X"d5", X"d4", X"d2", X"d3", X"d9", X"ce", X"c9", X"d5", X"da", X"d7", X"e0", X"e5", X"e1", X"ec", X"e4", X"e3", X"e2", X"e2", X"dc", X"dd", X"db", X"df", X"df", X"d9", X"d7", X"d2", X"d5", X"cc", X"cf", X"ce", X"cc", X"d7", X"d4", X"cc", X"c3", X"d2", X"d0", X"d8", X"d2", X"db", X"d8", X"d7", X"dd", X"f2", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"e0", X"c4", X"bf", X"c2", X"b0", X"bc", X"b2", X"b8", X"aa", X"a7", X"a7", X"a3", X"96", X"94", X"8a", X"93", X"94", X"9e", X"a2", X"a9", X"b8", X"cf", X"db", X"f3", X"ff", X"ff", X"ff", X"ff", X"ff", X"fb", X"c2", X"be", X"b5", X"bb", X"c0", X"be", X"b8", X"b2", X"b5", X"b1", X"b1", X"ac", X"ad", X"a7", X"aa", X"b2", X"aa", X"a9", X"9b", X"9e", X"9f", X"9f", X"a5", X"9c", X"9a", X"9e", X"97", X"93", X"93", X"99", X"90", X"99", X"91", X"98", X"95", X"99", X"9c", X"9b", X"9c", X"92", X"a1", X"9b", X"a0", X"a7", X"99", X"a4", X"a3", X"9d", X"a2", X"9f", X"96", X"9e", X"9a", X"97", X"97", X"95", X"9a", X"8e", X"8e", X"90", X"8c", X"85", X"83", X"82", X"7f", X"77", X"76", X"75", X"73", X"73", X"75", X"65", X"67", X"5f", X"52", X"55", X"5a", X"4e", X"41", X"35", X"31", X"23", X"1c", X"1e", X"19", X"0f", X"10", X"13", X"0d", X"07", X"0a", X"0b", X"0e", X"09", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"06", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"06", X"08", X"07", X"0d", X"0e", X"07", X"0c", X"11", X"1a", X"1c", X"25", X"25", X"27", X"3b", X"47", X"60", X"86", X"96", X"94", X"99", X"9f", X"9e", X"a0", X"a1", X"94", X"9b", X"9d", X"a1", X"a4", X"a8", X"a6", X"b1", X"b4", X"bd", X"c2", X"be", X"c7", X"cb", X"c1", X"c3", X"c2", X"c0", X"bf", X"c4", X"c1", X"c4", X"c1", X"be", X"c6", X"c3", X"c1", X"cc", X"cb", X"c9", X"d3", X"d6", X"cb", X"d1", X"c5", X"ce", X"c7", X"d0", X"d4", X"d5", X"dc", X"e4", X"df", X"e5", X"e4", X"d8", X"e0", X"df", X"d9", X"e6", X"d9", X"da", X"da", X"d9", X"d6", X"ca", X"cf", X"ce", X"c8", X"c2", X"c7", X"c7", X"d0", X"c7", X"ca", X"d0", X"c6", X"d2", X"d3", X"d1", X"cf", X"d7", X"d9", X"f2", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ee", X"d7", X"bf", X"af", X"9c", X"9b", X"96", X"94", X"95", X"8d", X"8e", X"7e", X"77", X"7b", X"79", X"78", X"84", X"78", X"7d", X"85", X"85", X"88", X"8e", X"96", X"a4", X"ae", X"bd", X"d5", X"e9", X"ff", X"ff", X"ff", X"fb", X"bd", X"b9", X"b1", X"c0", X"ba", X"b7", X"bf", X"b5", X"ae", X"b1", X"ad", X"ac", X"a7", X"ab", X"a6", X"a1", X"a2", X"a9", X"a3", X"9f", X"9c", X"a1", X"a5", X"99", X"94", X"a0", X"99", X"9b", X"98", X"9a", X"9d", X"97", X"90", X"94", X"98", X"99", X"90", X"94", X"96", X"95", X"94", X"a0", X"a2", X"a5", X"a1", X"a3", X"98", X"9b", X"a4", X"9f", X"96", X"9d", X"96", X"94", X"92", X"8f", X"96", X"8c", X"8e", X"89", X"84", X"7a", X"81", X"71", X"7a", X"75", X"7a", X"7f", X"75", X"78", X"66", X"64", X"5d", X"60", X"58", X"60", X"5f", X"55", X"44", X"3a", X"2f", X"2a", X"1f", X"1e", X"19", X"11", X"0f", X"12", X"12", X"0e", X"07", X"09", X"09", X"07", X"0a", X"11", X"03", X"09", X"06", X"05", X"03", X"0a", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"12", X"05", X"03", X"14", X"0d", X"0b", X"13", X"14", X"12", X"23", X"26", X"22", X"2c", X"32", X"44", X"5b", X"80", X"92", X"91", X"9e", X"9a", X"a2", X"a6", X"9c", X"9d", X"a2", X"a0", X"9e", X"a9", X"a3", X"a7", X"aa", X"af", X"be", X"bf", X"c0", X"c5", X"c1", X"c5", X"bf", X"b6", X"bb", X"c0", X"b9", X"bd", X"bc", X"c5", X"bd", X"c5", X"bd", X"b7", X"c7", X"c9", X"c2", X"c3", X"c5", X"c4", X"ca", X"c9", X"c3", X"ca", X"cc", X"cd", X"d5", X"d4", X"d7", X"de", X"d9", X"df", X"d0", X"db", X"df", X"d4", X"da", X"da", X"dc", X"dc", X"dc", X"d8", X"d8", X"d2", X"cd", X"c9", X"ce", X"ca", X"c8", X"c5", X"ce", X"c9", X"cb", X"d3", X"ce", X"d0", X"d1", X"d1", X"d1", X"d7", X"ee", X"ff", X"ff", X"ff", X"ff", X"ee", X"d2", X"b4", X"a1", X"90", X"87", X"80", X"76", X"76", X"6e", X"70", X"6f", X"69", X"5e", X"60", X"5f", X"60", X"60", X"61", X"62", X"61", X"67", X"67", X"75", X"7d", X"83", X"8d", X"8f", X"9f", X"b7", X"c0", X"dc", X"ff", X"ff", X"f9", X"bd", X"ac", X"a9", X"b7", X"b8", X"b1", X"bb", X"aa", X"ab", X"ab", X"a0", X"a5", X"a2", X"a6", X"a9", X"a5", X"a0", X"9b", X"9f", X"a0", X"97", X"98", X"94", X"9a", X"93", X"99", X"96", X"91", X"97", X"92", X"99", X"99", X"95", X"96", X"96", X"96", X"94", X"94", X"93", X"98", X"9e", X"9b", X"99", X"a0", X"9e", X"9f", X"a4", X"97", X"9e", X"94", X"93", X"97", X"92", X"90", X"91", X"8e", X"8f", X"87", X"86", X"8a", X"77", X"70", X"76", X"75", X"75", X"6f", X"73", X"7b", X"76", X"72", X"71", X"6b", X"68", X"5f", X"5e", X"64", X"5d", X"55", X"4e", X"44", X"2d", X"2b", X"28", X"21", X"20", X"1e", X"0c", X"10", X"14", X"10", X"08", X"0d", X"0a", X"0b", X"06", X"05", X"07", X"02", X"06", X"05", X"08", X"04", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"07", X"06", X"05", X"0b", X"14", X"0d", X"15", X"1d", X"21", X"28", X"28", X"37", X"41", X"61", X"7d", X"88", X"93", X"9a", X"99", X"a8", X"a5", X"a5", X"ac", X"ab", X"a1", X"a0", X"a3", X"a7", X"aa", X"ab", X"b0", X"c0", X"b8", X"c4", X"bc", X"ba", X"c1", X"ba", X"c0", X"c0", X"bd", X"c0", X"bf", X"c1", X"b6", X"bc", X"bf", X"b9", X"bb", X"bf", X"bf", X"bb", X"c4", X"c0", X"c3", X"bc", X"bf", X"c4", X"c2", X"bf", X"cd", X"ce", X"ce", X"cc", X"d2", X"d6", X"d3", X"cf", X"d1", X"d7", X"d4", X"da", X"cf", X"ce", X"d4", X"d2", X"d5", X"cc", X"ce", X"c6", X"ca", X"cb", X"c7", X"ca", X"c5", X"ca", X"b9", X"ca", X"ce", X"c4", X"cd", X"c9", X"ce", X"d4", X"d0", X"e1", X"ff", X"ff", X"f5", X"d0", X"b0", X"a7", X"96", X"8a", X"7c", X"6d", X"64", X"64", X"5d", X"59", X"54", X"58", X"55", X"54", X"52", X"4d", X"50", X"50", X"56", X"45", X"50", X"54", X"4f", X"5a", X"61", X"63", X"72", X"80", X"8a", X"96", X"aa", X"bd", X"ee", X"ff", X"ea", X"b5", X"ae", X"a8", X"ac", X"ad", X"ae", X"b5", X"b5", X"aa", X"a3", X"a1", X"97", X"9b", X"98", X"95", X"97", X"9f", X"98", X"95", X"9b", X"98", X"94", X"95", X"98", X"9a", X"95", X"97", X"94", X"94", X"95", X"93", X"8d", X"8d", X"8c", X"91", X"94", X"92", X"8e", X"99", X"99", X"95", X"93", X"97", X"95", X"90", X"98", X"97", X"91", X"a1", X"98", X"8b", X"92", X"8c", X"8d", X"86", X"86", X"89", X"7c", X"79", X"76", X"6e", X"70", X"69", X"6b", X"74", X"71", X"73", X"78", X"6c", X"6d", X"70", X"66", X"6f", X"61", X"63", X"68", X"58", X"5c", X"40", X"3e", X"36", X"2e", X"26", X"16", X"1f", X"1c", X"13", X"0a", X"13", X"0c", X"09", X"05", X"04", X"06", X"08", X"0c", X"0d", X"06", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"0c", X"0b", X"06", X"0c", X"10", X"12", X"10", X"17", X"20", X"28", X"33", X"2e", X"39", X"43", X"51", X"77", X"85", X"88", X"94", X"90", X"9e", X"a4", X"a6", X"ac", X"b3", X"ab", X"ab", X"b2", X"a8", X"b1", X"b9", X"b4", X"b9", X"bb", X"c3", X"c1", X"bf", X"be", X"c1", X"bf", X"bf", X"b9", X"c0", X"be", X"b7", X"b9", X"b3", X"b8", X"c1", X"b6", X"bb", X"b7", X"b6", X"bd", X"c0", X"ba", X"b8", X"b5", X"b7", X"c2", X"c7", X"c6", X"c4", X"c4", X"cd", X"d0", X"ca", X"ce", X"c6", X"c4", X"c9", X"c3", X"cd", X"cb", X"c6", X"d1", X"cb", X"d3", X"cd", X"c4", X"c7", X"ce", X"ca", X"ca", X"be", X"bf", X"be", X"c2", X"bc", X"c3", X"c7", X"c5", X"cb", X"c8", X"ba", X"c4", X"d5", X"ea", X"d5", X"bc", X"b1", X"9f", X"97", X"83", X"72", X"69", X"60", X"51", X"52", X"46", X"4b", X"45", X"3e", X"3d", X"3f", X"40", X"32", X"45", X"3f", X"44", X"47", X"43", X"41", X"48", X"4e", X"5c", X"60", X"5f", X"67", X"74", X"80", X"93", X"b2", X"e0", X"ff", X"e0", X"b3", X"a7", X"a4", X"aa", X"ab", X"b6", X"ac", X"a9", X"a6", X"a2", X"9d", X"a4", X"9c", X"9f", X"9a", X"99", X"9c", X"98", X"97", X"94", X"90", X"9c", X"8f", X"94", X"92", X"94", X"8b", X"96", X"9b", X"94", X"92", X"91", X"86", X"8a", X"8f", X"8b", X"95", X"8a", X"84", X"99", X"98", X"90", X"9f", X"94", X"94", X"90", X"97", X"9a", X"90", X"93", X"8f", X"86", X"88", X"87", X"84", X"7d", X"7b", X"68", X"6d", X"72", X"65", X"6c", X"6c", X"62", X"6b", X"64", X"6f", X"75", X"70", X"71", X"6c", X"6b", X"6c", X"61", X"5f", X"65", X"5c", X"51", X"4e", X"3b", X"37", X"26", X"1e", X"27", X"17", X"15", X"11", X"14", X"16", X"09", X"0b", X"08", X"06", X"0c", X"0d", X"08", X"11", X"06", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"07", X"0b", X"0e", X"07", X"0f", X"11", X"17", X"1a", X"2a", X"34", X"39", X"31", X"3b", X"42", X"51", X"6d", X"84", X"89", X"90", X"9b", X"9e", X"a6", X"9e", X"a5", X"a5", X"ad", X"b3", X"b6", X"b8", X"b6", X"b8", X"b9", X"c2", X"be", X"c2", X"c0", X"c3", X"bf", X"be", X"be", X"be", X"bd", X"ba", X"bc", X"b8", X"be", X"b6", X"b2", X"b4", X"ab", X"b2", X"b6", X"b3", X"b4", X"b6", X"b3", X"ab", X"b1", X"bb", X"ac", X"b8", X"be", X"b5", X"c8", X"c7", X"c4", X"c0", X"cb", X"c6", X"c6", X"c6", X"c4", X"cb", X"c6", X"cc", X"ca", X"c2", X"c6", X"c6", X"cc", X"c2", X"b9", X"c0", X"bb", X"c3", X"c3", X"bc", X"b4", X"be", X"bb", X"be", X"bc", X"bf", X"bd", X"ba", X"b9", X"c7", X"d3", X"ba", X"99", X"8a", X"89", X"81", X"6f", X"5d", X"53", X"49", X"3e", X"43", X"37", X"3c", X"39", X"33", X"34", X"32", X"3b", X"36", X"32", X"35", X"3b", X"30", X"40", X"3d", X"45", X"40", X"4b", X"4d", X"52", X"55", X"60", X"6f", X"8a", X"9c", X"c1", X"ed", X"d2", X"b0", X"ab", X"a9", X"b1", X"ad", X"a7", X"af", X"a0", X"a3", X"a9", X"a0", X"98", X"97", X"99", X"9d", X"91", X"94", X"90", X"91", X"9a", X"94", X"99", X"9b", X"9c", X"8a", X"98", X"8c", X"85", X"8c", X"8e", X"8a", X"92", X"8b", X"92", X"8d", X"91", X"90", X"91", X"93", X"91", X"9a", X"93", X"94", X"95", X"95", X"93", X"96", X"90", X"8f", X"8f", X"89", X"88", X"80", X"78", X"7d", X"71", X"74", X"75", X"6e", X"77", X"68", X"61", X"64", X"69", X"61", X"6f", X"6b", X"71", X"70", X"74", X"6e", X"75", X"69", X"61", X"5d", X"69", X"5b", X"56", X"4c", X"34", X"30", X"2d", X"1d", X"1f", X"22", X"16", X"12", X"11", X"0f", X"08", X"07", X"09", X"09", X"0f", X"09", X"08", X"03", X"05", X"0a", X"05", X"03", X"04", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"06", X"09", X"05", X"10", X"06", X"0d", X"0e", X"14", X"24", X"2e", X"36", X"3b", X"3f", X"37", X"3e", X"51", X"68", X"84", X"8b", X"85", X"8e", X"98", X"a0", X"a1", X"a2", X"a3", X"ae", X"b6", X"b9", X"b8", X"b5", X"c0", X"b2", X"c5", X"c2", X"bb", X"c3", X"c4", X"c1", X"c4", X"bf", X"ba", X"bc", X"b5", X"b0", X"b1", X"b1", X"af", X"af", X"b6", X"b0", X"ac", X"ab", X"b4", X"ac", X"b2", X"ad", X"b6", X"b5", X"ab", X"b1", X"af", X"b0", X"b1", X"b3", X"b2", X"b1", X"b8", X"c5", X"bf", X"be", X"c2", X"bc", X"bc", X"bd", X"bd", X"cc", X"c3", X"ba", X"c4", X"c3", X"bc", X"bf", X"c2", X"b9", X"b6", X"b8", X"b7", X"b2", X"b4", X"b8", X"b4", X"ba", X"ae", X"b6", X"b7", X"b6", X"b5", X"b9", X"b7", X"86", X"84", X"72", X"65", X"54", X"53", X"46", X"3f", X"39", X"3c", X"38", X"2f", X"30", X"2a", X"2c", X"26", X"2a", X"29", X"2f", X"2c", X"2e", X"2a", X"2f", X"30", X"37", X"3d", X"31", X"3a", X"3f", X"49", X"54", X"60", X"6b", X"8c", X"a0", X"cf", X"c2", X"aa", X"a3", X"a8", X"a5", X"a6", X"a0", X"a5", X"a9", X"9f", X"9e", X"96", X"90", X"97", X"8d", X"98", X"8e", X"8d", X"96", X"92", X"8d", X"91", X"94", X"8f", X"91", X"94", X"92", X"92", X"8a", X"8b", X"8f", X"8b", X"8e", X"8f", X"8e", X"88", X"8d", X"8a", X"8e", X"9d", X"92", X"98", X"8f", X"90", X"94", X"91", X"91", X"95", X"8b", X"8b", X"89", X"84", X"84", X"7b", X"73", X"74", X"6f", X"67", X"6d", X"60", X"60", X"60", X"60", X"66", X"52", X"5d", X"5e", X"69", X"6a", X"6a", X"70", X"71", X"67", X"62", X"5d", X"5f", X"65", X"5f", X"52", X"4b", X"3d", X"34", X"30", X"29", X"1d", X"12", X"10", X"12", X"0b", X"0f", X"0a", X"08", X"06", X"03", X"02", X"09", X"05", X"04", X"02", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"08", X"08", X"0f", X"0b", X"05", X"0a", X"11", X"12", X"19", X"1d", X"21", X"2c", X"39", X"42", X"46", X"3e", X"47", X"4e", X"65", X"77", X"88", X"80", X"84", X"84", X"92", X"98", X"9b", X"a0", X"a2", X"a9", X"b3", X"b5", X"be", X"cd", X"c5", X"c6", X"c1", X"c4", X"bf", X"c4", X"c1", X"ba", X"bd", X"ba", X"b3", X"b0", X"b8", X"b0", X"ae", X"ad", X"b3", X"b2", X"b3", X"a5", X"b0", X"a3", X"a8", X"ac", X"a6", X"b0", X"ad", X"a5", X"a7", X"b2", X"af", X"b0", X"ac", X"b8", X"b0", X"b4", X"b4", X"ba", X"b4", X"bb", X"b9", X"b7", X"b6", X"bd", X"b7", X"c1", X"c1", X"b7", X"c0", X"b5", X"ad", X"b8", X"b4", X"b1", X"b3", X"b8", X"b1", X"b0", X"b1", X"ae", X"af", X"ac", X"b2", X"b5", X"ad", X"a4", X"b3", X"a1", X"78", X"74", X"5f", X"56", X"4e", X"3f", X"36", X"31", X"3b", X"2c", X"22", X"26", X"2c", X"2d", X"26", X"20", X"24", X"24", X"22", X"21", X"20", X"29", X"28", X"30", X"27", X"29", X"32", X"38", X"39", X"42", X"40", X"50", X"64", X"76", X"93", X"b2", X"af", X"aa", X"af", X"a1", X"a9", X"a5", X"9f", X"ab", X"9f", X"a1", X"9b", X"9c", X"98", X"91", X"94", X"8d", X"94", X"95", X"94", X"94", X"8d", X"8f", X"94", X"8c", X"8b", X"89", X"99", X"94", X"96", X"8d", X"8e", X"8c", X"8b", X"94", X"95", X"8e", X"96", X"8f", X"8f", X"8c", X"8c", X"97", X"8f", X"8d", X"8b", X"8d", X"8b", X"87", X"83", X"8b", X"80", X"7b", X"7e", X"75", X"7e", X"6c", X"72", X"69", X"62", X"63", X"5c", X"5b", X"5f", X"5e", X"5e", X"65", X"57", X"62", X"65", X"65", X"70", X"6e", X"6c", X"60", X"55", X"57", X"64", X"66", X"5b", X"48", X"43", X"31", X"29", X"24", X"1e", X"11", X"17", X"11", X"18", X"0c", X"0a", X"06", X"0b", X"03", X"09", X"06", X"05", X"08", X"0c", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"0b", X"0c", X"0b", X"04", X"0d", X"0f", X"0e", X"13", X"1d", X"1a", X"27", X"2f", X"3a", X"41", X"3d", X"3d", X"41", X"47", X"65", X"84", X"8a", X"86", X"81", X"82", X"87", X"98", X"98", X"98", X"9d", X"a5", X"a7", X"aa", X"ba", X"bc", X"bb", X"ba", X"be", X"c6", X"c0", X"c2", X"c1", X"c4", X"c5", X"b9", X"b4", X"b8", X"b1", X"ae", X"ae", X"ae", X"ad", X"ac", X"b1", X"b0", X"b0", X"a9", X"a9", X"ab", X"a5", X"a7", X"a0", X"a8", X"a9", X"ae", X"a9", X"a8", X"af", X"a6", X"b1", X"ab", X"af", X"b5", X"a9", X"ac", X"b1", X"bc", X"b5", X"b6", X"be", X"bb", X"b7", X"b5", X"b4", X"bb", X"b0", X"ae", X"b5", X"b5", X"b0", X"ab", X"aa", X"b1", X"aa", X"a8", X"a8", X"a4", X"ac", X"ab", X"a8", X"aa", X"a5", X"91", X"7d", X"65", X"5a", X"4a", X"44", X"37", X"39", X"21", X"28", X"25", X"24", X"28", X"25", X"1f", X"22", X"24", X"25", X"24", X"26", X"21", X"20", X"26", X"22", X"24", X"26", X"26", X"21", X"2f", X"3e", X"40", X"3c", X"49", X"59", X"6c", X"7e", X"a8", X"aa", X"a6", X"af", X"a4", X"9f", X"a0", X"a0", X"a2", X"9c", X"97", X"9d", X"99", X"91", X"92", X"92", X"8e", X"91", X"8f", X"93", X"8f", X"95", X"91", X"8e", X"8f", X"91", X"97", X"94", X"95", X"8f", X"97", X"8d", X"94", X"98", X"92", X"98", X"8f", X"8f", X"99", X"91", X"89", X"99", X"98", X"8f", X"8a", X"94", X"8b", X"88", X"7f", X"7c", X"79", X"79", X"78", X"70", X"6f", X"6e", X"6b", X"66", X"60", X"64", X"66", X"61", X"53", X"61", X"57", X"59", X"5c", X"65", X"66", X"64", X"6f", X"6b", X"6d", X"62", X"57", X"4e", X"5a", X"5e", X"54", X"59", X"50", X"3e", X"32", X"26", X"2a", X"21", X"1a", X"16", X"16", X"11", X"0d", X"0f", X"0b", X"0c", X"07", X"03", X"08", X"06", X"10", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"05", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"04", X"06", X"05", X"03", X"0f", X"06", X"0a", X"11", X"0f", X"0e", X"0e", X"1a", X"16", X"1f", X"1f", X"2a", X"38", X"41", X"3d", X"41", X"3d", X"49", X"61", X"77", X"85", X"89", X"7e", X"71", X"74", X"89", X"89", X"91", X"97", X"9a", X"a4", X"a8", X"a7", X"b3", X"b5", X"be", X"b6", X"bb", X"be", X"be", X"bb", X"b6", X"ba", X"b6", X"b7", X"b5", X"b8", X"ad", X"b2", X"ac", X"ae", X"b0", X"a9", X"a7", X"a9", X"aa", X"9f", X"a4", X"a6", X"a2", X"9b", X"a3", X"a9", X"a5", X"a5", X"ac", X"a0", X"a6", X"a2", X"a2", X"ae", X"aa", X"a4", X"a5", X"ab", X"aa", X"a9", X"ae", X"ae", X"a6", X"aa", X"ad", X"ac", X"ac", X"ae", X"a6", X"a7", X"a9", X"ad", X"a9", X"a8", X"a6", X"a1", X"a9", X"ad", X"a6", X"a5", X"a1", X"9c", X"97", X"9d", X"85", X"7c", X"60", X"45", X"3b", X"32", X"32", X"27", X"23", X"20", X"15", X"1f", X"15", X"18", X"19", X"1e", X"16", X"20", X"1d", X"14", X"17", X"21", X"1c", X"1e", X"24", X"17", X"26", X"29", X"2d", X"30", X"2c", X"2f", X"3e", X"5b", X"67", X"7d", X"a0", X"9d", X"a3", X"a1", X"a2", X"a1", X"96", X"a2", X"9e", X"9b", X"93", X"91", X"8d", X"94", X"94", X"95", X"91", X"8f", X"91", X"8b", X"8c", X"9a", X"90", X"92", X"93", X"8a", X"99", X"9b", X"9c", X"90", X"97", X"a0", X"91", X"9b", X"8a", X"90", X"91", X"92", X"90", X"97", X"90", X"94", X"94", X"8c", X"8d", X"89", X"89", X"86", X"7c", X"79", X"79", X"72", X"70", X"69", X"65", X"68", X"64", X"61", X"5a", X"58", X"58", X"53", X"50", X"52", X"59", X"5b", X"54", X"5e", X"60", X"60", X"6a", X"63", X"64", X"52", X"4c", X"46", X"56", X"64", X"56", X"5b", X"45", X"3e", X"36", X"31", X"20", X"20", X"16", X"15", X"10", X"0d", X"0d", X"0b", X"06", X"0b", X"04", X"05", X"07", X"05", X"03", X"00", X"0d", X"05", X"03", X"05", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"06", X"03", X"0c", X"06", X"08", X"0f", X"0a", X"0f", X"16", X"1a", X"21", X"28", X"29", X"34", X"36", X"3a", X"43", X"3e", X"3f", X"4b", X"59", X"76", X"87", X"87", X"7f", X"7c", X"76", X"7d", X"83", X"8c", X"8f", X"98", X"ab", X"9b", X"a4", X"aa", X"a5", X"af", X"ae", X"b3", X"b5", X"b8", X"b6", X"c0", X"c2", X"be", X"af", X"b6", X"ae", X"b2", X"ab", X"b0", X"b2", X"ae", X"ae", X"aa", X"a7", X"a8", X"a1", X"9e", X"96", X"a5", X"a3", X"97", X"a0", X"9d", X"9f", X"9c", X"a5", X"a5", X"a1", X"a2", X"a5", X"a3", X"9f", X"9d", X"aa", X"aa", X"a4", X"ab", X"ae", X"a3", X"a6", X"a6", X"a5", X"a5", X"a8", X"a1", X"a9", X"a4", X"a0", X"a8", X"a3", X"a5", X"9f", X"ab", X"aa", X"a3", X"9f", X"a0", X"96", X"9b", X"95", X"81", X"69", X"53", X"49", X"3a", X"32", X"2d", X"28", X"1e", X"1b", X"17", X"20", X"15", X"18", X"1a", X"11", X"16", X"17", X"17", X"1a", X"15", X"19", X"12", X"17", X"13", X"1b", X"1a", X"1f", X"23", X"1b", X"30", X"31", X"38", X"4c", X"63", X"7c", X"96", X"a3", X"a6", X"9e", X"9d", X"a2", X"93", X"98", X"9c", X"97", X"96", X"93", X"8f", X"89", X"94", X"92", X"8d", X"94", X"8b", X"96", X"8d", X"95", X"8d", X"92", X"91", X"98", X"9b", X"94", X"95", X"9c", X"9b", X"a0", X"9b", X"a2", X"9c", X"95", X"9a", X"96", X"8d", X"91", X"93", X"96", X"94", X"89", X"90", X"78", X"7d", X"7e", X"72", X"6f", X"6a", X"70", X"69", X"67", X"65", X"66", X"62", X"56", X"58", X"4e", X"55", X"55", X"59", X"59", X"5e", X"5a", X"52", X"69", X"53", X"64", X"5d", X"61", X"5f", X"54", X"59", X"4d", X"54", X"60", X"61", X"5a", X"4b", X"3a", X"33", X"20", X"22", X"1e", X"16", X"13", X"16", X"15", X"05", X"02", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"04", X"06", X"05", X"05", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"06", X"07", X"07", X"0d", X"11", X"0e", X"15", X"16", X"19", X"1f", X"27", X"24", X"34", X"39", X"3c", X"3f", X"3a", X"3f", X"4a", X"5b", X"6f", X"7b", X"81", X"7f", X"76", X"6c", X"75", X"77", X"7f", X"85", X"8a", X"9e", X"99", X"97", X"a0", X"a4", X"a4", X"a3", X"b2", X"b5", X"ae", X"b4", X"b5", X"bd", X"c4", X"b0", X"b1", X"ae", X"ae", X"a7", X"b3", X"b4", X"b9", X"b0", X"a9", X"a6", X"a0", X"98", X"9d", X"9f", X"9c", X"a0", X"a0", X"9d", X"a0", X"a1", X"9f", X"a1", X"a3", X"a0", X"a1", X"a5", X"a7", X"9e", X"a5", X"a1", X"a5", X"a2", X"a9", X"9b", X"a3", X"9d", X"9e", X"a2", X"a0", X"a3", X"a0", X"9f", X"9d", X"a4", X"a6", X"a2", X"a4", X"9f", X"9f", X"9f", X"9e", X"9e", X"96", X"96", X"9a", X"94", X"84", X"66", X"4c", X"2f", X"33", X"2c", X"21", X"27", X"23", X"20", X"19", X"11", X"12", X"14", X"18", X"18", X"10", X"11", X"17", X"18", X"14", X"1c", X"16", X"13", X"14", X"1b", X"1b", X"21", X"25", X"30", X"27", X"2b", X"2a", X"49", X"5e", X"80", X"a1", X"a7", X"a2", X"a0", X"96", X"9b", X"92", X"94", X"9c", X"91", X"8c", X"90", X"8a", X"9b", X"8c", X"8f", X"92", X"89", X"8b", X"8f", X"94", X"93", X"95", X"94", X"96", X"97", X"9a", X"9e", X"a0", X"a9", X"a3", X"9a", X"9a", X"9b", X"9a", X"92", X"90", X"93", X"86", X"8a", X"8b", X"86", X"90", X"80", X"79", X"7d", X"78", X"70", X"6b", X"70", X"67", X"63", X"64", X"60", X"59", X"60", X"5f", X"5a", X"57", X"4f", X"59", X"50", X"50", X"54", X"4d", X"52", X"59", X"57", X"5e", X"67", X"57", X"63", X"52", X"4f", X"54", X"5b", X"5e", X"63", X"57", X"59", X"4d", X"45", X"3b", X"27", X"25", X"22", X"1c", X"15", X"15", X"14", X"12", X"06", X"06", X"06", X"03", X"0d", X"06", X"05", X"07", X"00", X"0a", X"05", X"03", X"07", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"02", X"06", X"05", X"04", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"0d", X"09", X"06", X"07", X"07", X"0a", X"0e", X"13", X"17", X"1b", X"22", X"27", X"2c", X"34", X"36", X"37", X"39", X"3a", X"45", X"4a", X"5a", X"75", X"75", X"74", X"74", X"6d", X"72", X"73", X"70", X"75", X"82", X"85", X"90", X"8d", X"95", X"99", X"a2", X"a1", X"9e", X"a6", X"a9", X"aa", X"b3", X"b7", X"af", X"b5", X"ae", X"b3", X"ae", X"b2", X"af", X"ac", X"ae", X"ad", X"a7", X"ad", X"a5", X"9e", X"99", X"96", X"97", X"9d", X"9e", X"a2", X"99", X"9e", X"9e", X"8d", X"9b", X"a0", X"9e", X"97", X"a0", X"97", X"9b", X"98", X"9e", X"a9", X"9c", X"a2", X"9b", X"9d", X"91", X"9f", X"9f", X"a0", X"a1", X"a5", X"9b", X"9b", X"96", X"99", X"9f", X"9b", X"9b", X"95", X"96", X"96", X"98", X"96", X"90", X"91", X"8b", X"79", X"68", X"4d", X"3b", X"31", X"28", X"1e", X"1d", X"14", X"15", X"13", X"10", X"10", X"10", X"0b", X"17", X"15", X"05", X"13", X"09", X"0c", X"09", X"0f", X"13", X"09", X"0d", X"10", X"1a", X"16", X"2b", X"23", X"1e", X"23", X"3b", X"67", X"80", X"9d", X"9e", X"99", X"96", X"96", X"91", X"8d", X"96", X"8d", X"8f", X"89", X"98", X"8f", X"8e", X"99", X"91", X"8c", X"8d", X"8f", X"85", X"89", X"8c", X"8f", X"91", X"8d", X"9d", X"a2", X"a1", X"a0", X"a0", X"a0", X"a0", X"9b", X"9d", X"9b", X"99", X"90", X"8f", X"8a", X"89", X"87", X"82", X"7a", X"7c", X"7f", X"72", X"67", X"6d", X"65", X"68", X"66", X"61", X"58", X"62", X"4f", X"5a", X"51", X"55", X"5e", X"50", X"4c", X"4b", X"4a", X"51", X"4f", X"4c", X"55", X"57", X"59", X"5a", X"5a", X"51", X"50", X"4d", X"4f", X"4e", X"5b", X"5c", X"60", X"54", X"4b", X"40", X"3c", X"2d", X"23", X"26", X"1b", X"15", X"10", X"07", X"08", X"07", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"01", X"0d", X"0a", X"09", X"11", X"11", X"16", X"1c", X"1f", X"22", X"25", X"34", X"36", X"33", X"37", X"39", X"39", X"47", X"5c", X"70", X"76", X"78", X"6f", X"65", X"6d", X"6d", X"71", X"6e", X"6e", X"71", X"7b", X"8c", X"83", X"91", X"99", X"9b", X"99", X"a4", X"a7", X"a8", X"ae", X"b4", X"a9", X"ae", X"a8", X"b3", X"b3", X"ab", X"b3", X"b2", X"b0", X"b1", X"ad", X"a7", X"a3", X"a0", X"98", X"99", X"9c", X"a0", X"8f", X"98", X"9b", X"9b", X"90", X"95", X"9e", X"94", X"98", X"96", X"a0", X"9d", X"9c", X"96", X"9e", X"9a", X"90", X"93", X"91", X"a0", X"95", X"96", X"94", X"9f", X"9a", X"9c", X"95", X"8e", X"92", X"91", X"94", X"92", X"96", X"94", X"99", X"91", X"9b", X"94", X"8e", X"85", X"85", X"81", X"62", X"4a", X"3b", X"2d", X"1f", X"15", X"12", X"19", X"10", X"0f", X"09", X"0e", X"0b", X"0c", X"0d", X"0c", X"0a", X"09", X"09", X"0b", X"09", X"08", X"0d", X"0e", X"10", X"15", X"0f", X"15", X"19", X"20", X"1b", X"20", X"34", X"65", X"95", X"9f", X"a1", X"9e", X"97", X"95", X"99", X"8d", X"90", X"8f", X"95", X"92", X"98", X"91", X"8d", X"8b", X"84", X"92", X"8a", X"8a", X"8d", X"8a", X"8f", X"97", X"89", X"94", X"95", X"9b", X"9f", X"9f", X"a3", X"9d", X"97", X"97", X"92", X"92", X"98", X"8a", X"8a", X"80", X"80", X"78", X"7b", X"79", X"70", X"70", X"70", X"66", X"63", X"64", X"60", X"54", X"56", X"5d", X"52", X"58", X"4f", X"50", X"51", X"53", X"49", X"52", X"50", X"4a", X"4c", X"4c", X"4c", X"4f", X"50", X"53", X"4b", X"51", X"50", X"47", X"46", X"47", X"4f", X"52", X"64", X"5d", X"52", X"43", X"40", X"36", X"27", X"25", X"1b", X"0a", X"0e", X"0c", X"12", X"06", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"08", X"05", X"06", X"05", X"07", X"0e", X"06", X"0d", X"0e", X"1a", X"1e", X"22", X"20", X"2a", X"25", X"3a", X"39", X"3a", X"3e", X"41", X"46", X"56", X"6f", X"78", X"73", X"71", X"73", X"6c", X"6d", X"6f", X"73", X"6e", X"6b", X"70", X"7b", X"80", X"8d", X"96", X"97", X"9a", X"9d", X"a5", X"ac", X"ac", X"a5", X"b0", X"ae", X"b1", X"b4", X"b7", X"b1", X"b1", X"b2", X"b5", X"b9", X"b2", X"a0", X"a1", X"9f", X"a2", X"9c", X"9a", X"a0", X"9a", X"97", X"97", X"97", X"8f", X"99", X"9d", X"98", X"9c", X"9c", X"a2", X"9a", X"91", X"9c", X"98", X"a3", X"99", X"95", X"8c", X"9a", X"a0", X"95", X"96", X"9a", X"91", X"99", X"95", X"92", X"8e", X"8b", X"99", X"89", X"93", X"90", X"8b", X"8a", X"92", X"8e", X"8a", X"8f", X"8b", X"82", X"6d", X"51", X"40", X"2c", X"1e", X"1b", X"0b", X"0b", X"08", X"09", X"09", X"10", X"13", X"0d", X"09", X"11", X"0b", X"0d", X"0e", X"0d", X"05", X"0a", X"0d", X"0d", X"12", X"09", X"06", X"10", X"1c", X"20", X"20", X"29", X"2a", X"62", X"8d", X"9c", X"a2", X"9b", X"99", X"97", X"97", X"8f", X"93", X"8e", X"94", X"8b", X"8c", X"95", X"8e", X"81", X"86", X"87", X"8b", X"88", X"88", X"85", X"94", X"81", X"89", X"96", X"9f", X"9e", X"96", X"9b", X"91", X"90", X"93", X"90", X"94", X"8c", X"8c", X"7f", X"7d", X"7a", X"6b", X"71", X"6d", X"69", X"6f", X"70", X"67", X"6d", X"5c", X"58", X"5b", X"5e", X"58", X"58", X"59", X"51", X"52", X"4d", X"4c", X"53", X"4e", X"4f", X"45", X"50", X"4e", X"57", X"59", X"4f", X"55", X"4e", X"52", X"49", X"4d", X"49", X"4b", X"4a", X"4f", X"47", X"60", X"55", X"51", X"4f", X"3e", X"33", X"2e", X"23", X"1c", X"16", X"0d", X"08", X"09", X"03", X"00", X"06", X"06", X"03", X"05", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"10", X"06", X"0b", X"09", X"0f", X"12", X"14", X"17", X"22", X"21", X"2d", X"33", X"33", X"38", X"3a", X"37", X"3f", X"41", X"55", X"6c", X"71", X"76", X"6b", X"6f", X"70", X"68", X"72", X"73", X"67", X"6f", X"77", X"74", X"7a", X"7e", X"86", X"8d", X"92", X"9a", X"9d", X"a4", X"a2", X"a6", X"ab", X"b3", X"b5", X"b5", X"b4", X"b4", X"b1", X"b1", X"b2", X"b1", X"b1", X"ab", X"ab", X"a7", X"a5", X"a4", X"9e", X"98", X"9f", X"98", X"93", X"99", X"95", X"96", X"98", X"9b", X"a0", X"9c", X"9c", X"91", X"98", X"99", X"91", X"a0", X"97", X"97", X"99", X"93", X"92", X"94", X"88", X"95", X"89", X"92", X"9b", X"8e", X"90", X"92", X"8d", X"92", X"98", X"8d", X"8f", X"8f", X"8a", X"86", X"84", X"82", X"83", X"89", X"71", X"5b", X"45", X"25", X"18", X"0d", X"10", X"13", X"0b", X"0f", X"07", X"06", X"12", X"04", X"05", X"06", X"06", X"07", X"14", X"10", X"0c", X"07", X"06", X"06", X"0a", X"17", X"15", X"12", X"1b", X"16", X"19", X"1c", X"2b", X"5d", X"8d", X"9e", X"96", X"98", X"94", X"8d", X"8c", X"90", X"8b", X"8f", X"8a", X"8c", X"8f", X"84", X"8b", X"8b", X"87", X"8f", X"87", X"88", X"85", X"86", X"8b", X"89", X"8c", X"8c", X"99", X"8d", X"94", X"8f", X"8e", X"8f", X"8e", X"88", X"87", X"85", X"81", X"76", X"6c", X"70", X"62", X"6d", X"72", X"6c", X"64", X"69", X"64", X"65", X"59", X"62", X"51", X"56", X"51", X"55", X"4a", X"53", X"53", X"48", X"52", X"4b", X"4a", X"50", X"4c", X"49", X"4f", X"4c", X"50", X"52", X"5c", X"52", X"4c", X"47", X"4a", X"47", X"47", X"46", X"51", X"55", X"64", X"58", X"59", X"4b", X"42", X"3a", X"28", X"24", X"21", X"1a", X"18", X"0c", X"06", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"14", X"15", X"1d", X"18", X"1e", X"24", X"31", X"31", X"37", X"40", X"33", X"36", X"40", X"49", X"61", X"64", X"65", X"6c", X"67", X"69", X"76", X"72", X"70", X"68", X"60", X"68", X"68", X"70", X"74", X"78", X"76", X"79", X"85", X"8e", X"94", X"99", X"9f", X"a2", X"9b", X"a7", X"a8", X"b2", X"a8", X"b0", X"b8", X"b2", X"b6", X"b2", X"ac", X"b0", X"ab", X"a9", X"a8", X"a7", X"a6", X"9e", X"a5", X"a0", X"a0", X"a0", X"a1", X"9d", X"a8", X"98", X"96", X"94", X"95", X"94", X"99", X"9e", X"9b", X"a0", X"98", X"96", X"93", X"9d", X"8b", X"92", X"93", X"92", X"88", X"95", X"8c", X"92", X"86", X"95", X"8d", X"8b", X"8b", X"91", X"87", X"98", X"86", X"87", X"89", X"7e", X"7f", X"75", X"59", X"39", X"20", X"12", X"09", X"0a", X"0b", X"05", X"03", X"07", X"06", X"06", X"03", X"00", X"08", X"09", X"05", X"05", X"06", X"09", X"05", X"0b", X"06", X"05", X"0d", X"05", X"0b", X"06", X"11", X"16", X"18", X"2c", X"56", X"81", X"95", X"90", X"8e", X"8a", X"89", X"8d", X"8e", X"83", X"85", X"84", X"81", X"86", X"87", X"8a", X"82", X"86", X"80", X"82", X"85", X"84", X"85", X"89", X"83", X"85", X"8c", X"8e", X"8f", X"8c", X"81", X"84", X"7f", X"7f", X"81", X"71", X"73", X"6f", X"75", X"6f", X"64", X"5f", X"64", X"64", X"64", X"64", X"60", X"66", X"55", X"55", X"4d", X"59", X"57", X"4f", X"4b", X"43", X"48", X"4d", X"4b", X"4e", X"49", X"49", X"52", X"44", X"48", X"42", X"52", X"53", X"52", X"59", X"4e", X"52", X"47", X"3a", X"43", X"3a", X"40", X"4b", X"59", X"64", X"62", X"58", X"4d", X"44", X"32", X"21", X"26", X"15", X"18", X"0b", X"0f", X"05", X"07", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"0d", X"06", X"10", X"16", X"1a", X"17", X"1f", X"26", X"2f", X"30", X"3f", X"33", X"35", X"31", X"3f", X"41", X"51", X"58", X"64", X"63", X"67", X"68", X"69", X"6e", X"6a", X"73", X"6e", X"67", X"6f", X"68", X"6f", X"6f", X"6c", X"7a", X"7a", X"75", X"80", X"86", X"8c", X"94", X"9b", X"9d", X"aa", X"a4", X"ad", X"ad", X"b0", X"b6", X"b5", X"bd", X"b9", X"af", X"b8", X"b1", X"ad", X"b0", X"af", X"af", X"a9", X"a4", X"ab", X"ab", X"ab", X"a9", X"a6", X"a6", X"9a", X"9e", X"a0", X"a3", X"9a", X"a0", X"9d", X"9d", X"a6", X"94", X"97", X"96", X"8f", X"9d", X"97", X"91", X"9a", X"93", X"98", X"91", X"91", X"8b", X"8e", X"8d", X"8f", X"94", X"85", X"86", X"88", X"83", X"82", X"85", X"7f", X"76", X"76", X"62", X"37", X"19", X"1b", X"0a", X"09", X"09", X"05", X"0b", X"0a", X"0b", X"05", X"04", X"00", X"07", X"08", X"03", X"04", X"08", X"05", X"06", X"07", X"0b", X"0a", X"06", X"0c", X"0f", X"0b", X"11", X"17", X"11", X"27", X"4a", X"7d", X"8f", X"82", X"8e", X"8d", X"82", X"87", X"81", X"84", X"85", X"84", X"81", X"79", X"7f", X"7a", X"7d", X"7a", X"85", X"86", X"83", X"89", X"81", X"7a", X"8c", X"7e", X"86", X"89", X"87", X"86", X"75", X"79", X"78", X"6f", X"6e", X"70", X"73", X"70", X"6a", X"6d", X"65", X"65", X"64", X"65", X"6e", X"64", X"5f", X"62", X"52", X"56", X"57", X"59", X"4f", X"54", X"53", X"4d", X"4b", X"4b", X"4b", X"46", X"44", X"41", X"48", X"4b", X"4a", X"4e", X"52", X"54", X"4e", X"50", X"4c", X"48", X"4a", X"43", X"46", X"3c", X"3e", X"41", X"54", X"62", X"5f", X"57", X"48", X"41", X"35", X"2a", X"20", X"22", X"1b", X"0f", X"11", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"08", X"06", X"05", X"0e", X"09", X"0b", X"14", X"15", X"28", X"24", X"2c", X"32", X"35", X"42", X"33", X"31", X"3f", X"49", X"4e", X"62", X"5f", X"5d", X"66", X"61", X"66", X"6c", X"6e", X"70", X"69", X"71", X"75", X"68", X"6f", X"73", X"69", X"73", X"71", X"73", X"75", X"7b", X"7a", X"83", X"87", X"8b", X"9f", X"97", X"a1", X"aa", X"b4", X"b4", X"b8", X"b2", X"b9", X"ae", X"b5", X"af", X"b6", X"b7", X"b5", X"b5", X"a9", X"ac", X"b0", X"a9", X"a6", X"ae", X"b1", X"a3", X"a8", X"a5", X"a6", X"a5", X"a4", X"a0", X"a3", X"ab", X"9a", X"a5", X"9e", X"9c", X"9f", X"96", X"97", X"9c", X"9f", X"92", X"95", X"98", X"92", X"8e", X"95", X"8f", X"8d", X"8f", X"85", X"8b", X"8e", X"8a", X"8f", X"84", X"82", X"85", X"75", X"59", X"32", X"1a", X"0e", X"0f", X"0c", X"06", X"05", X"03", X"0b", X"0e", X"05", X"03", X"00", X"06", X"05", X"0a", X"00", X"06", X"05", X"03", X"00", X"06", X"0b", X"06", X"0c", X"0e", X"10", X"14", X"0d", X"12", X"22", X"49", X"7d", X"8d", X"8a", X"83", X"7c", X"7b", X"7d", X"7f", X"81", X"80", X"7e", X"75", X"81", X"77", X"7d", X"81", X"7e", X"7a", X"84", X"7c", X"85", X"82", X"7d", X"78", X"7a", X"79", X"7e", X"7b", X"76", X"70", X"6d", X"74", X"6e", X"6b", X"65", X"69", X"69", X"6a", X"68", X"61", X"64", X"63", X"64", X"63", X"5b", X"60", X"60", X"4e", X"55", X"54", X"54", X"53", X"52", X"4b", X"50", X"4e", X"4b", X"4c", X"4a", X"4c", X"4d", X"48", X"4a", X"47", X"49", X"57", X"4c", X"4a", X"4a", X"4c", X"55", X"44", X"3b", X"3c", X"40", X"43", X"47", X"4f", X"60", X"5b", X"4e", X"44", X"45", X"37", X"27", X"23", X"19", X"11", X"10", X"06", X"05", X"05", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0a", X"00", X"0a", X"14", X"12", X"20", X"23", X"2a", X"39", X"38", X"3d", X"35", X"36", X"3b", X"40", X"52", X"5d", X"5e", X"5d", X"5b", X"5b", X"60", X"5e", X"66", X"62", X"67", X"69", X"68", X"72", X"68", X"70", X"64", X"6c", X"6f", X"75", X"6b", X"69", X"6e", X"78", X"77", X"81", X"8c", X"88", X"94", X"a0", X"a0", X"a8", X"aa", X"a5", X"ab", X"a7", X"a6", X"a1", X"ae", X"b0", X"b5", X"af", X"ad", X"ae", X"ac", X"a8", X"a8", X"b1", X"ae", X"b2", X"ac", X"a6", X"ad", X"a7", X"a6", X"a7", X"a5", X"a3", X"a8", X"a0", X"a0", X"9d", X"a0", X"9c", X"a0", X"9e", X"99", X"95", X"9b", X"95", X"94", X"99", X"96", X"97", X"85", X"95", X"90", X"8d", X"8e", X"85", X"84", X"81", X"86", X"7b", X"7d", X"5d", X"2d", X"15", X"05", X"0d", X"03", X"06", X"05", X"05", X"01", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"08", X"0f", X"06", X"0e", X"11", X"0e", X"14", X"18", X"38", X"70", X"81", X"84", X"7f", X"7f", X"71", X"7c", X"70", X"7c", X"80", X"7d", X"74", X"78", X"72", X"74", X"75", X"79", X"70", X"6f", X"7a", X"72", X"76", X"78", X"6d", X"6d", X"72", X"69", X"6b", X"6f", X"68", X"6d", X"70", X"6a", X"66", X"65", X"62", X"5f", X"64", X"62", X"62", X"5f", X"60", X"5f", X"55", X"5f", X"55", X"58", X"58", X"56", X"4b", X"4f", X"4a", X"4e", X"4d", X"4e", X"42", X"43", X"3b", X"51", X"45", X"4b", X"51", X"44", X"49", X"4b", X"4b", X"52", X"4d", X"4d", X"4a", X"48", X"39", X"37", X"3b", X"35", X"41", X"41", X"4e", X"66", X"52", X"50", X"4c", X"3b", X"32", X"2b", X"1e", X"1a", X"1a", X"0b", X"16", X"05", X"06", X"01", X"06", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"04", X"06", X"0a", X"17", X"19", X"25", X"26", X"39", X"36", X"3a", X"3a", X"3b", X"3d", X"43", X"47", X"58", X"59", X"56", X"5d", X"52", X"5c", X"5d", X"62", X"6c", X"6a", X"6f", X"6e", X"6a", X"70", X"72", X"6e", X"6e", X"6a", X"6a", X"6d", X"69", X"72", X"70", X"72", X"6f", X"70", X"7a", X"7b", X"84", X"8c", X"91", X"90", X"97", X"98", X"a3", X"a5", X"9d", X"a0", X"aa", X"a3", X"b4", X"a7", X"ac", X"ac", X"ad", X"ac", X"aa", X"b2", X"aa", X"a9", X"af", X"a5", X"aa", X"a7", X"a2", X"aa", X"a8", X"a5", X"aa", X"a5", X"a1", X"9c", X"9c", X"9e", X"9b", X"92", X"98", X"99", X"99", X"96", X"92", X"8c", X"8e", X"97", X"8d", X"8f", X"85", X"8b", X"8e", X"8a", X"7b", X"82", X"7e", X"77", X"60", X"32", X"18", X"0d", X"04", X"01", X"06", X"05", X"05", X"05", X"06", X"07", X"06", X"03", X"07", X"05", X"08", X"00", X"06", X"05", X"04", X"04", X"06", X"09", X"07", X"0c", X"0d", X"0a", X"06", X"08", X"0e", X"1c", X"3c", X"6e", X"78", X"7d", X"79", X"78", X"6d", X"78", X"75", X"73", X"74", X"6e", X"79", X"75", X"71", X"6e", X"6d", X"73", X"70", X"79", X"71", X"6d", X"61", X"71", X"73", X"66", X"6b", X"6a", X"67", X"63", X"5c", X"64", X"5c", X"69", X"65", X"64", X"62", X"5f", X"60", X"60", X"61", X"52", X"56", X"5c", X"56", X"51", X"5b", X"53", X"4a", X"52", X"5a", X"4b", X"54", X"56", X"4c", X"46", X"42", X"4b", X"53", X"45", X"48", X"42", X"45", X"48", X"4c", X"4e", X"52", X"4c", X"3e", X"43", X"47", X"47", X"45", X"3a", X"46", X"35", X"41", X"41", X"55", X"5a", X"51", X"50", X"49", X"47", X"36", X"2f", X"18", X"14", X"12", X"12", X"0e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"09", X"08", X"0d", X"12", X"19", X"29", X"28", X"2f", X"3f", X"3b", X"3b", X"3a", X"3d", X"46", X"50", X"5f", X"57", X"5a", X"58", X"51", X"56", X"59", X"5d", X"5c", X"63", X"6e", X"6b", X"73", X"61", X"6b", X"73", X"74", X"78", X"78", X"72", X"73", X"63", X"6d", X"67", X"6c", X"6e", X"73", X"73", X"71", X"7e", X"75", X"82", X"81", X"88", X"96", X"8d", X"92", X"9e", X"a2", X"98", X"9f", X"9f", X"9c", X"a0", X"a4", X"ae", X"a4", X"ae", X"aa", X"a6", X"a4", X"a9", X"a1", X"a1", X"a6", X"a4", X"a8", X"a1", X"a6", X"9d", X"9c", X"99", X"9a", X"97", X"9b", X"8c", X"97", X"94", X"94", X"9b", X"94", X"9c", X"95", X"90", X"91", X"8d", X"7d", X"80", X"86", X"84", X"7e", X"81", X"80", X"6c", X"5d", X"2f", X"18", X"08", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"06", X"06", X"00", X"06", X"06", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"08", X"0f", X"00", X"10", X"0e", X"09", X"0c", X"07", X"16", X"32", X"5f", X"75", X"82", X"77", X"75", X"6c", X"75", X"74", X"70", X"74", X"75", X"75", X"76", X"6b", X"69", X"75", X"78", X"73", X"71", X"6b", X"6d", X"6a", X"6d", X"6e", X"6b", X"66", X"65", X"69", X"5f", X"68", X"61", X"61", X"60", X"64", X"62", X"60", X"62", X"60", X"59", X"57", X"58", X"55", X"5b", X"59", X"61", X"5d", X"5e", X"54", X"4f", X"5b", X"4e", X"54", X"4f", X"43", X"47", X"47", X"55", X"52", X"55", X"51", X"4b", X"4c", X"4d", X"4c", X"49", X"4b", X"4a", X"38", X"4d", X"3f", X"41", X"41", X"41", X"37", X"3e", X"3c", X"4b", X"51", X"5d", X"50", X"4f", X"3f", X"35", X"2a", X"26", X"1e", X"19", X"12", X"08", X"0e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"06", X"09", X"0f", X"1b", X"28", X"2e", X"33", X"39", X"35", X"2c", X"33", X"3e", X"4c", X"62", X"5a", X"52", X"50", X"4f", X"53", X"52", X"54", X"57", X"55", X"64", X"62", X"5c", X"69", X"64", X"6e", X"74", X"7b", X"84", X"77", X"6e", X"6f", X"68", X"68", X"72", X"66", X"6e", X"6d", X"6a", X"68", X"67", X"77", X"71", X"79", X"79", X"7e", X"7a", X"88", X"8f", X"8b", X"8e", X"88", X"92", X"90", X"9c", X"96", X"93", X"99", X"9c", X"98", X"9a", X"96", X"9a", X"8b", X"88", X"97", X"94", X"94", X"9a", X"98", X"92", X"8c", X"92", X"90", X"88", X"89", X"89", X"8d", X"85", X"90", X"85", X"7d", X"84", X"82", X"83", X"7c", X"83", X"83", X"81", X"7b", X"82", X"82", X"76", X"6c", X"54", X"28", X"0b", X"05", X"0a", X"07", X"06", X"05", X"03", X"04", X"06", X"05", X"04", X"01", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0a", X"06", X"0c", X"0b", X"09", X"0b", X"13", X"2a", X"61", X"80", X"7d", X"76", X"73", X"6d", X"72", X"6f", X"6d", X"6e", X"6e", X"66", X"71", X"6d", X"6b", X"6d", X"66", X"6f", X"70", X"70", X"6b", X"66", X"6a", X"67", X"64", X"66", X"66", X"65", X"62", X"65", X"56", X"5b", X"61", X"64", X"5f", X"53", X"5b", X"59", X"4e", X"4d", X"58", X"4e", X"54", X"54", X"53", X"50", X"58", X"4e", X"51", X"56", X"4f", X"4e", X"4e", X"4e", X"4a", X"4c", X"48", X"57", X"49", X"4d", X"4e", X"47", X"47", X"48", X"4e", X"45", X"39", X"41", X"3d", X"45", X"44", X"38", X"41", X"32", X"41", X"40", X"44", X"5b", X"54", X"48", X"44", X"3e", X"37", X"2d", X"24", X"23", X"1c", X"13", X"08", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"08", X"06", X"07", X"0c", X"11", X"1e", X"23", X"2e", X"37", X"37", X"47", X"36", X"37", X"3d", X"44", X"52", X"50", X"57", X"54", X"50", X"56", X"5b", X"5b", X"5b", X"56", X"5d", X"5b", X"5d", X"61", X"65", X"64", X"6f", X"70", X"74", X"6d", X"79", X"78", X"6f", X"69", X"6b", X"6a", X"69", X"68", X"62", X"68", X"64", X"6b", X"68", X"6d", X"71", X"73", X"73", X"7a", X"86", X"86", X"81", X"7b", X"7f", X"85", X"7b", X"81", X"88", X"91", X"8f", X"8d", X"8e", X"91", X"8c", X"8a", X"83", X"90", X"8a", X"8c", X"86", X"8d", X"84", X"87", X"89", X"84", X"87", X"7c", X"80", X"84", X"84", X"80", X"7a", X"82", X"7b", X"7e", X"7e", X"81", X"7b", X"78", X"78", X"70", X"75", X"72", X"6b", X"6c", X"54", X"2b", X"18", X"0e", X"0a", X"08", X"06", X"05", X"03", X"01", X"06", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"0e", X"06", X"07", X"13", X"0d", X"0c", X"10", X"2e", X"60", X"74", X"79", X"72", X"70", X"68", X"72", X"67", X"74", X"6f", X"6b", X"6a", X"69", X"6a", X"72", X"67", X"6b", X"66", X"6b", X"68", X"6a", X"66", X"69", X"68", X"64", X"67", X"64", X"5d", X"61", X"59", X"55", X"5a", X"59", X"5a", X"5f", X"55", X"56", X"5d", X"56", X"54", X"55", X"59", X"5a", X"5d", X"4f", X"52", X"5d", X"50", X"4a", X"54", X"4f", X"53", X"4e", X"48", X"4d", X"40", X"4e", X"48", X"4e", X"4c", X"4b", X"52", X"4c", X"48", X"44", X"41", X"3e", X"3e", X"3b", X"3a", X"3f", X"3e", X"3e", X"3f", X"3e", X"46", X"4a", X"56", X"50", X"47", X"3d", X"36", X"31", X"2d", X"2b", X"1b", X"1a", X"0b", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"03", X"06", X"06", X"05", X"00", X"0a", X"05", X"08", X"11", X"1b", X"21", X"2e", X"37", X"39", X"41", X"43", X"3e", X"42", X"49", X"51", X"4d", X"56", X"51", X"51", X"4b", X"58", X"58", X"58", X"58", X"58", X"5c", X"5a", X"57", X"5e", X"61", X"60", X"69", X"67", X"67", X"70", X"6a", X"70", X"79", X"6d", X"73", X"6d", X"67", X"6a", X"6e", X"71", X"6c", X"6a", X"67", X"71", X"70", X"72", X"70", X"75", X"7b", X"77", X"72", X"79", X"75", X"6e", X"7d", X"78", X"82", X"83", X"7a", X"83", X"84", X"80", X"82", X"7f", X"82", X"82", X"83", X"82", X"85", X"88", X"82", X"79", X"7b", X"7d", X"7e", X"7f", X"7b", X"7b", X"78", X"76", X"70", X"78", X"77", X"77", X"7a", X"73", X"7c", X"74", X"76", X"76", X"6f", X"6d", X"67", X"5a", X"2d", X"0e", X"0b", X"09", X"07", X"06", X"05", X"03", X"03", X"09", X"05", X"03", X"01", X"06", X"05", X"05", X"00", X"06", X"05", X"04", X"05", X"06", X"05", X"03", X"04", X"06", X"06", X"0a", X"0e", X"12", X"10", X"2e", X"5f", X"67", X"71", X"67", X"68", X"62", X"73", X"65", X"71", X"71", X"64", X"70", X"6a", X"6c", X"65", X"6b", X"69", X"65", X"6b", X"64", X"60", X"63", X"68", X"60", X"61", X"5e", X"5d", X"55", X"5c", X"5d", X"58", X"51", X"5a", X"59", X"64", X"59", X"59", X"54", X"54", X"53", X"52", X"5a", X"55", X"5e", X"4f", X"4e", X"4f", X"48", X"56", X"4a", X"48", X"4a", X"4e", X"4e", X"49", X"45", X"4f", X"47", X"4a", X"4c", X"50", X"4b", X"53", X"40", X"45", X"44", X"47", X"40", X"45", X"3b", X"43", X"39", X"3f", X"44", X"40", X"39", X"42", X"54", X"58", X"43", X"39", X"34", X"33", X"34", X"28", X"1e", X"17", X"19", X"0a", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"09", X"07", X"06", X"04", X"0f", X"15", X"1d", X"2b", X"31", X"35", X"44", X"44", X"3e", X"40", X"4a", X"51", X"49", X"4f", X"50", X"51", X"57", X"59", X"5b", X"4e", X"4d", X"5a", X"51", X"56", X"5c", X"57", X"54", X"5e", X"57", X"68", X"5a", X"62", X"63", X"6c", X"67", X"65", X"6d", X"67", X"6c", X"71", X"6f", X"68", X"6b", X"64", X"62", X"72", X"6e", X"71", X"6d", X"77", X"70", X"70", X"70", X"76", X"6c", X"73", X"71", X"78", X"84", X"81", X"82", X"76", X"84", X"80", X"7c", X"76", X"7c", X"7d", X"82", X"7d", X"84", X"79", X"82", X"7e", X"82", X"7b", X"79", X"7e", X"7b", X"74", X"6f", X"77", X"76", X"73", X"73", X"73", X"75", X"71", X"78", X"6e", X"6a", X"73", X"6d", X"66", X"67", X"50", X"31", X"08", X"09", X"03", X"05", X"06", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"0a", X"07", X"0a", X"08", X"06", X"10", X"26", X"4d", X"6e", X"64", X"65", X"6a", X"61", X"6f", X"6b", X"62", X"69", X"6e", X"6c", X"70", X"65", X"6a", X"61", X"66", X"6d", X"64", X"61", X"61", X"5e", X"64", X"5d", X"64", X"5b", X"5c", X"5a", X"58", X"56", X"58", X"58", X"56", X"50", X"52", X"5a", X"53", X"58", X"57", X"50", X"53", X"59", X"51", X"50", X"51", X"52", X"56", X"4c", X"50", X"52", X"4f", X"4b", X"4e", X"4d", X"48", X"4c", X"46", X"43", X"4c", X"4e", X"55", X"50", X"47", X"44", X"3d", X"3f", X"38", X"3e", X"41", X"3d", X"45", X"3c", X"3b", X"36", X"3e", X"34", X"40", X"4e", X"40", X"34", X"34", X"2d", X"30", X"2a", X"23", X"1b", X"1a", X"0e", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"03", X"0a", X"15", X"1c", X"2a", X"38", X"35", X"44", X"3c", X"3d", X"3b", X"41", X"4b", X"4f", X"4d", X"4c", X"4c", X"4f", X"55", X"51", X"55", X"58", X"4c", X"55", X"55", X"57", X"59", X"58", X"54", X"58", X"5a", X"56", X"5d", X"66", X"62", X"64", X"63", X"69", X"68", X"67", X"70", X"6f", X"6e", X"6f", X"61", X"6b", X"65", X"6f", X"64", X"73", X"79", X"76", X"78", X"72", X"66", X"6d", X"6c", X"70", X"6f", X"6e", X"7a", X"7d", X"76", X"74", X"70", X"71", X"7a", X"72", X"80", X"82", X"7e", X"7b", X"7e", X"7c", X"7a", X"7b", X"7f", X"7c", X"77", X"6e", X"73", X"75", X"73", X"73", X"71", X"6e", X"6f", X"70", X"6e", X"6b", X"74", X"70", X"67", X"66", X"66", X"65", X"56", X"33", X"0f", X"0c", X"05", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"0a", X"03", X"02", X"06", X"05", X"1f", X"4e", X"69", X"6f", X"65", X"63", X"60", X"64", X"64", X"64", X"65", X"67", X"64", X"67", X"6e", X"6c", X"55", X"60", X"64", X"60", X"62", X"5d", X"5b", X"58", X"5c", X"52", X"56", X"59", X"58", X"55", X"55", X"56", X"5a", X"56", X"56", X"55", X"55", X"5e", X"59", X"57", X"54", X"59", X"5b", X"57", X"56", X"54", X"4e", X"49", X"48", X"51", X"49", X"49", X"49", X"44", X"4c", X"4f", X"49", X"48", X"4a", X"4d", X"49", X"4a", X"44", X"48", X"3c", X"3f", X"48", X"44", X"3c", X"36", X"36", X"41", X"41", X"46", X"3c", X"39", X"35", X"3d", X"3b", X"37", X"31", X"24", X"2d", X"2d", X"2e", X"1f", X"1e", X"13", X"0b", X"09", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"03", X"00", X"07", X"05", X"08", X"0f", X"0d", X"24", X"21", X"2f", X"3a", X"42", X"49", X"46", X"46", X"46", X"51", X"5b", X"57", X"54", X"49", X"4d", X"49", X"53", X"56", X"5c", X"5a", X"5d", X"5b", X"5b", X"56", X"56", X"5d", X"5c", X"57", X"60", X"51", X"59", X"62", X"5d", X"5e", X"5d", X"5f", X"65", X"67", X"6b", X"6a", X"6f", X"6f", X"66", X"6b", X"6a", X"6a", X"6f", X"7d", X"72", X"71", X"69", X"68", X"69", X"73", X"6c", X"70", X"73", X"77", X"74", X"78", X"7e", X"7a", X"6f", X"74", X"70", X"7b", X"75", X"7b", X"77", X"79", X"7d", X"74", X"76", X"7d", X"71", X"78", X"73", X"77", X"6b", X"76", X"7a", X"68", X"67", X"6a", X"6d", X"70", X"76", X"67", X"67", X"62", X"69", X"66", X"5b", X"56", X"32", X"12", X"09", X"03", X"02", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"08", X"0a", X"0a", X"09", X"08", X"1f", X"4d", X"60", X"68", X"63", X"6a", X"61", X"65", X"61", X"6c", X"6a", X"69", X"6c", X"5c", X"63", X"63", X"6c", X"5d", X"66", X"5d", X"62", X"5f", X"56", X"5b", X"5d", X"59", X"55", X"61", X"53", X"5c", X"60", X"59", X"53", X"52", X"56", X"4e", X"55", X"52", X"56", X"54", X"5d", X"5d", X"5b", X"55", X"52", X"56", X"57", X"56", X"52", X"47", X"4b", X"46", X"4e", X"4d", X"43", X"4f", X"48", X"4a", X"3f", X"47", X"4e", X"50", X"4c", X"45", X"3e", X"49", X"41", X"3b", X"3e", X"43", X"45", X"4a", X"3b", X"3e", X"41", X"3b", X"47", X"35", X"3b", X"33", X"2a", X"2f", X"2d", X"25", X"2e", X"20", X"17", X"16", X"14", X"0d", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"0a", X"07", X"09", X"1b", X"26", X"27", X"35", X"41", X"3c", X"46", X"49", X"58", X"61", X"68", X"61", X"5c", X"53", X"59", X"4d", X"55", X"50", X"4b", X"55", X"56", X"55", X"58", X"54", X"57", X"5e", X"5c", X"5c", X"59", X"53", X"56", X"55", X"5d", X"58", X"5d", X"63", X"5d", X"5b", X"69", X"63", X"69", X"72", X"6b", X"6e", X"64", X"6c", X"6a", X"72", X"67", X"6f", X"69", X"66", X"6e", X"64", X"6b", X"72", X"75", X"76", X"74", X"6d", X"6b", X"70", X"66", X"70", X"72", X"77", X"77", X"76", X"76", X"79", X"74", X"76", X"76", X"76", X"6f", X"72", X"6e", X"6e", X"72", X"6d", X"74", X"6c", X"6d", X"71", X"73", X"66", X"66", X"62", X"64", X"64", X"67", X"67", X"5c", X"59", X"32", X"18", X"07", X"03", X"02", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"08", X"03", X"01", X"07", X"13", X"12", X"4d", X"5b", X"64", X"60", X"6c", X"61", X"65", X"65", X"67", X"64", X"5d", X"65", X"66", X"65", X"66", X"61", X"63", X"62", X"5e", X"5e", X"54", X"56", X"56", X"50", X"52", X"48", X"5a", X"51", X"58", X"5a", X"54", X"5b", X"5b", X"56", X"59", X"4f", X"58", X"59", X"5a", X"55", X"58", X"59", X"57", X"56", X"4f", X"54", X"51", X"4f", X"4b", X"4c", X"47", X"40", X"46", X"45", X"4e", X"3f", X"47", X"44", X"46", X"45", X"43", X"46", X"42", X"3d", X"3e", X"3d", X"41", X"43", X"43", X"3c", X"41", X"3f", X"36", X"3f", X"38", X"3e", X"2f", X"2b", X"36", X"23", X"27", X"29", X"25", X"24", X"1f", X"18", X"13", X"04", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"02", X"06", X"05", X"03", X"0a", X"0e", X"19", X"25", X"29", X"3d", X"35", X"44", X"4b", X"4e", X"5e", X"6f", X"77", X"70", X"5f", X"4f", X"50", X"4d", X"52", X"51", X"56", X"58", X"58", X"4e", X"5a", X"59", X"5a", X"5a", X"53", X"59", X"54", X"53", X"51", X"4a", X"5a", X"5c", X"58", X"4f", X"5d", X"58", X"5e", X"64", X"66", X"6f", X"69", X"67", X"6a", X"6a", X"70", X"6e", X"74", X"6f", X"6f", X"61", X"6f", X"69", X"6b", X"75", X"74", X"6e", X"6f", X"6a", X"72", X"6c", X"6e", X"67", X"6b", X"75", X"69", X"76", X"73", X"6d", X"78", X"73", X"77", X"6d", X"6e", X"6c", X"72", X"73", X"71", X"6b", X"77", X"6c", X"6f", X"67", X"71", X"6f", X"6d", X"6f", X"60", X"68", X"60", X"58", X"68", X"4d", X"34", X"11", X"0d", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"04", X"0a", X"0a", X"0a", X"1c", X"48", X"5e", X"6a", X"62", X"65", X"5c", X"64", X"5e", X"66", X"5a", X"5d", X"5e", X"6a", X"63", X"64", X"5d", X"61", X"64", X"63", X"5f", X"55", X"54", X"55", X"57", X"54", X"52", X"54", X"4f", X"50", X"58", X"53", X"53", X"4e", X"4f", X"50", X"50", X"50", X"4b", X"5d", X"59", X"53", X"56", X"47", X"55", X"4b", X"4f", X"49", X"4e", X"4e", X"4f", X"43", X"3d", X"53", X"48", X"44", X"40", X"49", X"49", X"47", X"4a", X"3a", X"46", X"43", X"3d", X"3f", X"3b", X"40", X"3d", X"3f", X"3f", X"38", X"37", X"44", X"3c", X"36", X"3b", X"33", X"37", X"2f", X"2e", X"29", X"2c", X"22", X"27", X"1d", X"19", X"0e", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"0c", X"05", X"03", X"09", X"06", X"14", X"1c", X"31", X"39", X"43", X"49", X"47", X"42", X"57", X"6a", X"7b", X"83", X"6e", X"64", X"53", X"4e", X"4c", X"55", X"4f", X"53", X"55", X"51", X"59", X"4e", X"57", X"56", X"54", X"54", X"58", X"55", X"57", X"5e", X"55", X"51", X"5a", X"5b", X"5a", X"5c", X"59", X"5e", X"66", X"62", X"5c", X"63", X"6c", X"67", X"6e", X"74", X"62", X"6a", X"65", X"6a", X"69", X"6d", X"69", X"6e", X"73", X"6d", X"6c", X"6e", X"68", X"63", X"69", X"69", X"70", X"6e", X"6a", X"71", X"73", X"6c", X"7c", X"6e", X"73", X"73", X"68", X"6c", X"71", X"67", X"6f", X"6a", X"6b", X"65", X"70", X"6e", X"6a", X"69", X"69", X"63", X"61", X"5b", X"61", X"68", X"64", X"62", X"44", X"12", X"07", X"07", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"07", X"05", X"05", X"04", X"07", X"05", X"10", X"3c", X"5f", X"62", X"6b", X"65", X"5e", X"67", X"66", X"63", X"62", X"60", X"60", X"64", X"63", X"66", X"59", X"5f", X"59", X"5c", X"58", X"56", X"5a", X"48", X"53", X"54", X"51", X"54", X"4d", X"50", X"4b", X"50", X"55", X"58", X"55", X"50", X"4b", X"4f", X"53", X"51", X"52", X"54", X"57", X"56", X"5d", X"49", X"53", X"54", X"4a", X"4e", X"4a", X"50", X"4c", X"50", X"4e", X"4a", X"42", X"4b", X"47", X"47", X"48", X"3e", X"44", X"3b", X"36", X"3b", X"46", X"46", X"3f", X"40", X"37", X"42", X"3d", X"3f", X"3c", X"39", X"3b", X"30", X"30", X"35", X"29", X"25", X"23", X"1e", X"25", X"19", X"11", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"07", X"0a", X"07", X"18", X"24", X"2d", X"37", X"43", X"4c", X"48", X"57", X"5b", X"6c", X"82", X"79", X"5e", X"56", X"4e", X"50", X"5a", X"59", X"58", X"57", X"57", X"53", X"54", X"5d", X"5b", X"5c", X"59", X"50", X"58", X"5b", X"5d", X"52", X"63", X"5b", X"50", X"56", X"5e", X"5a", X"5e", X"63", X"59", X"5f", X"63", X"67", X"68", X"6c", X"6d", X"69", X"6c", X"62", X"60", X"68", X"69", X"6f", X"71", X"70", X"6e", X"6d", X"62", X"6c", X"68", X"6a", X"64", X"65", X"6e", X"74", X"6b", X"71", X"72", X"6f", X"68", X"6e", X"6e", X"65", X"6b", X"66", X"6a", X"6d", X"65", X"6c", X"6f", X"67", X"6d", X"6a", X"6a", X"68", X"68", X"69", X"6b", X"66", X"62", X"99", X"a0", X"53", X"17", X"06", X"03", X"01", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"05", X"02", X"06", X"07", X"11", X"3f", X"58", X"5a", X"60", X"5d", X"5e", X"65", X"59", X"62", X"5f", X"65", X"62", X"69", X"60", X"57", X"58", X"5b", X"4f", X"58", X"53", X"57", X"51", X"53", X"4a", X"49", X"56", X"51", X"53", X"54", X"51", X"53", X"50", X"4b", X"4d", X"44", X"4b", X"45", X"46", X"50", X"4f", X"56", X"54", X"4c", X"50", X"4a", X"55", X"4c", X"3f", X"42", X"50", X"4f", X"4f", X"50", X"46", X"4b", X"4e", X"3e", X"47", X"49", X"44", X"44", X"3a", X"3e", X"3d", X"42", X"40", X"44", X"46", X"39", X"44", X"41", X"3d", X"40", X"40", X"3a", X"38", X"36", X"35", X"2e", X"2c", X"2e", X"2b", X"19", X"1c", X"20", X"0d", X"12", X"08", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"0c", X"14", X"14", X"31", X"3d", X"44", X"4e", X"41", X"54", X"55", X"64", X"70", X"7b", X"6c", X"56", X"53", X"51", X"4a", X"54", X"54", X"56", X"50", X"53", X"56", X"4e", X"55", X"58", X"4e", X"58", X"5c", X"53", X"52", X"53", X"54", X"57", X"50", X"55", X"56", X"57", X"56", X"54", X"54", X"62", X"59", X"62", X"62", X"66", X"6c", X"66", X"6a", X"62", X"65", X"68", X"65", X"6a", X"6e", X"6a", X"6e", X"69", X"67", X"6e", X"5b", X"69", X"6a", X"66", X"69", X"66", X"61", X"6c", X"69", X"6f", X"69", X"6e", X"6b", X"6a", X"65", X"67", X"5e", X"62", X"6b", X"6d", X"79", X"6d", X"6c", X"65", X"6b", X"6a", X"65", X"5d", X"62", X"62", X"67", X"a2", X"b1", X"59", X"1f", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"06", X"06", X"05", X"0d", X"39", X"56", X"60", X"63", X"62", X"5e", X"5f", X"5a", X"61", X"64", X"5e", X"5e", X"63", X"5c", X"5e", X"59", X"57", X"5e", X"54", X"4a", X"50", X"52", X"4f", X"4b", X"50", X"50", X"53", X"52", X"56", X"54", X"54", X"4f", X"51", X"4d", X"4b", X"4e", X"47", X"46", X"4d", X"4b", X"4a", X"4c", X"4b", X"54", X"47", X"51", X"4f", X"47", X"45", X"49", X"4b", X"4e", X"50", X"47", X"4a", X"4d", X"46", X"4a", X"47", X"38", X"38", X"3c", X"43", X"3f", X"3e", X"43", X"3c", X"3d", X"3e", X"3d", X"3c", X"33", X"39", X"39", X"35", X"3a", X"27", X"2c", X"31", X"2c", X"26", X"20", X"1a", X"23", X"11", X"15", X"13", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"0a", X"06", X"13", X"0d", X"1a", X"29", X"2f", X"44", X"49", X"4d", X"4d", X"53", X"5a", X"65", X"68", X"5e", X"52", X"57", X"4c", X"52", X"5a", X"55", X"50", X"59", X"51", X"59", X"55", X"55", X"57", X"52", X"52", X"5a", X"5e", X"53", X"5d", X"53", X"50", X"57", X"55", X"58", X"57", X"56", X"57", X"51", X"59", X"61", X"54", X"5d", X"66", X"64", X"62", X"5f", X"62", X"66", X"69", X"6e", X"6f", X"6c", X"6b", X"67", X"6f", X"69", X"65", X"63", X"65", X"65", X"64", X"65", X"69", X"62", X"6a", X"6e", X"69", X"5f", X"68", X"6a", X"63", X"63", X"66", X"5c", X"65", X"6a", X"66", X"6a", X"61", X"70", X"6d", X"6c", X"65", X"63", X"5f", X"64", X"5f", X"65", X"82", X"6b", X"3d", X"18", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"07", X"09", X"05", X"03", X"02", X"0e", X"08", X"0b", X"34", X"4f", X"56", X"5c", X"5f", X"62", X"5d", X"5f", X"65", X"65", X"62", X"5d", X"5f", X"52", X"56", X"50", X"5c", X"53", X"54", X"52", X"4e", X"4e", X"51", X"4b", X"4f", X"4d", X"50", X"53", X"58", X"53", X"4f", X"50", X"4c", X"55", X"4b", X"51", X"49", X"45", X"49", X"49", X"4c", X"51", X"4b", X"53", X"4a", X"46", X"55", X"4f", X"48", X"43", X"47", X"50", X"45", X"55", X"56", X"49", X"46", X"43", X"4b", X"3c", X"42", X"41", X"3a", X"3d", X"45", X"46", X"3d", X"42", X"47", X"47", X"3e", X"3a", X"35", X"39", X"3d", X"33", X"3d", X"2d", X"31", X"2c", X"21", X"24", X"16", X"22", X"1b", X"17", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"05", X"03", X"00", X"06", X"08", X"11", X"13", X"24", X"24", X"39", X"50", X"4d", X"52", X"50", X"4f", X"58", X"58", X"58", X"57", X"4c", X"4b", X"5a", X"4f", X"5a", X"54", X"4d", X"51", X"57", X"55", X"52", X"59", X"55", X"55", X"59", X"50", X"50", X"54", X"5e", X"58", X"54", X"57", X"56", X"50", X"54", X"56", X"52", X"5b", X"54", X"64", X"58", X"5b", X"5e", X"57", X"60", X"5b", X"64", X"65", X"60", X"6f", X"69", X"68", X"6c", X"61", X"64", X"68", X"63", X"6c", X"66", X"69", X"6b", X"64", X"5e", X"66", X"60", X"6b", X"67", X"60", X"5e", X"5c", X"5b", X"66", X"5e", X"63", X"69", X"66", X"66", X"69", X"6e", X"6c", X"6a", X"66", X"5e", X"68", X"60", X"5f", X"65", X"6a", X"57", X"39", X"12", X"0c", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"0f", X"06", X"06", X"0a", X"30", X"5e", X"5d", X"5e", X"5e", X"5d", X"5c", X"5d", X"65", X"5b", X"5c", X"5a", X"60", X"56", X"58", X"52", X"54", X"5b", X"51", X"52", X"4f", X"4c", X"53", X"48", X"52", X"54", X"51", X"49", X"52", X"4c", X"46", X"51", X"4b", X"51", X"4a", X"46", X"4a", X"4c", X"4e", X"51", X"4c", X"4e", X"48", X"50", X"4b", X"4c", X"4d", X"45", X"46", X"4c", X"4d", X"48", X"4a", X"49", X"4a", X"4b", X"4a", X"48", X"45", X"3e", X"3d", X"43", X"45", X"42", X"3e", X"39", X"43", X"3f", X"46", X"3e", X"40", X"39", X"45", X"34", X"3e", X"38", X"2f", X"31", X"30", X"2a", X"22", X"1f", X"1a", X"1b", X"18", X"09", X"09", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"11", X"10", X"12", X"27", X"33", X"4e", X"57", X"57", X"57", X"4f", X"56", X"52", X"4d", X"4c", X"56", X"5d", X"4b", X"59", X"55", X"53", X"48", X"50", X"5d", X"56", X"54", X"5a", X"58", X"51", X"53", X"55", X"56", X"4a", X"57", X"54", X"51", X"50", X"51", X"56", X"55", X"4f", X"53", X"51", X"5a", X"57", X"54", X"5c", X"4d", X"5b", X"5c", X"60", X"5f", X"61", X"58", X"58", X"60", X"60", X"64", X"63", X"5f", X"68", X"60", X"5f", X"6a", X"65", X"62", X"63", X"5f", X"5f", X"66", X"5a", X"62", X"64", X"63", X"60", X"5f", X"60", X"5d", X"62", X"62", X"65", X"63", X"6b", X"6f", X"6e", X"6a", X"62", X"5b", X"58", X"5b", X"5e", X"61", X"5d", X"51", X"38", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"08", X"09", X"29", X"4a", X"57", X"5c", X"5d", X"5d", X"5b", X"57", X"56", X"59", X"60", X"58", X"56", X"5a", X"54", X"4b", X"51", X"4b", X"4b", X"4e", X"47", X"4b", X"4b", X"4a", X"50", X"4d", X"52", X"45", X"4b", X"45", X"46", X"44", X"4f", X"43", X"45", X"49", X"46", X"42", X"42", X"44", X"42", X"43", X"4f", X"41", X"4b", X"48", X"4f", X"44", X"49", X"4b", X"42", X"45", X"4a", X"41", X"46", X"44", X"44", X"44", X"42", X"3e", X"3d", X"43", X"3b", X"3a", X"43", X"41", X"45", X"4b", X"3f", X"40", X"44", X"3c", X"40", X"34", X"38", X"35", X"3a", X"2d", X"2b", X"23", X"20", X"1e", X"1d", X"1a", X"1b", X"11", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"0a", X"13", X"23", X"31", X"44", X"4e", X"56", X"59", X"54", X"56", X"4d", X"4b", X"50", X"51", X"53", X"4e", X"50", X"49", X"57", X"55", X"57", X"61", X"4c", X"52", X"56", X"53", X"4d", X"5c", X"4e", X"58", X"54", X"54", X"60", X"4d", X"4e", X"5d", X"59", X"58", X"4f", X"52", X"58", X"54", X"56", X"53", X"4f", X"56", X"4d", X"57", X"59", X"5b", X"64", X"5b", X"64", X"5e", X"59", X"63", X"60", X"64", X"65", X"62", X"63", X"63", X"5c", X"6c", X"65", X"65", X"65", X"67", X"64", X"5c", X"5c", X"5f", X"64", X"5e", X"5e", X"5d", X"58", X"5b", X"66", X"69", X"66", X"77", X"65", X"63", X"5f", X"57", X"5a", X"65", X"5f", X"5b", X"56", X"5d", X"3a", X"1a", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"08", X"0b", X"00", X"06", X"05", X"0a", X"27", X"4b", X"50", X"63", X"57", X"56", X"59", X"57", X"5b", X"62", X"4c", X"56", X"58", X"5a", X"4d", X"51", X"47", X"48", X"4e", X"4d", X"52", X"4d", X"4d", X"52", X"47", X"46", X"4d", X"4b", X"43", X"4a", X"48", X"45", X"45", X"44", X"4a", X"4d", X"4b", X"48", X"45", X"4b", X"48", X"40", X"47", X"44", X"47", X"50", X"4d", X"4b", X"44", X"47", X"4f", X"4b", X"47", X"49", X"47", X"47", X"47", X"4a", X"3b", X"48", X"3e", X"39", X"3f", X"38", X"42", X"41", X"46", X"42", X"44", X"3b", X"3b", X"35", X"33", X"3a", X"33", X"39", X"30", X"2d", X"39", X"2a", X"26", X"1f", X"11", X"1c", X"0f", X"11", X"07", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"16", X"23", X"27", X"3c", X"4b", X"54", X"5c", X"50", X"47", X"4e", X"53", X"4d", X"58", X"54", X"5b", X"51", X"50", X"55", X"51", X"4f", X"58", X"53", X"54", X"59", X"54", X"52", X"50", X"55", X"4c", X"53", X"57", X"53", X"57", X"54", X"53", X"55", X"53", X"4f", X"54", X"58", X"5c", X"50", X"50", X"52", X"4b", X"54", X"52", X"53", X"58", X"59", X"5a", X"54", X"57", X"5b", X"5d", X"60", X"64", X"63", X"5f", X"61", X"65", X"63", X"65", X"5d", X"67", X"63", X"5b", X"64", X"61", X"5d", X"61", X"50", X"62", X"58", X"69", X"5f", X"62", X"64", X"6a", X"6a", X"68", X"64", X"62", X"61", X"5e", X"5f", X"5e", X"62", X"5e", X"5a", X"50", X"3b", X"11", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"0e", X"22", X"4f", X"59", X"58", X"5f", X"5d", X"57", X"50", X"59", X"5a", X"51", X"52", X"55", X"47", X"54", X"47", X"4a", X"4f", X"44", X"4e", X"51", X"49", X"4f", X"48", X"54", X"4c", X"4d", X"4a", X"49", X"4e", X"49", X"44", X"4a", X"49", X"4a", X"45", X"44", X"4c", X"45", X"4c", X"48", X"41", X"47", X"4a", X"46", X"4a", X"50", X"43", X"41", X"4d", X"48", X"47", X"4e", X"48", X"4a", X"4d", X"48", X"42", X"4c", X"47", X"43", X"44", X"43", X"45", X"3e", X"46", X"46", X"3f", X"47", X"3f", X"35", X"3c", X"44", X"34", X"3a", X"33", X"39", X"26", X"2a", X"23", X"26", X"23", X"1a", X"15", X"10", X"18", X"0e", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"07", X"1a", X"1e", X"24", X"42", X"4f", X"54", X"5b", X"4e", X"4b", X"4a", X"4f", X"4e", X"50", X"51", X"52", X"55", X"58", X"55", X"4c", X"52", X"55", X"53", X"50", X"51", X"53", X"4d", X"54", X"4d", X"56", X"4e", X"51", X"56", X"53", X"52", X"53", X"58", X"52", X"55", X"50", X"4c", X"52", X"4e", X"57", X"50", X"47", X"4f", X"4c", X"4b", X"4e", X"4d", X"54", X"55", X"59", X"58", X"52", X"56", X"58", X"5f", X"5d", X"57", X"59", X"63", X"54", X"5c", X"5e", X"58", X"61", X"5e", X"63", X"64", X"5d", X"58", X"5f", X"59", X"59", X"5d", X"5f", X"62", X"62", X"67", X"5f", X"5c", X"58", X"54", X"53", X"52", X"58", X"57", X"55", X"4e", X"3e", X"11", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"1b", X"50", X"4b", X"5e", X"52", X"4b", X"4e", X"47", X"56", X"51", X"4f", X"52", X"4e", X"4e", X"43", X"46", X"45", X"47", X"4f", X"47", X"43", X"46", X"43", X"4c", X"4f", X"49", X"4c", X"47", X"42", X"43", X"45", X"40", X"40", X"45", X"45", X"43", X"3c", X"46", X"47", X"42", X"45", X"4a", X"3e", X"46", X"43", X"3f", X"4d", X"47", X"50", X"53", X"51", X"50", X"4d", X"4e", X"51", X"44", X"51", X"44", X"41", X"43", X"3d", X"43", X"3f", X"3a", X"44", X"3e", X"46", X"3d", X"3e", X"40", X"41", X"3a", X"3c", X"33", X"31", X"33", X"30", X"2d", X"26", X"24", X"23", X"17", X"10", X"0d", X"0e", X"0c", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0b", X"00", X"09", X"0c", X"16", X"1f", X"35", X"3e", X"5b", X"56", X"4c", X"4d", X"4c", X"53", X"4e", X"54", X"4e", X"50", X"4b", X"51", X"4e", X"5b", X"57", X"50", X"52", X"58", X"55", X"52", X"58", X"4c", X"55", X"4a", X"4e", X"56", X"4e", X"4e", X"54", X"50", X"4b", X"54", X"51", X"4f", X"57", X"4f", X"5a", X"53", X"4d", X"4b", X"4f", X"4f", X"4d", X"55", X"4b", X"55", X"59", X"5c", X"56", X"54", X"56", X"5b", X"5e", X"5b", X"5b", X"5e", X"5e", X"5d", X"57", X"5a", X"5b", X"5a", X"59", X"5a", X"5c", X"64", X"5e", X"59", X"56", X"5f", X"57", X"5f", X"5e", X"61", X"6c", X"5e", X"57", X"5d", X"4f", X"4b", X"4b", X"55", X"4f", X"4d", X"5a", X"33", X"19", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0b", X"06", X"05", X"07", X"1e", X"45", X"55", X"53", X"49", X"48", X"53", X"49", X"5a", X"50", X"4d", X"4e", X"49", X"49", X"4d", X"44", X"3e", X"44", X"3c", X"49", X"4d", X"48", X"4d", X"4d", X"4b", X"47", X"4c", X"4e", X"44", X"49", X"48", X"3d", X"46", X"49", X"3d", X"46", X"46", X"48", X"3e", X"43", X"3d", X"41", X"40", X"45", X"43", X"4a", X"4d", X"4d", X"4c", X"51", X"57", X"55", X"55", X"49", X"52", X"52", X"4f", X"46", X"48", X"44", X"4d", X"45", X"3f", X"3c", X"44", X"3e", X"39", X"3f", X"40", X"3a", X"3b", X"33", X"3c", X"35", X"36", X"33", X"30", X"28", X"2b", X"24", X"1e", X"16", X"14", X"13", X"08", X"0f", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"02", X"08", X"10", X"17", X"16", X"23", X"3c", X"45", X"49", X"44", X"4b", X"45", X"4d", X"5b", X"52", X"4e", X"5a", X"57", X"59", X"55", X"59", X"59", X"58", X"4e", X"52", X"55", X"4d", X"55", X"52", X"4c", X"4f", X"4d", X"50", X"55", X"4f", X"54", X"4e", X"52", X"53", X"58", X"51", X"4f", X"50", X"45", X"51", X"4f", X"4d", X"4f", X"4f", X"4a", X"51", X"4f", X"47", X"4d", X"53", X"4e", X"49", X"55", X"59", X"54", X"52", X"58", X"56", X"5e", X"5f", X"56", X"5b", X"5a", X"63", X"56", X"5a", X"60", X"5d", X"65", X"5e", X"5b", X"5f", X"5a", X"62", X"6a", X"5d", X"64", X"5c", X"5b", X"54", X"52", X"52", X"5e", X"52", X"49", X"51", X"48", X"36", X"0f", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0d", X"06", X"09", X"0a", X"1b", X"41", X"4c", X"58", X"53", X"4d", X"48", X"48", X"4f", X"4c", X"45", X"4c", X"52", X"52", X"51", X"48", X"41", X"45", X"4d", X"45", X"49", X"47", X"47", X"4d", X"51", X"58", X"4e", X"4c", X"4d", X"46", X"48", X"3a", X"44", X"41", X"45", X"48", X"43", X"49", X"45", X"40", X"42", X"43", X"47", X"49", X"4a", X"4f", X"54", X"4e", X"56", X"5a", X"62", X"5a", X"54", X"5b", X"4a", X"4d", X"46", X"4a", X"46", X"4d", X"4f", X"46", X"48", X"47", X"46", X"4b", X"41", X"3b", X"40", X"41", X"38", X"37", X"39", X"32", X"34", X"36", X"2f", X"2b", X"2a", X"27", X"22", X"19", X"18", X"18", X"12", X"0e", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"02", X"06", X"0d", X"0e", X"11", X"22", X"2b", X"38", X"43", X"47", X"44", X"48", X"4c", X"4f", X"56", X"52", X"56", X"55", X"56", X"4d", X"55", X"56", X"50", X"4b", X"5b", X"4f", X"48", X"51", X"58", X"4b", X"50", X"55", X"54", X"48", X"46", X"4d", X"4f", X"4c", X"4c", X"52", X"48", X"46", X"4e", X"4c", X"4b", X"4c", X"53", X"4d", X"4b", X"4a", X"4c", X"4c", X"4f", X"4f", X"4b", X"4c", X"52", X"4d", X"54", X"52", X"50", X"51", X"55", X"53", X"4e", X"4a", X"53", X"59", X"52", X"5e", X"59", X"61", X"5d", X"5a", X"4f", X"56", X"5e", X"57", X"5c", X"61", X"5b", X"5c", X"5a", X"4b", X"55", X"59", X"58", X"49", X"4e", X"50", X"48", X"54", X"36", X"0f", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"06", X"0d", X"05", X"11", X"3e", X"4e", X"4f", X"4f", X"4c", X"51", X"4c", X"52", X"4c", X"46", X"4a", X"4b", X"44", X"46", X"44", X"4c", X"49", X"47", X"52", X"4f", X"47", X"4b", X"48", X"50", X"57", X"51", X"52", X"50", X"45", X"40", X"46", X"45", X"45", X"44", X"3c", X"47", X"3b", X"44", X"42", X"3d", X"45", X"42", X"43", X"41", X"48", X"54", X"4e", X"53", X"5b", X"4f", X"54", X"52", X"4e", X"4d", X"3d", X"42", X"41", X"45", X"3f", X"50", X"40", X"46", X"3c", X"3d", X"45", X"41", X"3c", X"38", X"3d", X"3b", X"36", X"35", X"2a", X"35", X"2e", X"31", X"2b", X"29", X"26", X"20", X"1d", X"17", X"12", X"0c", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"03", X"06", X"05", X"0b", X"17", X"22", X"25", X"33", X"37", X"40", X"45", X"50", X"4e", X"53", X"52", X"53", X"55", X"56", X"51", X"54", X"54", X"4b", X"54", X"4e", X"4d", X"50", X"4c", X"4a", X"4d", X"4b", X"4e", X"4f", X"4e", X"4d", X"46", X"4d", X"50", X"4f", X"54", X"50", X"43", X"48", X"53", X"47", X"4f", X"4d", X"42", X"52", X"41", X"4e", X"43", X"4d", X"4b", X"49", X"48", X"51", X"4f", X"4c", X"50", X"42", X"4a", X"55", X"4c", X"4c", X"58", X"54", X"5e", X"52", X"5a", X"55", X"4d", X"5a", X"57", X"5c", X"5f", X"60", X"60", X"60", X"5a", X"58", X"5c", X"56", X"54", X"58", X"4e", X"57", X"56", X"54", X"52", X"50", X"4d", X"4c", X"39", X"19", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"12", X"3e", X"48", X"55", X"4f", X"43", X"49", X"49", X"50", X"42", X"42", X"41", X"45", X"4e", X"45", X"4a", X"41", X"4d", X"4e", X"48", X"46", X"52", X"5c", X"52", X"54", X"45", X"54", X"4d", X"4e", X"45", X"42", X"4c", X"3c", X"40", X"44", X"44", X"49", X"43", X"4a", X"44", X"41", X"3d", X"49", X"40", X"4a", X"4b", X"47", X"49", X"45", X"50", X"52", X"51", X"54", X"41", X"47", X"41", X"47", X"44", X"4a", X"46", X"40", X"48", X"45", X"40", X"43", X"45", X"3e", X"3f", X"38", X"33", X"37", X"2f", X"38", X"33", X"35", X"34", X"2f", X"31", X"25", X"2d", X"13", X"13", X"1a", X"0f", X"03", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"08", X"04", X"0f", X"1c", X"1f", X"2a", X"35", X"3d", X"47", X"49", X"50", X"53", X"51", X"51", X"51", X"56", X"52", X"4d", X"54", X"53", X"4f", X"50", X"54", X"51", X"49", X"53", X"54", X"5a", X"4d", X"4d", X"4d", X"4f", X"4f", X"4d", X"50", X"43", X"47", X"4a", X"57", X"52", X"4d", X"47", X"4b", X"48", X"55", X"49", X"4d", X"51", X"48", X"49", X"50", X"4c", X"50", X"49", X"50", X"52", X"50", X"50", X"51", X"4e", X"4d", X"50", X"51", X"5b", X"54", X"58", X"5a", X"50", X"54", X"5b", X"54", X"58", X"5a", X"5e", X"61", X"57", X"5c", X"5c", X"5f", X"59", X"56", X"56", X"50", X"51", X"53", X"4d", X"4f", X"4e", X"4a", X"46", X"38", X"1c", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"07", X"1a", X"34", X"44", X"4d", X"4e", X"47", X"46", X"45", X"4f", X"48", X"47", X"47", X"44", X"45", X"4b", X"41", X"48", X"4a", X"4b", X"50", X"4f", X"53", X"54", X"51", X"4e", X"4a", X"57", X"4f", X"4b", X"4b", X"42", X"45", X"4d", X"4c", X"44", X"44", X"43", X"3e", X"45", X"42", X"47", X"44", X"47", X"48", X"46", X"49", X"43", X"3f", X"47", X"4c", X"43", X"4b", X"3f", X"4d", X"43", X"41", X"48", X"42", X"44", X"3f", X"44", X"48", X"47", X"48", X"3d", X"45", X"41", X"42", X"45", X"3c", X"3c", X"2b", X"37", X"35", X"35", X"2d", X"2f", X"27", X"27", X"20", X"19", X"18", X"17", X"11", X"0d", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"02", X"06", X"05", X"05", X"0b", X"13", X"1d", X"25", X"2b", X"38", X"46", X"4b", X"4a", X"50", X"4d", X"51", X"5a", X"50", X"53", X"52", X"4a", X"4e", X"4a", X"4b", X"49", X"4e", X"49", X"49", X"52", X"46", X"4c", X"51", X"56", X"4f", X"49", X"4a", X"4c", X"4e", X"4a", X"4c", X"4a", X"4c", X"49", X"45", X"4b", X"4b", X"50", X"47", X"3e", X"49", X"45", X"45", X"41", X"49", X"4d", X"51", X"50", X"48", X"4e", X"4b", X"56", X"42", X"52", X"4f", X"4b", X"4e", X"51", X"53", X"55", X"55", X"59", X"5b", X"5a", X"5f", X"54", X"56", X"55", X"59", X"5f", X"59", X"54", X"58", X"51", X"52", X"5b", X"50", X"4a", X"4d", X"50", X"52", X"4a", X"47", X"3e", X"14", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"07", X"3a", X"49", X"4d", X"46", X"47", X"46", X"41", X"44", X"42", X"45", X"44", X"45", X"49", X"46", X"47", X"44", X"4a", X"51", X"52", X"50", X"53", X"5a", X"56", X"4f", X"43", X"50", X"47", X"55", X"50", X"3e", X"4a", X"48", X"47", X"49", X"4a", X"44", X"43", X"46", X"3f", X"40", X"42", X"37", X"45", X"41", X"46", X"3e", X"3e", X"3f", X"3f", X"41", X"47", X"3d", X"3d", X"36", X"3b", X"44", X"42", X"44", X"3f", X"42", X"42", X"3e", X"3a", X"3a", X"3d", X"44", X"3b", X"35", X"37", X"34", X"35", X"2f", X"3d", X"35", X"35", X"2e", X"2d", X"30", X"1d", X"20", X"1b", X"12", X"0c", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"0d", X"0e", X"06", X"15", X"18", X"1d", X"3c", X"3a", X"47", X"45", X"4a", X"4e", X"4f", X"55", X"50", X"52", X"57", X"4f", X"48", X"4b", X"48", X"54", X"4d", X"4b", X"43", X"4b", X"46", X"42", X"4b", X"47", X"47", X"4d", X"4c", X"3e", X"4f", X"4c", X"45", X"4e", X"4b", X"54", X"48", X"49", X"4c", X"47", X"48", X"4f", X"43", X"40", X"48", X"4a", X"45", X"47", X"4a", X"46", X"4e", X"4f", X"48", X"4e", X"4b", X"46", X"4c", X"49", X"4f", X"56", X"4b", X"56", X"52", X"58", X"50", X"4d", X"5d", X"5f", X"52", X"5b", X"60", X"55", X"59", X"5a", X"5a", X"59", X"50", X"55", X"4f", X"4d", X"4f", X"4c", X"4b", X"4d", X"41", X"3e", X"1d", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"0c", X"36", X"47", X"50", X"4e", X"4b", X"46", X"48", X"3b", X"3d", X"43", X"43", X"4c", X"49", X"46", X"4a", X"57", X"4f", X"57", X"50", X"52", X"45", X"52", X"42", X"4e", X"40", X"48", X"44", X"4e", X"50", X"46", X"4f", X"49", X"42", X"4b", X"3c", X"48", X"4b", X"41", X"45", X"37", X"43", X"40", X"3d", X"3e", X"44", X"3b", X"3a", X"38", X"3d", X"3f", X"3f", X"3e", X"37", X"3f", X"3d", X"41", X"42", X"4c", X"3e", X"34", X"37", X"3b", X"3b", X"41", X"3a", X"38", X"3e", X"39", X"39", X"36", X"30", X"35", X"35", X"33", X"38", X"36", X"28", X"24", X"1b", X"1a", X"15", X"11", X"06", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0e", X"08", X"09", X"0b", X"14", X"22", X"2e", X"38", X"46", X"4c", X"41", X"54", X"4d", X"49", X"55", X"51", X"4d", X"4d", X"50", X"54", X"48", X"54", X"49", X"46", X"4d", X"4e", X"50", X"4a", X"46", X"46", X"48", X"45", X"47", X"54", X"4a", X"4a", X"45", X"49", X"4b", X"48", X"48", X"45", X"48", X"41", X"4c", X"4a", X"40", X"4d", X"49", X"47", X"4a", X"4e", X"4a", X"52", X"47", X"45", X"42", X"4a", X"48", X"4c", X"51", X"4d", X"51", X"59", X"47", X"51", X"54", X"47", X"53", X"56", X"5a", X"54", X"56", X"53", X"58", X"5e", X"5f", X"55", X"5b", X"4e", X"5d", X"50", X"55", X"51", X"52", X"53", X"53", X"54", X"4d", X"40", X"1a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"29", X"49", X"4d", X"4d", X"46", X"47", X"47", X"47", X"46", X"3c", X"44", X"44", X"47", X"4f", X"49", X"4c", X"48", X"4b", X"52", X"49", X"43", X"4e", X"43", X"4c", X"46", X"47", X"4f", X"4f", X"4b", X"48", X"41", X"46", X"41", X"45", X"39", X"41", X"47", X"3e", X"3a", X"42", X"36", X"44", X"48", X"3d", X"3d", X"40", X"3b", X"3e", X"40", X"38", X"3b", X"43", X"3f", X"41", X"44", X"42", X"3d", X"3c", X"3c", X"42", X"38", X"3e", X"37", X"39", X"3d", X"43", X"41", X"3a", X"3d", X"34", X"33", X"34", X"39", X"37", X"33", X"38", X"23", X"30", X"22", X"19", X"19", X"0b", X"0b", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"0a", X"05", X"06", X"06", X"07", X"15", X"19", X"1b", X"24", X"2d", X"3f", X"49", X"46", X"4f", X"52", X"46", X"48", X"49", X"52", X"4e", X"52", X"49", X"49", X"4b", X"4c", X"4f", X"47", X"46", X"49", X"4d", X"49", X"4e", X"46", X"44", X"4c", X"47", X"4b", X"47", X"45", X"4e", X"49", X"48", X"46", X"46", X"4e", X"3e", X"48", X"47", X"43", X"49", X"46", X"40", X"4c", X"4d", X"4a", X"4d", X"4d", X"49", X"42", X"4a", X"49", X"49", X"48", X"43", X"4e", X"52", X"58", X"53", X"55", X"55", X"52", X"50", X"53", X"60", X"5b", X"60", X"60", X"64", X"5b", X"51", X"60", X"51", X"4e", X"56", X"5c", X"58", X"52", X"4e", X"50", X"48", X"45", X"41", X"1f", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0c", X"31", X"48", X"49", X"51", X"45", X"45", X"3f", X"43", X"49", X"43", X"46", X"42", X"4d", X"4b", X"54", X"54", X"53", X"50", X"44", X"46", X"40", X"42", X"45", X"41", X"45", X"4c", X"53", X"53", X"4a", X"40", X"45", X"3d", X"3c", X"3c", X"4a", X"41", X"43", X"3f", X"3c", X"35", X"38", X"31", X"3f", X"3a", X"37", X"44", X"2e", X"3c", X"3a", X"39", X"40", X"3d", X"3c", X"3e", X"3b", X"39", X"3f", X"3f", X"3c", X"3d", X"3f", X"39", X"36", X"3a", X"44", X"41", X"38", X"3a", X"3c", X"30", X"30", X"3e", X"36", X"32", X"31", X"35", X"2b", X"24", X"1b", X"1a", X"17", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"09", X"05", X"0a", X"10", X"0e", X"1a", X"18", X"27", X"37", X"39", X"45", X"47", X"4e", X"50", X"4b", X"4a", X"51", X"4e", X"4c", X"48", X"4f", X"4a", X"45", X"45", X"44", X"48", X"47", X"4b", X"44", X"4a", X"41", X"4e", X"46", X"43", X"44", X"49", X"41", X"43", X"46", X"46", X"47", X"42", X"48", X"48", X"4f", X"49", X"3f", X"44", X"45", X"4a", X"48", X"4b", X"48", X"42", X"3c", X"4d", X"49", X"42", X"43", X"46", X"52", X"39", X"55", X"47", X"44", X"52", X"4b", X"57", X"51", X"4f", X"54", X"53", X"50", X"5a", X"57", X"58", X"5d", X"53", X"56", X"54", X"53", X"51", X"48", X"52", X"53", X"52", X"4a", X"4b", X"41", X"3c", X"17", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"28", X"42", X"49", X"44", X"3f", X"41", X"3e", X"48", X"43", X"46", X"47", X"4a", X"4c", X"4a", X"46", X"54", X"4f", X"53", X"52", X"53", X"3e", X"45", X"47", X"4a", X"46", X"4c", X"53", X"50", X"45", X"41", X"3f", X"43", X"45", X"42", X"39", X"35", X"3b", X"38", X"33", X"39", X"36", X"3b", X"37", X"33", X"36", X"39", X"34", X"39", X"3d", X"3c", X"37", X"3c", X"3d", X"39", X"35", X"3d", X"3a", X"35", X"3a", X"32", X"34", X"3f", X"31", X"31", X"3d", X"40", X"43", X"38", X"2d", X"37", X"2e", X"39", X"31", X"36", X"2e", X"31", X"25", X"2e", X"12", X"16", X"0b", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"08", X"0c", X"11", X"15", X"11", X"14", X"1b", X"2e", X"3a", X"44", X"4c", X"4a", X"4a", X"48", X"4a", X"4c", X"4f", X"4e", X"4e", X"48", X"50", X"3f", X"4a", X"4d", X"42", X"4e", X"49", X"4c", X"46", X"44", X"49", X"44", X"46", X"4d", X"47", X"3f", X"45", X"43", X"42", X"41", X"41", X"43", X"47", X"44", X"45", X"4e", X"47", X"47", X"45", X"3e", X"45", X"49", X"49", X"4d", X"4b", X"45", X"43", X"45", X"41", X"4a", X"4a", X"48", X"49", X"45", X"54", X"56", X"54", X"57", X"58", X"50", X"5d", X"5a", X"4e", X"59", X"5b", X"51", X"53", X"51", X"53", X"4a", X"51", X"52", X"59", X"4e", X"4e", X"50", X"4c", X"45", X"41", X"22", X"08", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"16", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"2c", X"44", X"4f", X"4d", X"46", X"45", X"46", X"49", X"45", X"3d", X"3e", X"47", X"47", X"4e", X"4c", X"4d", X"53", X"58", X"56", X"4b", X"42", X"44", X"48", X"4f", X"4e", X"54", X"47", X"4a", X"3e", X"46", X"3d", X"3b", X"38", X"40", X"3d", X"39", X"38", X"2e", X"34", X"3e", X"37", X"37", X"3b", X"38", X"3c", X"3a", X"30", X"32", X"36", X"3d", X"3d", X"3b", X"34", X"3b", X"3c", X"39", X"37", X"3b", X"37", X"33", X"35", X"37", X"3e", X"38", X"41", X"3d", X"3e", X"3b", X"3e", X"40", X"39", X"34", X"3b", X"35", X"2d", X"29", X"32", X"25", X"13", X"11", X"0b", X"0a", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"0b", X"11", X"11", X"16", X"1f", X"24", X"38", X"42", X"49", X"51", X"4f", X"4b", X"4a", X"4c", X"45", X"48", X"46", X"4b", X"4d", X"4f", X"44", X"42", X"47", X"46", X"41", X"42", X"4a", X"44", X"45", X"4a", X"4f", X"46", X"40", X"45", X"48", X"47", X"44", X"43", X"43", X"47", X"43", X"41", X"44", X"45", X"42", X"3c", X"41", X"4a", X"47", X"4d", X"46", X"4a", X"46", X"44", X"47", X"49", X"4a", X"4a", X"48", X"4b", X"49", X"46", X"4d", X"48", X"4b", X"54", X"54", X"57", X"54", X"52", X"56", X"59", X"58", X"51", X"52", X"53", X"4f", X"4b", X"56", X"53", X"4e", X"4d", X"50", X"4f", X"46", X"41", X"3b", X"1e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"02", X"2b", X"3c", X"45", X"51", X"42", X"44", X"3e", X"41", X"44", X"4b", X"47", X"48", X"45", X"4a", X"45", X"4c", X"5a", X"5b", X"4e", X"50", X"46", X"46", X"42", X"49", X"47", X"49", X"3f", X"44", X"3a", X"41", X"42", X"3d", X"33", X"3d", X"40", X"3c", X"3a", X"38", X"34", X"32", X"38", X"35", X"39", X"35", X"3c", X"33", X"40", X"39", X"35", X"3a", X"38", X"38", X"37", X"31", X"39", X"3b", X"3a", X"36", X"33", X"32", X"35", X"38", X"38", X"40", X"40", X"33", X"34", X"3c", X"3b", X"48", X"39", X"3e", X"33", X"32", X"28", X"32", X"2e", X"2e", X"20", X"0d", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0a", X"17", X"13", X"1c", X"24", X"31", X"44", X"49", X"49", X"4b", X"53", X"53", X"4e", X"4c", X"52", X"48", X"47", X"45", X"44", X"42", X"45", X"3e", X"44", X"47", X"45", X"46", X"45", X"41", X"3f", X"49", X"41", X"49", X"4a", X"45", X"3d", X"47", X"40", X"42", X"45", X"46", X"4a", X"42", X"42", X"3a", X"3e", X"44", X"42", X"42", X"44", X"41", X"3e", X"46", X"43", X"4a", X"3a", X"45", X"46", X"43", X"42", X"47", X"41", X"47", X"41", X"4a", X"50", X"50", X"53", X"54", X"4e", X"56", X"51", X"53", X"4c", X"49", X"56", X"4e", X"57", X"4c", X"52", X"53", X"4a", X"4d", X"56", X"4d", X"3f", X"3e", X"24", X"0f", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"25", X"48", X"49", X"47", X"4a", X"47", X"45", X"4a", X"4b", X"46", X"46", X"44", X"47", X"4a", X"52", X"48", X"51", X"4c", X"4e", X"4f", X"48", X"45", X"48", X"3d", X"42", X"46", X"39", X"48", X"3d", X"42", X"3d", X"3a", X"3e", X"41", X"3a", X"39", X"39", X"3b", X"2f", X"33", X"2f", X"32", X"36", X"32", X"3a", X"35", X"38", X"34", X"37", X"3a", X"36", X"36", X"31", X"35", X"3a", X"35", X"2d", X"36", X"37", X"35", X"3f", X"3a", X"39", X"39", X"34", X"32", X"39", X"3a", X"33", X"37", X"34", X"34", X"2b", X"30", X"32", X"28", X"26", X"1d", X"11", X"0f", X"0f", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"04", X"0f", X"08", X"0e", X"12", X"10", X"1c", X"21", X"2d", X"49", X"4c", X"4f", X"4f", X"4b", X"4f", X"50", X"51", X"48", X"4b", X"4e", X"4b", X"4e", X"46", X"49", X"44", X"4a", X"4e", X"43", X"4b", X"43", X"44", X"4b", X"4b", X"3e", X"45", X"49", X"42", X"4e", X"46", X"3d", X"3e", X"40", X"42", X"47", X"4e", X"3e", X"49", X"40", X"43", X"47", X"47", X"4b", X"50", X"4b", X"46", X"3c", X"40", X"40", X"43", X"42", X"44", X"44", X"47", X"40", X"42", X"44", X"4b", X"50", X"4d", X"51", X"55", X"52", X"53", X"4e", X"48", X"52", X"4e", X"44", X"52", X"4e", X"4d", X"4d", X"48", X"4e", X"47", X"53", X"54", X"46", X"3b", X"2a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"1e", X"3c", X"49", X"45", X"45", X"44", X"40", X"50", X"4e", X"44", X"45", X"49", X"45", X"54", X"4a", X"4f", X"51", X"44", X"4b", X"3d", X"3e", X"3c", X"40", X"43", X"3d", X"44", X"3e", X"3d", X"3b", X"3c", X"36", X"38", X"30", X"35", X"32", X"30", X"3e", X"3b", X"3b", X"3f", X"37", X"3e", X"36", X"3b", X"3f", X"31", X"32", X"33", X"31", X"33", X"3a", X"33", X"36", X"35", X"37", X"34", X"33", X"34", X"37", X"32", X"3c", X"33", X"34", X"35", X"37", X"34", X"3c", X"38", X"38", X"3a", X"32", X"37", X"35", X"34", X"36", X"2c", X"22", X"20", X"16", X"08", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"05", X"00", X"0a", X"05", X"06", X"12", X"18", X"11", X"1a", X"2a", X"33", X"4c", X"52", X"4f", X"4b", X"46", X"47", X"4b", X"47", X"4c", X"49", X"4e", X"4a", X"45", X"48", X"43", X"47", X"40", X"4e", X"47", X"3d", X"44", X"44", X"48", X"3e", X"4a", X"47", X"49", X"44", X"4a", X"44", X"49", X"45", X"44", X"3b", X"41", X"49", X"47", X"48", X"42", X"44", X"4c", X"43", X"44", X"4a", X"44", X"47", X"4b", X"41", X"43", X"4b", X"41", X"49", X"43", X"45", X"43", X"48", X"4d", X"45", X"48", X"42", X"4b", X"53", X"57", X"55", X"52", X"57", X"55", X"5d", X"4f", X"4c", X"54", X"4c", X"4c", X"4f", X"49", X"4a", X"4b", X"41", X"31", X"25", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"1f", X"40", X"46", X"4f", X"43", X"4d", X"44", X"53", X"52", X"49", X"3c", X"43", X"45", X"42", X"43", X"43", X"47", X"44", X"38", X"42", X"41", X"41", X"3b", X"46", X"3c", X"43", X"3c", X"3d", X"3b", X"3f", X"36", X"38", X"40", X"38", X"35", X"38", X"37", X"2e", X"38", X"35", X"36", X"38", X"38", X"38", X"33", X"42", X"3d", X"33", X"3c", X"3b", X"35", X"36", X"3f", X"2e", X"34", X"38", X"38", X"3c", X"3b", X"3f", X"39", X"32", X"33", X"3a", X"3e", X"38", X"39", X"38", X"37", X"2e", X"34", X"36", X"36", X"2b", X"28", X"30", X"28", X"28", X"16", X"16", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"09", X"02", X"0f", X"11", X"16", X"1e", X"2c", X"42", X"4d", X"4a", X"4b", X"52", X"40", X"3f", X"43", X"46", X"42", X"4e", X"44", X"45", X"48", X"4d", X"45", X"49", X"48", X"47", X"3c", X"4b", X"42", X"3a", X"49", X"45", X"45", X"47", X"47", X"46", X"49", X"3c", X"46", X"43", X"47", X"3b", X"40", X"41", X"3d", X"43", X"4a", X"44", X"45", X"43", X"41", X"48", X"3e", X"43", X"3f", X"3f", X"4c", X"39", X"40", X"44", X"48", X"49", X"44", X"49", X"4a", X"42", X"47", X"46", X"49", X"51", X"51", X"4d", X"53", X"47", X"4d", X"4d", X"47", X"4f", X"50", X"4b", X"4b", X"4a", X"4f", X"4b", X"46", X"34", X"29", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"16", X"3a", X"46", X"45", X"4c", X"47", X"3e", X"48", X"48", X"41", X"45", X"44", X"35", X"42", X"42", X"39", X"3b", X"35", X"40", X"3e", X"3c", X"43", X"43", X"3b", X"3b", X"3e", X"35", X"42", X"37", X"3d", X"3b", X"36", X"37", X"3a", X"36", X"3c", X"34", X"34", X"33", X"38", X"30", X"36", X"2f", X"3a", X"38", X"35", X"35", X"32", X"3a", X"40", X"37", X"37", X"31", X"35", X"27", X"33", X"32", X"31", X"33", X"31", X"34", X"43", X"35", X"3b", X"4a", X"3d", X"40", X"39", X"38", X"34", X"38", X"32", X"39", X"2e", X"2a", X"30", X"25", X"18", X"14", X"07", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0c", X"09", X"06", X"0c", X"21", X"1e", X"27", X"3c", X"3b", X"4a", X"4a", X"4c", X"4c", X"4c", X"4d", X"48", X"4a", X"41", X"43", X"46", X"3c", X"45", X"3f", X"44", X"4a", X"46", X"44", X"45", X"44", X"4a", X"39", X"46", X"48", X"3c", X"46", X"43", X"42", X"4a", X"3d", X"46", X"40", X"49", X"42", X"45", X"3f", X"45", X"45", X"44", X"3e", X"44", X"41", X"45", X"3c", X"3c", X"43", X"45", X"40", X"46", X"4d", X"41", X"3e", X"42", X"3e", X"44", X"48", X"41", X"45", X"47", X"47", X"44", X"45", X"48", X"51", X"56", X"56", X"4d", X"48", X"4e", X"47", X"52", X"4e", X"4f", X"50", X"41", X"43", X"3a", X"25", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"19", X"3a", X"4a", X"47", X"41", X"4b", X"41", X"4e", X"4a", X"3f", X"43", X"3f", X"3d", X"3e", X"37", X"39", X"3c", X"3b", X"3e", X"3c", X"35", X"3b", X"36", X"41", X"34", X"3b", X"40", X"42", X"36", X"40", X"34", X"3a", X"35", X"33", X"2d", X"39", X"32", X"37", X"38", X"3b", X"36", X"3a", X"39", X"30", X"35", X"31", X"2e", X"2e", X"34", X"30", X"37", X"36", X"33", X"2e", X"36", X"35", X"32", X"38", X"33", X"2e", X"39", X"36", X"3a", X"46", X"4d", X"4b", X"4a", X"3f", X"35", X"2d", X"37", X"2b", X"2b", X"35", X"28", X"29", X"24", X"14", X"1a", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"11", X"09", X"16", X"11", X"21", X"34", X"3f", X"46", X"4a", X"4f", X"46", X"47", X"46", X"48", X"4a", X"50", X"4d", X"44", X"45", X"41", X"4b", X"48", X"45", X"51", X"4c", X"45", X"44", X"46", X"42", X"3f", X"41", X"49", X"43", X"49", X"42", X"47", X"4d", X"47", X"4f", X"3d", X"3e", X"41", X"4b", X"41", X"46", X"46", X"41", X"49", X"3e", X"4a", X"45", X"46", X"3e", X"47", X"41", X"4a", X"43", X"47", X"48", X"41", X"46", X"48", X"3d", X"4b", X"4a", X"3f", X"3f", X"44", X"45", X"48", X"46", X"4c", X"52", X"52", X"4b", X"50", X"4c", X"4c", X"4a", X"49", X"4b", X"4d", X"44", X"41", X"29", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"0c", X"37", X"4c", X"48", X"41", X"45", X"3b", X"46", X"47", X"48", X"38", X"42", X"41", X"3f", X"3b", X"3f", X"45", X"3e", X"3e", X"45", X"3d", X"3c", X"41", X"3e", X"39", X"40", X"3c", X"35", X"45", X"42", X"37", X"3a", X"3e", X"3d", X"33", X"36", X"38", X"36", X"35", X"34", X"33", X"38", X"37", X"3a", X"38", X"41", X"38", X"31", X"3e", X"35", X"39", X"36", X"31", X"2e", X"2a", X"32", X"33", X"35", X"38", X"31", X"33", X"3a", X"39", X"49", X"52", X"4e", X"49", X"41", X"3d", X"3a", X"3a", X"37", X"3e", X"3c", X"2a", X"28", X"18", X"1f", X"13", X"0b", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"06", X"07", X"0c", X"10", X"14", X"1e", X"25", X"32", X"3b", X"45", X"50", X"41", X"41", X"3e", X"44", X"4e", X"50", X"46", X"44", X"49", X"3f", X"45", X"47", X"45", X"47", X"3d", X"48", X"4a", X"42", X"44", X"45", X"3c", X"49", X"40", X"49", X"3d", X"46", X"44", X"43", X"42", X"3a", X"42", X"47", X"3b", X"3e", X"41", X"45", X"3e", X"3e", X"39", X"39", X"42", X"47", X"36", X"45", X"40", X"46", X"45", X"44", X"46", X"46", X"3f", X"34", X"4a", X"3e", X"44", X"49", X"44", X"43", X"45", X"47", X"47", X"4a", X"3c", X"3f", X"43", X"43", X"45", X"4a", X"4e", X"45", X"47", X"42", X"41", X"40", X"26", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"08", X"3e", X"40", X"53", X"49", X"44", X"43", X"47", X"40", X"36", X"3e", X"39", X"3a", X"3c", X"3a", X"34", X"3a", X"30", X"3b", X"3d", X"3f", X"3f", X"3e", X"39", X"35", X"3f", X"35", X"3c", X"39", X"3d", X"3f", X"39", X"36", X"36", X"37", X"2f", X"37", X"36", X"3d", X"3b", X"36", X"34", X"37", X"31", X"38", X"36", X"33", X"32", X"37", X"38", X"32", X"2f", X"2d", X"2b", X"2f", X"27", X"34", X"33", X"35", X"30", X"32", X"39", X"3c", X"3b", X"3d", X"43", X"4a", X"45", X"47", X"38", X"35", X"2f", X"2d", X"32", X"2f", X"2a", X"1e", X"16", X"06", X"02", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"07", X"17", X"0e", X"16", X"1f", X"26", X"2e", X"43", X"3e", X"48", X"47", X"4b", X"51", X"45", X"42", X"4a", X"3d", X"46", X"48", X"47", X"44", X"44", X"4a", X"4e", X"44", X"41", X"42", X"41", X"47", X"46", X"46", X"3f", X"48", X"45", X"44", X"3c", X"40", X"3e", X"44", X"3b", X"40", X"43", X"40", X"3e", X"3e", X"3d", X"42", X"46", X"40", X"49", X"44", X"40", X"3d", X"48", X"43", X"47", X"49", X"38", X"3f", X"41", X"3d", X"46", X"40", X"39", X"3d", X"48", X"43", X"45", X"40", X"44", X"3d", X"49", X"47", X"40", X"41", X"45", X"4b", X"42", X"43", X"48", X"4e", X"42", X"3e", X"33", X"2d", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"10", X"30", X"49", X"4e", X"40", X"41", X"3e", X"39", X"3c", X"3f", X"37", X"35", X"35", X"35", X"3e", X"35", X"39", X"39", X"3a", X"3c", X"3e", X"3d", X"40", X"39", X"3a", X"3b", X"36", X"38", X"45", X"3a", X"3b", X"3d", X"3a", X"3e", X"38", X"36", X"43", X"3b", X"37", X"34", X"38", X"37", X"37", X"31", X"3c", X"30", X"30", X"32", X"3a", X"33", X"35", X"2f", X"32", X"38", X"34", X"37", X"35", X"33", X"32", X"30", X"3a", X"32", X"36", X"3e", X"48", X"3a", X"3c", X"3e", X"43", X"35", X"31", X"38", X"2e", X"2a", X"2b", X"22", X"1a", X"17", X"08", X"09", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"08", X"08", X"0c", X"14", X"1d", X"27", X"41", X"49", X"47", X"49", X"3d", X"49", X"50", X"43", X"49", X"4e", X"4a", X"45", X"41", X"3e", X"3d", X"44", X"3d", X"4d", X"43", X"44", X"4c", X"43", X"4a", X"41", X"43", X"48", X"4d", X"47", X"43", X"42", X"3f", X"45", X"41", X"41", X"49", X"42", X"49", X"47", X"38", X"43", X"44", X"3e", X"43", X"46", X"3d", X"41", X"45", X"44", X"46", X"3b", X"3e", X"41", X"44", X"3b", X"41", X"44", X"45", X"46", X"45", X"3a", X"43", X"4b", X"4b", X"3e", X"46", X"49", X"41", X"48", X"47", X"49", X"41", X"48", X"39", X"46", X"49", X"40", X"3a", X"43", X"29", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"0f", X"38", X"47", X"41", X"45", X"3e", X"38", X"40", X"3d", X"3e", X"3c", X"41", X"33", X"32", X"39", X"3e", X"3f", X"3d", X"42", X"40", X"3a", X"43", X"39", X"3c", X"38", X"41", X"40", X"3d", X"35", X"3f", X"3a", X"36", X"42", X"37", X"36", X"37", X"35", X"32", X"34", X"3a", X"39", X"30", X"32", X"31", X"38", X"31", X"33", X"3a", X"30", X"3d", X"39", X"3a", X"34", X"33", X"2d", X"33", X"36", X"3a", X"3f", X"35", X"35", X"35", X"35", X"39", X"41", X"40", X"43", X"4c", X"45", X"43", X"30", X"31", X"30", X"2c", X"2f", X"30", X"1a", X"17", X"05", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"0a", X"0a", X"0f", X"16", X"1e", X"25", X"34", X"3b", X"44", X"42", X"42", X"46", X"45", X"46", X"44", X"4b", X"45", X"41", X"49", X"47", X"44", X"43", X"4b", X"3e", X"45", X"41", X"48", X"4d", X"41", X"42", X"4e", X"43", X"44", X"40", X"45", X"46", X"3f", X"46", X"47", X"3f", X"3a", X"3b", X"44", X"3e", X"3b", X"45", X"45", X"45", X"3e", X"43", X"33", X"41", X"43", X"3e", X"45", X"38", X"41", X"40", X"46", X"3a", X"3b", X"3f", X"44", X"47", X"40", X"49", X"40", X"3f", X"43", X"38", X"45", X"42", X"38", X"38", X"3a", X"49", X"3f", X"3f", X"40", X"49", X"41", X"43", X"39", X"37", X"2b", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"35", X"3a", X"43", X"45", X"43", X"35", X"44", X"42", X"2e", X"40", X"37", X"42", X"3b", X"37", X"3a", X"34", X"3b", X"36", X"30", X"36", X"33", X"34", X"34", X"36", X"3b", X"33", X"3b", X"36", X"40", X"3c", X"3b", X"39", X"30", X"34", X"37", X"35", X"38", X"36", X"35", X"34", X"33", X"34", X"35", X"32", X"32", X"2f", X"2e", X"35", X"37", X"33", X"35", X"30", X"31", X"39", X"36", X"3c", X"39", X"39", X"34", X"35", X"41", X"39", X"42", X"45", X"4c", X"42", X"45", X"3e", X"30", X"2b", X"2d", X"2d", X"25", X"25", X"26", X"14", X"0d", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"0b", X"0b", X"1b", X"17", X"19", X"2e", X"2e", X"40", X"49", X"47", X"4c", X"48", X"3a", X"41", X"46", X"42", X"38", X"43", X"42", X"3f", X"3c", X"3f", X"44", X"48", X"3a", X"3f", X"41", X"3b", X"46", X"45", X"44", X"42", X"41", X"44", X"3f", X"4b", X"3a", X"43", X"3e", X"40", X"3e", X"40", X"40", X"3e", X"49", X"44", X"40", X"45", X"3b", X"44", X"42", X"43", X"3c", X"43", X"3b", X"43", X"43", X"37", X"3a", X"3c", X"42", X"40", X"43", X"38", X"34", X"3d", X"3b", X"3d", X"3f", X"3e", X"41", X"39", X"3b", X"33", X"3e", X"3f", X"42", X"3c", X"38", X"37", X"36", X"35", X"32", X"23", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"2e", X"3f", X"3b", X"3f", X"3c", X"38", X"3f", X"34", X"38", X"30", X"3b", X"32", X"38", X"36", X"3b", X"3a", X"35", X"3c", X"42", X"3b", X"41", X"3a", X"41", X"37", X"3b", X"38", X"34", X"3a", X"39", X"32", X"38", X"3e", X"3d", X"37", X"38", X"35", X"33", X"2a", X"39", X"30", X"3b", X"31", X"2f", X"36", X"37", X"32", X"2f", X"36", X"37", X"31", X"2b", X"2c", X"2f", X"37", X"3b", X"3a", X"40", X"39", X"3c", X"36", X"3d", X"3d", X"46", X"3d", X"3c", X"40", X"3b", X"34", X"35", X"2d", X"33", X"36", X"34", X"2e", X"1d", X"15", X"07", X"05", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"07", X"07", X"06", X"18", X"1b", X"25", X"2f", X"32", X"3d", X"45", X"4a", X"45", X"42", X"4a", X"48", X"42", X"43", X"44", X"49", X"40", X"49", X"41", X"45", X"3f", X"41", X"45", X"44", X"3e", X"3c", X"48", X"43", X"47", X"40", X"41", X"48", X"3f", X"48", X"42", X"44", X"41", X"39", X"37", X"47", X"3c", X"43", X"41", X"38", X"37", X"45", X"41", X"44", X"45", X"34", X"3e", X"43", X"43", X"45", X"3f", X"45", X"37", X"41", X"3f", X"37", X"3e", X"45", X"3b", X"3c", X"43", X"39", X"3e", X"37", X"43", X"40", X"35", X"3b", X"35", X"35", X"35", X"3d", X"3a", X"40", X"39", X"2f", X"2b", X"0e", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"28", X"42", X"3b", X"44", X"40", X"3d", X"39", X"35", X"3a", X"32", X"3c", X"38", X"39", X"37", X"32", X"36", X"3a", X"39", X"3e", X"36", X"33", X"3e", X"37", X"35", X"3f", X"37", X"3a", X"34", X"44", X"32", X"42", X"40", X"3c", X"3d", X"3b", X"38", X"39", X"2c", X"31", X"32", X"3a", X"33", X"38", X"35", X"31", X"31", X"38", X"3b", X"38", X"31", X"35", X"35", X"3d", X"3d", X"3b", X"3a", X"3a", X"3b", X"37", X"3a", X"42", X"3d", X"4b", X"42", X"44", X"3e", X"3f", X"33", X"34", X"33", X"2f", X"2f", X"25", X"29", X"1f", X"0b", X"0d", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"0b", X"0c", X"16", X"22", X"28", X"2a", X"3a", X"3e", X"41", X"41", X"41", X"45", X"44", X"47", X"48", X"44", X"45", X"44", X"45", X"46", X"3f", X"45", X"41", X"48", X"49", X"44", X"41", X"3b", X"4a", X"41", X"3e", X"45", X"40", X"41", X"38", X"3f", X"3d", X"40", X"3c", X"45", X"3b", X"3c", X"3c", X"3c", X"40", X"3c", X"36", X"3d", X"3b", X"38", X"36", X"3a", X"45", X"3a", X"41", X"48", X"44", X"36", X"41", X"42", X"3f", X"43", X"40", X"47", X"3c", X"42", X"48", X"3e", X"38", X"41", X"40", X"41", X"3b", X"3d", X"36", X"3a", X"39", X"40", X"3b", X"2d", X"36", X"2f", X"2e", X"10", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"0b", X"28", X"3c", X"3f", X"3c", X"37", X"2f", X"34", X"38", X"3a", X"38", X"39", X"31", X"34", X"35", X"32", X"3c", X"3a", X"3c", X"3e", X"3e", X"3e", X"37", X"35", X"39", X"3f", X"30", X"39", X"45", X"39", X"3e", X"35", X"34", X"3e", X"31", X"33", X"3b", X"31", X"3e", X"3c", X"3b", X"3c", X"3b", X"39", X"3b", X"3d", X"34", X"2d", X"3d", X"3b", X"34", X"39", X"30", X"3e", X"3f", X"3b", X"34", X"42", X"40", X"3d", X"47", X"40", X"42", X"43", X"3f", X"3c", X"3c", X"3c", X"32", X"35", X"32", X"37", X"2e", X"2b", X"24", X"1e", X"0d", X"05", X"0c", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"05", X"04", X"14", X"19", X"1c", X"16", X"25", X"39", X"42", X"40", X"40", X"49", X"46", X"49", X"41", X"3f", X"41", X"47", X"3e", X"3a", X"40", X"41", X"43", X"39", X"47", X"3f", X"50", X"43", X"3e", X"3d", X"4b", X"3d", X"44", X"42", X"40", X"45", X"47", X"46", X"39", X"42", X"35", X"39", X"3c", X"3a", X"36", X"39", X"3a", X"3d", X"3e", X"41", X"40", X"39", X"3f", X"3a", X"42", X"3d", X"39", X"41", X"42", X"3b", X"38", X"44", X"47", X"3a", X"40", X"44", X"46", X"42", X"3a", X"3a", X"3a", X"3f", X"34", X"3a", X"35", X"36", X"35", X"2e", X"34", X"33", X"36", X"29", X"27", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"26", X"32", X"42", X"30", X"32", X"32", X"34", X"3d", X"3a", X"3c", X"39", X"34", X"35", X"3c", X"30", X"3c", X"3b", X"32", X"3f", X"3d", X"3a", X"3a", X"38", X"38", X"3c", X"42", X"37", X"3b", X"35", X"39", X"34", X"3b", X"3b", X"39", X"39", X"3b", X"30", X"35", X"36", X"36", X"38", X"33", X"37", X"35", X"36", X"3a", X"3a", X"36", X"3a", X"33", X"32", X"37", X"3b", X"3d", X"34", X"32", X"3f", X"3d", X"41", X"41", X"40", X"44", X"45", X"3e", X"3e", X"3b", X"3a", X"2e", X"30", X"30", X"34", X"2d", X"27", X"17", X"15", X"0d", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"0d", X"14", X"1f", X"20", X"30", X"3b", X"33", X"42", X"41", X"46", X"51", X"46", X"41", X"41", X"41", X"47", X"43", X"40", X"47", X"47", X"3e", X"45", X"36", X"4e", X"43", X"40", X"45", X"40", X"3c", X"45", X"3e", X"39", X"45", X"3d", X"40", X"3e", X"44", X"3f", X"3b", X"3e", X"3b", X"3b", X"3b", X"3b", X"3c", X"3d", X"37", X"35", X"3b", X"40", X"42", X"40", X"3d", X"3c", X"3b", X"3f", X"40", X"37", X"41", X"37", X"3e", X"40", X"40", X"38", X"3c", X"35", X"33", X"3f", X"3e", X"39", X"3a", X"3d", X"39", X"34", X"33", X"35", X"33", X"2b", X"2b", X"2d", X"25", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"09", X"26", X"40", X"3a", X"40", X"37", X"35", X"3c", X"36", X"38", X"3e", X"3b", X"3a", X"3a", X"3d", X"35", X"3a", X"35", X"40", X"38", X"34", X"3a", X"3f", X"3b", X"3c", X"3d", X"3c", X"42", X"3c", X"42", X"44", X"39", X"39", X"35", X"35", X"31", X"30", X"30", X"3a", X"36", X"38", X"3c", X"40", X"3f", X"41", X"37", X"41", X"45", X"3d", X"3c", X"39", X"36", X"31", X"3e", X"3d", X"33", X"41", X"40", X"3c", X"39", X"3d", X"49", X"43", X"42", X"3c", X"3b", X"3c", X"38", X"40", X"32", X"2f", X"2e", X"26", X"1d", X"18", X"20", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"03", X"05", X"06", X"05", X"03", X"01", X"11", X"12", X"18", X"1f", X"29", X"32", X"3e", X"3d", X"39", X"46", X"48", X"3b", X"3f", X"3e", X"40", X"43", X"37", X"3b", X"45", X"42", X"46", X"49", X"42", X"3e", X"44", X"3b", X"42", X"42", X"3e", X"49", X"3f", X"3d", X"47", X"38", X"44", X"3e", X"3b", X"40", X"3a", X"43", X"47", X"40", X"42", X"3c", X"43", X"3f", X"39", X"3f", X"3b", X"3f", X"3f", X"3b", X"39", X"3c", X"3d", X"35", X"3f", X"3b", X"3d", X"40", X"40", X"3c", X"40", X"43", X"39", X"40", X"37", X"43", X"41", X"43", X"35", X"3a", X"35", X"34", X"3a", X"39", X"35", X"27", X"2d", X"2c", X"26", X"12", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"23", X"36", X"48", X"36", X"3b", X"29", X"31", X"35", X"35", X"37", X"37", X"3f", X"3a", X"39", X"3b", X"3b", X"38", X"39", X"3f", X"41", X"38", X"3c", X"3a", X"3c", X"43", X"3e", X"3a", X"35", X"37", X"3b", X"38", X"3e", X"39", X"33", X"38", X"3f", X"3a", X"3f", X"34", X"3a", X"39", X"3e", X"39", X"3d", X"3e", X"34", X"43", X"3f", X"48", X"3b", X"3c", X"3f", X"3c", X"44", X"3c", X"44", X"44", X"3f", X"3b", X"40", X"41", X"46", X"44", X"3b", X"3b", X"3d", X"3e", X"36", X"39", X"31", X"30", X"21", X"1b", X"1b", X"12", X"0f", X"06", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"14", X"0c", X"15", X"23", X"29", X"32", X"39", X"43", X"44", X"42", X"45", X"3f", X"3d", X"39", X"3b", X"39", X"40", X"3b", X"3f", X"35", X"46", X"42", X"3b", X"3b", X"41", X"3b", X"43", X"3c", X"43", X"37", X"3d", X"43", X"4a", X"47", X"41", X"44", X"3d", X"38", X"32", X"40", X"3e", X"3e", X"42", X"37", X"36", X"3b", X"34", X"31", X"37", X"39", X"36", X"37", X"3a", X"35", X"43", X"42", X"3d", X"3d", X"39", X"3b", X"3e", X"3f", X"3a", X"40", X"3a", X"3b", X"3b", X"41", X"42", X"3c", X"40", X"34", X"36", X"33", X"35", X"37", X"2e", X"30", X"25", X"2d", X"11", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"1b", X"33", X"36", X"3d", X"3e", X"39", X"35", X"3f", X"34", X"3a", X"3d", X"3b", X"39", X"37", X"3a", X"36", X"35", X"40", X"38", X"3b", X"37", X"37", X"42", X"39", X"40", X"3f", X"37", X"37", X"41", X"35", X"41", X"39", X"33", X"3b", X"35", X"3a", X"38", X"35", X"3b", X"3f", X"3f", X"3c", X"34", X"33", X"44", X"3b", X"3e", X"3d", X"47", X"44", X"3d", X"4c", X"4b", X"3f", X"4a", X"42", X"40", X"3d", X"3e", X"3d", X"3c", X"44", X"44", X"43", X"42", X"41", X"32", X"2f", X"38", X"2b", X"2b", X"26", X"1c", X"12", X"0c", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"07", X"06", X"0c", X"1d", X"21", X"2a", X"3b", X"32", X"43", X"44", X"44", X"43", X"41", X"3e", X"3c", X"3e", X"3b", X"3e", X"43", X"3e", X"44", X"3c", X"3b", X"3d", X"42", X"3b", X"37", X"3f", X"41", X"42", X"3e", X"3f", X"43", X"43", X"3d", X"3a", X"3c", X"38", X"3e", X"3b", X"41", X"42", X"42", X"40", X"36", X"39", X"33", X"39", X"3c", X"39", X"3f", X"33", X"38", X"36", X"34", X"3a", X"3c", X"3c", X"33", X"34", X"3b", X"3e", X"35", X"47", X"3d", X"39", X"42", X"3a", X"3a", X"37", X"44", X"36", X"3e", X"36", X"2f", X"30", X"32", X"36", X"2c", X"30", X"23", X"12", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"07", X"1b", X"37", X"33", X"38", X"3a", X"2e", X"39", X"3c", X"3c", X"2e", X"32", X"38", X"3c", X"39", X"37", X"3a", X"31", X"3a", X"41", X"3a", X"3a", X"33", X"45", X"3b", X"3d", X"3d", X"3d", X"36", X"3c", X"3d", X"3a", X"3b", X"35", X"38", X"3b", X"40", X"3e", X"2f", X"45", X"3f", X"3e", X"42", X"3d", X"39", X"4d", X"45", X"42", X"4b", X"4f", X"47", X"48", X"52", X"4a", X"49", X"4f", X"43", X"44", X"45", X"41", X"3e", X"3f", X"46", X"3e", X"43", X"40", X"3b", X"3a", X"2f", X"26", X"32", X"30", X"21", X"19", X"11", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"15", X"17", X"20", X"29", X"2d", X"3e", X"48", X"49", X"4a", X"45", X"41", X"43", X"48", X"42", X"3e", X"44", X"43", X"46", X"3e", X"3c", X"43", X"45", X"41", X"4b", X"42", X"41", X"3d", X"42", X"44", X"40", X"3a", X"3f", X"42", X"41", X"37", X"3b", X"3b", X"3e", X"40", X"36", X"3b", X"36", X"31", X"42", X"33", X"3b", X"31", X"38", X"39", X"38", X"37", X"38", X"39", X"38", X"3b", X"37", X"42", X"3d", X"3a", X"3a", X"3e", X"3d", X"35", X"3b", X"40", X"3b", X"44", X"43", X"32", X"41", X"39", X"38", X"3d", X"36", X"39", X"32", X"2b", X"29", X"28", X"17", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"1d", X"32", X"3d", X"39", X"3b", X"2f", X"35", X"38", X"36", X"3c", X"3b", X"35", X"3e", X"42", X"37", X"39", X"3b", X"38", X"3a", X"35", X"39", X"3e", X"45", X"32", X"48", X"36", X"45", X"3a", X"42", X"3d", X"3f", X"3f", X"43", X"3f", X"35", X"3b", X"42", X"3d", X"3e", X"3e", X"40", X"41", X"47", X"48", X"4a", X"4e", X"52", X"5c", X"54", X"5e", X"59", X"57", X"5f", X"5a", X"5c", X"45", X"48", X"55", X"45", X"43", X"3d", X"49", X"49", X"44", X"3d", X"3e", X"36", X"38", X"31", X"26", X"24", X"1e", X"0e", X"0e", X"11", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0b", X"09", X"10", X"1b", X"17", X"27", X"2f", X"37", X"43", X"43", X"4a", X"42", X"42", X"3c", X"3a", X"39", X"44", X"48", X"39", X"48", X"3e", X"3e", X"47", X"41", X"44", X"46", X"40", X"49", X"43", X"37", X"47", X"41", X"3f", X"37", X"3a", X"3f", X"38", X"36", X"36", X"37", X"35", X"3e", X"3a", X"3d", X"3b", X"33", X"3b", X"36", X"32", X"3b", X"34", X"37", X"3f", X"41", X"39", X"39", X"3a", X"3d", X"36", X"43", X"3a", X"38", X"3d", X"42", X"3d", X"42", X"3a", X"40", X"3c", X"43", X"36", X"3d", X"3e", X"3c", X"30", X"28", X"34", X"34", X"2f", X"29", X"10", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"18", X"34", X"33", X"3a", X"40", X"33", X"39", X"39", X"3d", X"34", X"40", X"40", X"44", X"3b", X"38", X"39", X"36", X"3e", X"43", X"40", X"46", X"37", X"41", X"3a", X"44", X"43", X"3f", X"41", X"3b", X"3c", X"3b", X"40", X"3f", X"36", X"41", X"3b", X"40", X"45", X"43", X"43", X"4a", X"59", X"51", X"56", X"5d", X"57", X"5e", X"63", X"60", X"61", X"69", X"73", X"76", X"6d", X"67", X"61", X"5c", X"59", X"53", X"48", X"4b", X"44", X"48", X"44", X"3f", X"3f", X"33", X"36", X"30", X"24", X"1f", X"1b", X"14", X"0c", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"0e", X"16", X"1f", X"24", X"2f", X"39", X"44", X"41", X"49", X"42", X"3d", X"3f", X"41", X"48", X"42", X"3a", X"44", X"34", X"40", X"41", X"3f", X"4c", X"45", X"46", X"41", X"44", X"3f", X"37", X"3c", X"40", X"3c", X"3b", X"3d", X"3c", X"3b", X"35", X"37", X"3c", X"44", X"46", X"42", X"39", X"38", X"34", X"33", X"3d", X"39", X"36", X"3a", X"38", X"3d", X"3d", X"3a", X"30", X"3c", X"40", X"34", X"3e", X"3a", X"3c", X"34", X"37", X"3c", X"40", X"42", X"42", X"47", X"3f", X"46", X"33", X"3b", X"32", X"36", X"32", X"31", X"30", X"30", X"33", X"18", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"15", X"31", X"33", X"39", X"33", X"32", X"3d", X"40", X"35", X"38", X"33", X"41", X"3e", X"3a", X"3e", X"33", X"39", X"38", X"3f", X"42", X"44", X"3f", X"3d", X"3e", X"4d", X"3d", X"44", X"3c", X"45", X"3f", X"41", X"3f", X"4f", X"48", X"46", X"4e", X"40", X"4e", X"51", X"55", X"5e", X"63", X"66", X"66", X"6f", X"72", X"71", X"79", X"7b", X"72", X"7a", X"76", X"7c", X"78", X"78", X"78", X"6f", X"6c", X"60", X"5d", X"5b", X"4e", X"4f", X"43", X"3f", X"3f", X"2e", X"32", X"26", X"26", X"1e", X"1f", X"0c", X"06", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"0f", X"13", X"16", X"24", X"2b", X"37", X"3e", X"46", X"3d", X"42", X"3e", X"49", X"3f", X"36", X"42", X"3b", X"40", X"45", X"42", X"40", X"48", X"3e", X"37", X"44", X"42", X"41", X"40", X"42", X"3d", X"42", X"37", X"40", X"40", X"44", X"38", X"38", X"3b", X"35", X"41", X"37", X"38", X"36", X"3a", X"33", X"39", X"39", X"32", X"33", X"31", X"39", X"39", X"3b", X"3a", X"3c", X"3a", X"3a", X"39", X"3d", X"37", X"41", X"37", X"3c", X"3e", X"3c", X"3f", X"43", X"3d", X"38", X"3d", X"3d", X"3b", X"32", X"35", X"2c", X"38", X"2e", X"3c", X"2a", X"17", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0c", X"34", X"42", X"37", X"33", X"34", X"35", X"37", X"33", X"39", X"3a", X"43", X"44", X"40", X"3f", X"41", X"41", X"44", X"42", X"3d", X"44", X"44", X"40", X"41", X"43", X"44", X"4a", X"47", X"42", X"4b", X"4d", X"4c", X"50", X"53", X"4c", X"4b", X"5b", X"5b", X"65", X"6c", X"6a", X"72", X"75", X"7b", X"80", X"82", X"86", X"87", X"82", X"7a", X"80", X"83", X"84", X"83", X"84", X"78", X"79", X"80", X"79", X"70", X"5d", X"54", X"52", X"4b", X"41", X"3b", X"30", X"31", X"28", X"25", X"2f", X"12", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0a", X"0d", X"15", X"15", X"22", X"2b", X"40", X"3b", X"3f", X"41", X"3b", X"40", X"43", X"3b", X"46", X"40", X"43", X"45", X"42", X"3e", X"33", X"46", X"3d", X"3c", X"3b", X"3c", X"42", X"41", X"35", X"3c", X"3d", X"3a", X"3d", X"37", X"39", X"2f", X"3a", X"45", X"43", X"3f", X"3b", X"31", X"34", X"44", X"3a", X"3b", X"32", X"34", X"3b", X"40", X"3e", X"39", X"33", X"39", X"38", X"3e", X"3b", X"38", X"3d", X"3a", X"34", X"3c", X"3d", X"3a", X"3a", X"3b", X"35", X"37", X"39", X"3d", X"3c", X"39", X"2b", X"2f", X"2d", X"2b", X"27", X"2d", X"1c", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"17", X"2d", X"3c", X"37", X"35", X"34", X"3a", X"3c", X"32", X"3f", X"3a", X"3f", X"47", X"40", X"3e", X"41", X"39", X"37", X"45", X"41", X"43", X"36", X"4c", X"3c", X"49", X"42", X"46", X"44", X"46", X"46", X"52", X"59", X"56", X"5f", X"64", X"69", X"6a", X"6c", X"7c", X"74", X"78", X"8a", X"7f", X"82", X"8c", X"86", X"87", X"85", X"88", X"8d", X"7c", X"85", X"7e", X"83", X"86", X"85", X"7b", X"79", X"7b", X"73", X"6e", X"60", X"58", X"4a", X"44", X"3a", X"35", X"2d", X"25", X"20", X"0d", X"10", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"0b", X"15", X"19", X"25", X"2f", X"39", X"3c", X"46", X"41", X"3b", X"41", X"3a", X"3b", X"3f", X"3b", X"45", X"3c", X"3c", X"40", X"3c", X"3f", X"3f", X"3f", X"46", X"41", X"42", X"35", X"42", X"36", X"39", X"3e", X"3a", X"39", X"39", X"34", X"3e", X"38", X"3e", X"3a", X"30", X"3e", X"3d", X"38", X"35", X"3a", X"2f", X"31", X"31", X"35", X"3a", X"40", X"2f", X"35", X"33", X"37", X"31", X"36", X"38", X"34", X"37", X"35", X"3e", X"39", X"30", X"3b", X"3a", X"38", X"3b", X"35", X"36", X"36", X"32", X"39", X"29", X"28", X"2e", X"2b", X"14", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0e", X"30", X"37", X"32", X"37", X"3b", X"3d", X"37", X"38", X"37", X"47", X"41", X"45", X"3f", X"42", X"41", X"3f", X"41", X"44", X"49", X"44", X"45", X"48", X"45", X"46", X"4b", X"4e", X"4a", X"55", X"56", X"6b", X"67", X"6e", X"74", X"76", X"7d", X"7e", X"84", X"7c", X"82", X"89", X"8c", X"8d", X"85", X"88", X"86", X"8d", X"89", X"83", X"92", X"7e", X"87", X"8c", X"7e", X"84", X"7c", X"82", X"7a", X"7a", X"73", X"6d", X"68", X"64", X"50", X"42", X"36", X"33", X"28", X"28", X"18", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"03", X"07", X"0d", X"14", X"12", X"20", X"28", X"2f", X"36", X"43", X"46", X"4b", X"47", X"44", X"3f", X"40", X"40", X"41", X"3c", X"40", X"44", X"3a", X"3b", X"3d", X"44", X"45", X"3f", X"42", X"3c", X"3e", X"47", X"39", X"45", X"3b", X"3e", X"3a", X"32", X"38", X"39", X"3f", X"3e", X"34", X"37", X"39", X"3a", X"3f", X"34", X"35", X"3a", X"36", X"33", X"3e", X"3b", X"31", X"32", X"35", X"39", X"35", X"39", X"36", X"36", X"34", X"41", X"39", X"38", X"39", X"3d", X"3b", X"3b", X"34", X"34", X"2e", X"3b", X"38", X"35", X"36", X"2e", X"2e", X"27", X"1a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0f", X"33", X"32", X"3a", X"3c", X"3a", X"3b", X"3a", X"31", X"45", X"41", X"51", X"4f", X"45", X"4a", X"4b", X"44", X"4a", X"4e", X"47", X"52", X"4e", X"4d", X"55", X"55", X"59", X"5d", X"64", X"6d", X"71", X"77", X"7e", X"80", X"83", X"8b", X"8c", X"91", X"8c", X"83", X"90", X"89", X"8e", X"93", X"8f", X"8b", X"89", X"8f", X"8b", X"90", X"89", X"8c", X"88", X"7e", X"85", X"86", X"7c", X"84", X"7c", X"77", X"78", X"74", X"71", X"63", X"55", X"4d", X"39", X"33", X"28", X"20", X"16", X"14", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"09", X"12", X"14", X"20", X"26", X"2e", X"37", X"43", X"39", X"44", X"43", X"44", X"3a", X"3d", X"3d", X"39", X"38", X"36", X"39", X"43", X"3c", X"41", X"3e", X"3c", X"3f", X"3d", X"3f", X"3c", X"3e", X"3c", X"3d", X"3e", X"44", X"3c", X"31", X"2e", X"39", X"3c", X"33", X"36", X"3a", X"35", X"39", X"34", X"3e", X"38", X"3b", X"39", X"36", X"38", X"33", X"38", X"3b", X"37", X"39", X"31", X"33", X"35", X"34", X"3a", X"36", X"35", X"33", X"3b", X"3f", X"3a", X"34", X"3e", X"34", X"38", X"34", X"33", X"2b", X"2e", X"29", X"2a", X"22", X"1b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"30", X"34", X"3f", X"44", X"3b", X"43", X"43", X"44", X"49", X"4c", X"4d", X"4c", X"4a", X"52", X"49", X"4b", X"56", X"56", X"56", X"54", X"57", X"65", X"62", X"6e", X"73", X"71", X"7d", X"7c", X"81", X"8a", X"8d", X"86", X"8b", X"8f", X"8f", X"94", X"95", X"93", X"8d", X"8e", X"92", X"90", X"8a", X"8a", X"8e", X"8a", X"8e", X"8e", X"87", X"8c", X"7f", X"81", X"7f", X"84", X"7d", X"85", X"74", X"7a", X"77", X"6f", X"6a", X"60", X"5a", X"4d", X"3b", X"2f", X"26", X"20", X"14", X"09", X"0a", X"09", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"06", X"06", X"13", X"11", X"1a", X"20", X"2e", X"36", X"39", X"3a", X"42", X"43", X"45", X"33", X"41", X"38", X"4e", X"37", X"38", X"42", X"4a", X"3d", X"39", X"38", X"3e", X"3a", X"41", X"41", X"39", X"3c", X"3a", X"3e", X"3e", X"45", X"2b", X"39", X"34", X"3c", X"3f", X"33", X"33", X"34", X"41", X"33", X"33", X"35", X"3a", X"40", X"38", X"34", X"3c", X"37", X"3d", X"30", X"3b", X"3b", X"32", X"33", X"3a", X"2c", X"3a", X"32", X"36", X"3c", X"36", X"38", X"3a", X"3a", X"33", X"39", X"37", X"35", X"34", X"2d", X"2d", X"28", X"24", X"2c", X"19", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"10", X"2d", X"38", X"40", X"40", X"32", X"4a", X"42", X"44", X"51", X"58", X"57", X"59", X"4f", X"53", X"5b", X"5e", X"64", X"63", X"6f", X"77", X"78", X"75", X"78", X"84", X"83", X"8f", X"93", X"92", X"96", X"94", X"97", X"91", X"9f", X"8f", X"95", X"99", X"94", X"96", X"8f", X"8f", X"90", X"8c", X"91", X"8f", X"7e", X"80", X"84", X"7f", X"8a", X"7d", X"87", X"84", X"7f", X"84", X"85", X"81", X"76", X"70", X"6b", X"6d", X"61", X"5e", X"55", X"42", X"38", X"2b", X"21", X"1a", X"0a", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"0e", X"08", X"0f", X"18", X"28", X"2e", X"39", X"40", X"44", X"45", X"44", X"3f", X"4a", X"3d", X"3d", X"44", X"42", X"38", X"3c", X"3f", X"43", X"3f", X"41", X"38", X"47", X"40", X"45", X"3b", X"34", X"3f", X"3b", X"3a", X"3d", X"3a", X"3a", X"3e", X"40", X"3d", X"38", X"30", X"39", X"2f", X"38", X"3d", X"38", X"3b", X"34", X"39", X"39", X"33", X"39", X"35", X"38", X"37", X"37", X"39", X"3c", X"32", X"3e", X"37", X"33", X"36", X"30", X"3e", X"36", X"3a", X"30", X"36", X"32", X"33", X"30", X"36", X"2e", X"38", X"2d", X"25", X"1e", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"10", X"3d", X"4d", X"42", X"44", X"44", X"50", X"53", X"53", X"5b", X"60", X"65", X"6f", X"6a", X"6b", X"72", X"78", X"7e", X"7d", X"7e", X"8c", X"8a", X"95", X"8b", X"93", X"93", X"91", X"93", X"9b", X"99", X"96", X"98", X"97", X"96", X"95", X"92", X"95", X"90", X"90", X"8e", X"92", X"8b", X"8b", X"8d", X"8f", X"87", X"87", X"8d", X"83", X"82", X"78", X"84", X"80", X"79", X"79", X"79", X"7e", X"7e", X"76", X"76", X"70", X"62", X"5a", X"4e", X"3c", X"31", X"2f", X"22", X"1a", X"0b", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"08", X"06", X"08", X"0a", X"0e", X"1e", X"1e", X"2b", X"3a", X"3b", X"3f", X"42", X"3a", X"39", X"46", X"3e", X"44", X"3d", X"44", X"3e", X"40", X"43", X"3c", X"43", X"3e", X"38", X"3d", X"3a", X"42", X"3e", X"3d", X"3f", X"38", X"36", X"44", X"40", X"3d", X"3f", X"38", X"3f", X"3d", X"39", X"3d", X"3b", X"2f", X"35", X"36", X"3e", X"38", X"39", X"3c", X"2f", X"37", X"34", X"33", X"3c", X"35", X"35", X"37", X"2b", X"37", X"36", X"3b", X"2b", X"36", X"3a", X"37", X"39", X"33", X"31", X"35", X"2c", X"34", X"33", X"2e", X"2b", X"2b", X"2c", X"21", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0f", X"3c", X"46", X"4c", X"55", X"57", X"64", X"68", X"68", X"6f", X"7c", X"75", X"84", X"85", X"8a", X"89", X"8c", X"96", X"92", X"91", X"98", X"99", X"96", X"90", X"97", X"9a", X"9d", X"9b", X"98", X"96", X"99", X"98", X"94", X"92", X"93", X"94", X"94", X"90", X"8e", X"8b", X"88", X"89", X"89", X"87", X"88", X"82", X"81", X"89", X"84", X"83", X"7e", X"82", X"7b", X"73", X"7a", X"77", X"75", X"7c", X"6f", X"6d", X"64", X"5e", X"57", X"40", X"3e", X"33", X"22", X"1c", X"0e", X"0d", X"06", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0e", X"12", X"21", X"20", X"34", X"30", X"3e", X"3a", X"38", X"3b", X"3c", X"3c", X"3e", X"44", X"3a", X"40", X"3b", X"34", X"46", X"3b", X"3f", X"40", X"43", X"39", X"40", X"3b", X"40", X"3e", X"3d", X"35", X"44", X"35", X"37", X"37", X"3c", X"37", X"36", X"40", X"3b", X"42", X"31", X"34", X"3c", X"38", X"39", X"33", X"30", X"2f", X"31", X"36", X"33", X"3b", X"32", X"36", X"32", X"2f", X"35", X"2f", X"2f", X"32", X"32", X"39", X"3a", X"35", X"2d", X"31", X"36", X"33", X"34", X"2f", X"2f", X"2d", X"2b", X"33", X"16", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"0f", X"42", X"61", X"5f", X"7a", X"6b", X"78", X"79", X"7a", X"84", X"84", X"8a", X"90", X"92", X"8e", X"94", X"8f", X"93", X"94", X"92", X"a1", X"9b", X"9b", X"9a", X"95", X"9f", X"94", X"96", X"96", X"98", X"95", X"96", X"8e", X"8f", X"8d", X"8d", X"99", X"90", X"89", X"8e", X"90", X"82", X"84", X"89", X"89", X"81", X"81", X"82", X"7c", X"7e", X"7a", X"82", X"7c", X"75", X"76", X"72", X"75", X"71", X"70", X"72", X"66", X"56", X"4f", X"4d", X"37", X"2f", X"22", X"16", X"0e", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"15", X"15", X"25", X"1b", X"29", X"2f", X"38", X"3f", X"41", X"38", X"43", X"47", X"42", X"49", X"42", X"44", X"45", X"44", X"42", X"42", X"3c", X"3b", X"3e", X"43", X"41", X"3c", X"46", X"45", X"3e", X"3f", X"3a", X"3e", X"3f", X"42", X"37", X"3e", X"3e", X"39", X"40", X"34", X"36", X"3a", X"3c", X"3d", X"32", X"34", X"2e", X"37", X"34", X"31", X"37", X"3b", X"37", X"39", X"35", X"32", X"3c", X"39", X"33", X"33", X"3a", X"36", X"35", X"34", X"39", X"3d", X"39", X"2e", X"30", X"32", X"33", X"33", X"2f", X"2d", X"25", X"07", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"1a", X"5a", X"79", X"82", X"84", X"83", X"89", X"8d", X"8f", X"8e", X"8f", X"97", X"95", X"9b", X"96", X"93", X"9d", X"92", X"95", X"96", X"98", X"95", X"97", X"96", X"9e", X"96", X"96", X"92", X"90", X"99", X"95", X"8a", X"91", X"8e", X"88", X"8d", X"8f", X"8a", X"81", X"86", X"8a", X"91", X"88", X"85", X"82", X"80", X"7b", X"85", X"88", X"7e", X"7a", X"72", X"78", X"77", X"72", X"70", X"74", X"6f", X"67", X"68", X"59", X"4c", X"4e", X"40", X"2a", X"24", X"23", X"0b", X"10", X"0a", X"0b", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"06", X"06", X"0a", X"0f", X"14", X"13", X"21", X"2b", X"2c", X"33", X"3e", X"3a", X"3a", X"44", X"3e", X"40", X"3d", X"46", X"46", X"3e", X"44", X"44", X"41", X"3c", X"48", X"3b", X"3c", X"44", X"45", X"45", X"44", X"42", X"43", X"42", X"3d", X"3a", X"42", X"42", X"4a", X"42", X"3d", X"3a", X"3b", X"3c", X"3f", X"39", X"3b", X"35", X"3b", X"39", X"37", X"38", X"35", X"35", X"3b", X"30", X"36", X"3e", X"36", X"35", X"37", X"36", X"33", X"34", X"39", X"42", X"35", X"38", X"39", X"33", X"39", X"2f", X"2d", X"2e", X"2f", X"29", X"27", X"2a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"10", X"59", X"84", X"8b", X"90", X"8e", X"8d", X"96", X"8b", X"90", X"92", X"8d", X"a0", X"99", X"93", X"93", X"9c", X"97", X"97", X"95", X"95", X"97", X"96", X"92", X"91", X"93", X"97", X"8f", X"8a", X"94", X"91", X"8e", X"90", X"88", X"8c", X"89", X"90", X"87", X"88", X"7e", X"87", X"88", X"7c", X"7e", X"84", X"7c", X"74", X"7a", X"7b", X"75", X"73", X"7e", X"7a", X"75", X"6f", X"6d", X"71", X"67", X"63", X"68", X"57", X"43", X"38", X"3b", X"2e", X"25", X"13", X"10", X"10", X"03", X"06", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0b", X"03", X"07", X"0b", X"0b", X"1c", X"21", X"2b", X"31", X"30", X"34", X"43", X"3f", X"4b", X"46", X"41", X"3f", X"45", X"49", X"42", X"46", X"46", X"45", X"42", X"3e", X"36", X"48", X"47", X"45", X"50", X"4d", X"43", X"43", X"45", X"46", X"45", X"4b", X"4c", X"3d", X"48", X"49", X"43", X"32", X"35", X"35", X"33", X"3a", X"3b", X"36", X"37", X"36", X"2b", X"38", X"3c", X"37", X"37", X"35", X"3a", X"36", X"36", X"3d", X"30", X"39", X"30", X"35", X"35", X"36", X"33", X"35", X"30", X"35", X"32", X"31", X"32", X"2f", X"2b", X"25", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"14", X"63", X"86", X"8f", X"8c", X"8d", X"8e", X"8f", X"90", X"93", X"8f", X"98", X"8e", X"97", X"9a", X"95", X"94", X"94", X"91", X"94", X"8e", X"97", X"8f", X"90", X"97", X"95", X"96", X"8e", X"8f", X"8d", X"80", X"8c", X"88", X"7f", X"82", X"84", X"7f", X"7a", X"7f", X"7d", X"7d", X"7d", X"7b", X"7a", X"7a", X"7b", X"7c", X"7b", X"6d", X"78", X"79", X"77", X"6d", X"71", X"74", X"65", X"74", X"6c", X"64", X"5e", X"5a", X"49", X"3a", X"32", X"23", X"22", X"13", X"0f", X"08", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"01", X"06", X"05", X"07", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"0d", X"05", X"0f", X"14", X"14", X"22", X"30", X"23", X"33", X"33", X"3b", X"44", X"47", X"43", X"4a", X"48", X"4b", X"49", X"45", X"45", X"43", X"44", X"44", X"44", X"3b", X"40", X"45", X"40", X"49", X"44", X"46", X"44", X"46", X"42", X"50", X"39", X"24", X"36", X"56", X"51", X"43", X"38", X"31", X"38", X"38", X"3c", X"37", X"34", X"2e", X"30", X"31", X"35", X"3d", X"35", X"3d", X"35", X"31", X"31", X"36", X"31", X"3b", X"33", X"33", X"36", X"3a", X"3f", X"2f", X"32", X"3c", X"32", X"34", X"32", X"2c", X"34", X"26", X"2b", X"09", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"10", X"60", X"86", X"95", X"98", X"92", X"8a", X"92", X"8d", X"8d", X"8f", X"8d", X"95", X"8e", X"94", X"98", X"95", X"88", X"95", X"96", X"8b", X"8d", X"91", X"8d", X"8e", X"87", X"8c", X"91", X"85", X"85", X"86", X"7e", X"7e", X"86", X"7a", X"86", X"7e", X"77", X"6e", X"71", X"7c", X"82", X"73", X"73", X"7e", X"74", X"75", X"79", X"77", X"79", X"76", X"74", X"6f", X"6c", X"68", X"68", X"70", X"60", X"5f", X"5a", X"52", X"48", X"34", X"2b", X"1e", X"14", X"0d", X"11", X"07", X"06", X"02", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"07", X"05", X"0b", X"0d", X"12", X"1d", X"24", X"2d", X"32", X"35", X"39", X"3f", X"42", X"49", X"51", X"45", X"53", X"4c", X"41", X"45", X"48", X"3d", X"47", X"40", X"45", X"45", X"41", X"3b", X"4c", X"42", X"40", X"4b", X"41", X"48", X"46", X"46", X"4c", X"4d", X"52", X"48", X"3f", X"3d", X"39", X"38", X"3d", X"35", X"35", X"38", X"33", X"33", X"36", X"30", X"31", X"30", X"31", X"39", X"3d", X"3c", X"3a", X"41", X"37", X"3a", X"39", X"38", X"2f", X"37", X"36", X"39", X"36", X"36", X"37", X"36", X"2e", X"2d", X"30", X"24", X"0f", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0e", X"54", X"89", X"8d", X"93", X"88", X"8e", X"8f", X"81", X"8f", X"8d", X"89", X"93", X"8d", X"95", X"92", X"8a", X"8d", X"87", X"86", X"82", X"87", X"8c", X"8e", X"87", X"89", X"8b", X"85", X"7e", X"7e", X"85", X"88", X"82", X"77", X"7c", X"80", X"7c", X"79", X"79", X"7e", X"7f", X"7a", X"78", X"79", X"70", X"6b", X"78", X"78", X"75", X"6d", X"70", X"66", X"75", X"65", X"64", X"68", X"6e", X"58", X"5b", X"56", X"48", X"42", X"32", X"2d", X"1f", X"11", X"0e", X"06", X"10", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0a", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"06", X"0b", X"10", X"13", X"1e", X"22", X"2d", X"3a", X"31", X"3b", X"41", X"43", X"45", X"43", X"51", X"59", X"4b", X"47", X"48", X"47", X"45", X"3c", X"41", X"44", X"3e", X"44", X"47", X"4b", X"40", X"47", X"44", X"40", X"50", X"49", X"43", X"3e", X"3e", X"47", X"37", X"38", X"38", X"2f", X"3d", X"3c", X"39", X"39", X"31", X"37", X"34", X"37", X"3c", X"36", X"34", X"33", X"39", X"38", X"31", X"3e", X"31", X"34", X"36", X"2f", X"38", X"3d", X"2d", X"3a", X"39", X"35", X"37", X"2e", X"28", X"32", X"27", X"25", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"55", X"7d", X"8f", X"97", X"88", X"8a", X"84", X"8a", X"85", X"8b", X"86", X"8e", X"84", X"8d", X"87", X"86", X"88", X"88", X"89", X"85", X"83", X"8a", X"7b", X"84", X"85", X"83", X"82", X"7e", X"76", X"7c", X"78", X"7c", X"7a", X"75", X"7e", X"73", X"76", X"72", X"73", X"70", X"77", X"79", X"6e", X"73", X"64", X"70", X"76", X"74", X"6d", X"6e", X"6a", X"6b", X"62", X"5f", X"5e", X"65", X"55", X"56", X"47", X"3f", X"30", X"31", X"1a", X"1f", X"09", X"0e", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"0a", X"0c", X"0a", X"14", X"26", X"20", X"30", X"2e", X"35", X"34", X"3a", X"43", X"45", X"49", X"49", X"59", X"57", X"52", X"45", X"43", X"41", X"48", X"38", X"3e", X"38", X"3d", X"43", X"4a", X"3e", X"3a", X"42", X"3b", X"43", X"43", X"42", X"3a", X"3c", X"41", X"38", X"33", X"34", X"37", X"31", X"39", X"41", X"3f", X"37", X"33", X"2b", X"34", X"38", X"3a", X"39", X"3b", X"35", X"3b", X"32", X"39", X"39", X"34", X"37", X"40", X"3a", X"36", X"3c", X"33", X"35", X"31", X"29", X"37", X"35", X"2d", X"3e", X"29", X"10", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"4b", X"85", X"8b", X"8d", X"84", X"89", X"86", X"8b", X"85", X"85", X"82", X"81", X"8b", X"89", X"85", X"83", X"86", X"88", X"86", X"7e", X"7d", X"7d", X"79", X"7c", X"7d", X"7b", X"76", X"7c", X"7b", X"7e", X"7b", X"78", X"76", X"78", X"77", X"74", X"6e", X"70", X"72", X"70", X"69", X"74", X"75", X"72", X"6b", X"6f", X"6a", X"66", X"6d", X"70", X"65", X"65", X"6b", X"66", X"65", X"5a", X"57", X"53", X"48", X"3d", X"2a", X"1e", X"1f", X"1b", X"0f", X"0a", X"09", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"08", X"0b", X"11", X"10", X"1f", X"20", X"28", X"2a", X"32", X"3c", X"3b", X"3d", X"42", X"4f", X"4e", X"53", X"54", X"55", X"4c", X"4c", X"3f", X"44", X"42", X"41", X"41", X"44", X"44", X"37", X"41", X"44", X"3f", X"42", X"42", X"3d", X"40", X"3d", X"48", X"3e", X"34", X"3e", X"38", X"42", X"45", X"36", X"3b", X"38", X"35", X"33", X"3e", X"33", X"2d", X"2f", X"3a", X"3e", X"3f", X"3d", X"3b", X"3a", X"3a", X"35", X"39", X"3c", X"2f", X"34", X"3b", X"39", X"37", X"3b", X"31", X"38", X"38", X"35", X"36", X"38", X"15", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"04", X"06", X"0d", X"4a", X"7d", X"7f", X"8b", X"85", X"88", X"7d", X"8b", X"7e", X"82", X"82", X"91", X"81", X"7e", X"83", X"84", X"7a", X"7e", X"7c", X"7d", X"7f", X"83", X"80", X"82", X"74", X"7b", X"7e", X"79", X"7b", X"75", X"74", X"73", X"73", X"76", X"70", X"70", X"70", X"67", X"70", X"6d", X"6d", X"75", X"6d", X"6a", X"6b", X"6f", X"66", X"6a", X"6d", X"66", X"71", X"64", X"5d", X"61", X"59", X"57", X"4a", X"4a", X"40", X"35", X"28", X"23", X"1e", X"13", X"13", X"0f", X"10", X"08", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"0e", X"0f", X"0b", X"10", X"1e", X"23", X"2d", X"34", X"36", X"32", X"3d", X"44", X"43", X"49", X"50", X"4c", X"4d", X"51", X"44", X"4c", X"44", X"42", X"44", X"43", X"40", X"40", X"45", X"45", X"4a", X"39", X"33", X"3a", X"39", X"40", X"3e", X"3a", X"3a", X"35", X"36", X"37", X"38", X"44", X"36", X"2f", X"35", X"35", X"3d", X"3b", X"3a", X"34", X"39", X"3c", X"35", X"30", X"31", X"33", X"30", X"34", X"36", X"3e", X"44", X"3b", X"3c", X"32", X"3b", X"3b", X"3a", X"2f", X"40", X"41", X"41", X"4a", X"40", X"1b", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"40", X"73", X"7a", X"84", X"82", X"87", X"7c", X"7b", X"7e", X"79", X"7c", X"80", X"7d", X"7d", X"79", X"83", X"78", X"7a", X"7e", X"80", X"7c", X"80", X"79", X"75", X"6e", X"78", X"6d", X"78", X"7e", X"77", X"7a", X"75", X"6b", X"77", X"70", X"6a", X"72", X"6f", X"73", X"71", X"71", X"6e", X"69", X"71", X"6e", X"69", X"70", X"67", X"61", X"61", X"62", X"65", X"54", X"55", X"4e", X"54", X"48", X"3f", X"38", X"2a", X"20", X"1f", X"13", X"14", X"0a", X"07", X"06", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"06", X"0c", X"15", X"11", X"22", X"25", X"29", X"30", X"38", X"37", X"3c", X"41", X"3c", X"47", X"48", X"4a", X"5b", X"4a", X"40", X"47", X"41", X"41", X"49", X"43", X"4e", X"3d", X"39", X"3b", X"3a", X"37", X"38", X"37", X"41", X"35", X"39", X"3d", X"3d", X"32", X"37", X"3f", X"3b", X"31", X"3e", X"33", X"30", X"39", X"2f", X"3c", X"36", X"31", X"39", X"3d", X"3f", X"35", X"37", X"37", X"3e", X"34", X"33", X"39", X"3a", X"3c", X"33", X"3f", X"3d", X"44", X"44", X"41", X"41", X"41", X"4e", X"4b", X"29", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"30", X"6e", X"7d", X"89", X"79", X"85", X"84", X"80", X"77", X"7a", X"7d", X"7b", X"84", X"7b", X"7e", X"79", X"77", X"83", X"77", X"7b", X"77", X"75", X"76", X"75", X"74", X"73", X"77", X"6f", X"77", X"70", X"69", X"6d", X"6b", X"73", X"76", X"71", X"62", X"6c", X"78", X"68", X"6b", X"6a", X"5e", X"6c", X"68", X"5e", X"6b", X"5d", X"66", X"60", X"61", X"5e", X"52", X"5a", X"52", X"4e", X"44", X"3d", X"39", X"26", X"1e", X"19", X"0e", X"0c", X"0c", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"01", X"06", X"05", X"0a", X"10", X"0e", X"1b", X"1e", X"24", X"2a", X"30", X"2f", X"35", X"3c", X"39", X"3d", X"48", X"44", X"48", X"48", X"44", X"4b", X"4a", X"42", X"4d", X"4e", X"45", X"44", X"3f", X"40", X"3c", X"40", X"35", X"39", X"35", X"3a", X"35", X"36", X"38", X"39", X"37", X"35", X"3c", X"3a", X"34", X"39", X"3d", X"37", X"36", X"36", X"41", X"38", X"3d", X"37", X"3c", X"35", X"45", X"3a", X"38", X"34", X"3b", X"3b", X"3f", X"41", X"3f", X"3e", X"43", X"3e", X"40", X"49", X"55", X"60", X"5f", X"69", X"63", X"2b", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"3a", X"71", X"7a", X"81", X"77", X"75", X"76", X"75", X"7b", X"7c", X"7e", X"75", X"7a", X"80", X"79", X"7b", X"73", X"81", X"7c", X"84", X"70", X"6f", X"79", X"75", X"70", X"76", X"74", X"78", X"74", X"6b", X"72", X"70", X"6e", X"72", X"6b", X"74", X"68", X"72", X"69", X"6e", X"72", X"6b", X"6c", X"65", X"6d", X"64", X"61", X"62", X"65", X"5e", X"62", X"54", X"52", X"56", X"43", X"4c", X"3f", X"33", X"39", X"25", X"12", X"13", X"0f", X"19", X"12", X"0d", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"09", X"05", X"03", X"14", X"0f", X"17", X"1f", X"21", X"25", X"2d", X"37", X"34", X"36", X"41", X"44", X"43", X"3e", X"47", X"44", X"42", X"44", X"42", X"3d", X"46", X"42", X"47", X"41", X"3e", X"45", X"3d", X"3b", X"3b", X"34", X"39", X"40", X"3d", X"3f", X"3e", X"42", X"35", X"33", X"35", X"36", X"33", X"3f", X"35", X"38", X"32", X"35", X"35", X"33", X"39", X"3b", X"3b", X"35", X"3d", X"33", X"3d", X"38", X"38", X"3b", X"3e", X"3f", X"3e", X"44", X"4b", X"4e", X"52", X"5b", X"60", X"6a", X"74", X"80", X"74", X"3d", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"06", X"2e", X"65", X"77", X"83", X"79", X"75", X"77", X"75", X"7c", X"71", X"76", X"79", X"75", X"7d", X"79", X"7e", X"72", X"7d", X"79", X"7c", X"74", X"6c", X"76", X"72", X"71", X"6e", X"6c", X"76", X"68", X"75", X"6e", X"75", X"6e", X"71", X"70", X"6b", X"6e", X"6b", X"60", X"67", X"68", X"69", X"66", X"66", X"5d", X"58", X"65", X"61", X"60", X"60", X"59", X"52", X"51", X"50", X"49", X"40", X"39", X"29", X"1e", X"23", X"19", X"22", X"0d", X"11", X"0b", X"06", X"06", X"06", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"0f", X"0c", X"0a", X"12", X"13", X"22", X"21", X"29", X"2c", X"2f", X"3a", X"41", X"36", X"39", X"40", X"4a", X"3d", X"49", X"45", X"4b", X"3f", X"47", X"43", X"43", X"44", X"3c", X"3d", X"41", X"3c", X"38", X"37", X"38", X"38", X"39", X"38", X"3b", X"35", X"34", X"37", X"37", X"34", X"32", X"39", X"37", X"31", X"31", X"34", X"39", X"38", X"32", X"37", X"36", X"34", X"37", X"41", X"37", X"3a", X"3a", X"41", X"44", X"43", X"4c", X"41", X"51", X"54", X"68", X"73", X"75", X"75", X"7f", X"78", X"74", X"49", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0c", X"25", X"63", X"75", X"79", X"76", X"70", X"70", X"73", X"6f", X"79", X"6e", X"7f", X"6a", X"74", X"76", X"75", X"73", X"72", X"73", X"70", X"6e", X"74", X"6f", X"6b", X"6f", X"6f", X"6b", X"63", X"66", X"68", X"73", X"69", X"68", X"68", X"68", X"62", X"6c", X"62", X"63", X"68", X"62", X"60", X"5f", X"5e", X"5f", X"5c", X"5e", X"5c", X"5b", X"54", X"4b", X"4b", X"45", X"4e", X"42", X"3c", X"3b", X"2e", X"26", X"22", X"12", X"0e", X"06", X"06", X"07", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"0d", X"05", X"05", X"09", X"09", X"0e", X"1b", X"1f", X"25", X"2d", X"38", X"36", X"31", X"32", X"42", X"43", X"43", X"45", X"3e", X"45", X"4f", X"46", X"40", X"49", X"40", X"3e", X"42", X"3d", X"43", X"3b", X"3c", X"38", X"43", X"3c", X"3a", X"33", X"33", X"39", X"38", X"36", X"39", X"3a", X"32", X"38", X"34", X"32", X"3a", X"2c", X"3a", X"37", X"31", X"32", X"39", X"3c", X"3d", X"3e", X"38", X"33", X"3e", X"39", X"46", X"47", X"50", X"59", X"63", X"70", X"7d", X"7e", X"85", X"81", X"84", X"83", X"76", X"48", X"0a", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"20", X"5f", X"75", X"7e", X"70", X"6c", X"70", X"6d", X"71", X"74", X"71", X"72", X"6d", X"73", X"6d", X"75", X"74", X"74", X"79", X"6b", X"6d", X"72", X"72", X"75", X"6f", X"7c", X"65", X"68", X"6a", X"6d", X"72", X"6f", X"67", X"62", X"69", X"61", X"64", X"69", X"69", X"69", X"68", X"67", X"57", X"63", X"5d", X"5f", X"64", X"5c", X"59", X"5c", X"55", X"56", X"4a", X"43", X"3c", X"3e", X"35", X"20", X"20", X"1a", X"12", X"16", X"0a", X"0b", X"0c", X"09", X"06", X"07", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"09", X"0e", X"11", X"06", X"0b", X"14", X"1a", X"1b", X"21", X"29", X"34", X"2f", X"3a", X"3f", X"3f", X"42", X"42", X"45", X"44", X"43", X"4a", X"41", X"49", X"47", X"3f", X"41", X"3e", X"3a", X"42", X"3f", X"45", X"43", X"3e", X"39", X"3a", X"3b", X"33", X"35", X"32", X"36", X"3a", X"38", X"30", X"37", X"3b", X"36", X"3e", X"2d", X"38", X"35", X"33", X"34", X"38", X"2e", X"40", X"36", X"3f", X"39", X"41", X"45", X"48", X"59", X"5a", X"64", X"68", X"7a", X"7d", X"83", X"86", X"85", X"88", X"81", X"7d", X"53", X"10", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"23", X"5c", X"70", X"75", X"70", X"6b", X"72", X"71", X"6a", X"6c", X"66", X"70", X"6a", X"70", X"75", X"6e", X"70", X"6d", X"73", X"77", X"6c", X"6d", X"73", X"6e", X"6b", X"74", X"6b", X"6d", X"68", X"70", X"66", X"6e", X"61", X"6c", X"6a", X"5f", X"62", X"60", X"60", X"66", X"61", X"64", X"66", X"5f", X"5d", X"5a", X"5f", X"5b", X"4d", X"52", X"50", X"4d", X"46", X"40", X"35", X"2b", X"2e", X"26", X"21", X"17", X"0f", X"1a", X"0f", X"05", X"0a", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"09", X"06", X"07", X"09", X"10", X"17", X"20", X"27", X"35", X"33", X"34", X"39", X"3c", X"3c", X"3b", X"3c", X"3b", X"4b", X"4a", X"46", X"48", X"47", X"3d", X"3a", X"3c", X"34", X"3b", X"36", X"3e", X"36", X"39", X"38", X"35", X"35", X"36", X"33", X"3b", X"36", X"3d", X"35", X"31", X"35", X"37", X"32", X"35", X"32", X"36", X"34", X"2f", X"36", X"31", X"37", X"36", X"35", X"37", X"3f", X"43", X"51", X"51", X"62", X"70", X"7f", X"7a", X"85", X"7e", X"8d", X"7e", X"80", X"84", X"83", X"72", X"4e", X"10", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"23", X"52", X"61", X"74", X"64", X"6b", X"68", X"6e", X"6d", X"66", X"6d", X"6d", X"73", X"71", X"6c", X"73", X"73", X"6f", X"6d", X"6c", X"68", X"6b", X"6a", X"67", X"6d", X"6e", X"60", X"70", X"68", X"66", X"64", X"66", X"65", X"64", X"64", X"64", X"5e", X"5f", X"66", X"5d", X"60", X"5f", X"61", X"5f", X"5b", X"58", X"4f", X"63", X"50", X"4a", X"4c", X"4a", X"3b", X"39", X"33", X"31", X"2e", X"23", X"1a", X"10", X"0e", X"09", X"0c", X"06", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"06", X"06", X"05", X"08", X"0e", X"18", X"15", X"26", X"23", X"2d", X"31", X"33", X"3a", X"3b", X"37", X"3d", X"3d", X"47", X"44", X"49", X"45", X"46", X"3f", X"40", X"3c", X"41", X"3e", X"3c", X"3d", X"3f", X"34", X"3c", X"3d", X"3c", X"3e", X"2e", X"37", X"39", X"3a", X"3a", X"37", X"3e", X"38", X"2f", X"34", X"3e", X"36", X"3f", X"32", X"39", X"3c", X"3d", X"38", X"38", X"34", X"40", X"54", X"5a", X"69", X"79", X"7d", X"82", X"87", X"83", X"80", X"89", X"86", X"86", X"88", X"83", X"7a", X"50", X"16", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"1e", X"57", X"6d", X"6e", X"67", X"64", X"76", X"6b", X"6d", X"6f", X"71", X"6d", X"6f", X"68", X"6c", X"73", X"6b", X"69", X"6c", X"6b", X"66", X"6a", X"62", X"65", X"62", X"64", X"6c", X"5e", X"68", X"63", X"6e", X"69", X"5d", X"61", X"5e", X"66", X"59", X"5d", X"61", X"5d", X"61", X"5c", X"61", X"5f", X"62", X"5d", X"54", X"52", X"50", X"4a", X"44", X"3f", X"3a", X"41", X"32", X"2e", X"25", X"19", X"1d", X"11", X"0b", X"10", X"08", X"05", X"09", X"09", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"09", X"06", X"0b", X"09", X"0d", X"11", X"19", X"22", X"30", X"25", X"2f", X"32", X"37", X"3e", X"43", X"42", X"3f", X"42", X"40", X"3e", X"4a", X"43", X"41", X"47", X"41", X"47", X"3e", X"3c", X"36", X"3a", X"44", X"38", X"3b", X"43", X"35", X"3c", X"36", X"33", X"33", X"37", X"41", X"35", X"3d", X"32", X"32", X"3a", X"34", X"37", X"3d", X"35", X"3b", X"3c", X"44", X"40", X"43", X"48", X"4d", X"6a", X"70", X"7c", X"89", X"86", X"8d", X"8a", X"8a", X"87", X"83", X"80", X"86", X"7d", X"7d", X"51", X"15", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"1c", X"59", X"6a", X"69", X"65", X"6b", X"64", X"6b", X"6b", X"6e", X"6a", X"65", X"5e", X"6e", X"66", X"6d", X"6b", X"6f", X"6d", X"6e", X"66", X"69", X"65", X"69", X"61", X"69", X"65", X"63", X"68", X"64", X"66", X"60", X"64", X"67", X"5c", X"62", X"60", X"61", X"68", X"5c", X"58", X"60", X"5a", X"58", X"55", X"51", X"54", X"51", X"4b", X"44", X"3e", X"3e", X"2f", X"30", X"30", X"26", X"1e", X"18", X"18", X"11", X"11", X"13", X"09", X"05", X"03", X"0e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"00", X"09", X"05", X"0b", X"10", X"0b", X"13", X"16", X"18", X"2a", X"34", X"2f", X"32", X"33", X"38", X"49", X"3a", X"47", X"42", X"47", X"3d", X"41", X"47", X"41", X"47", X"46", X"3d", X"39", X"39", X"38", X"36", X"3c", X"32", X"39", X"38", X"33", X"34", X"34", X"34", X"38", X"3f", X"3f", X"37", X"35", X"2f", X"31", X"35", X"32", X"2f", X"37", X"37", X"38", X"44", X"3b", X"43", X"4d", X"5f", X"67", X"86", X"89", X"87", X"82", X"86", X"89", X"8a", X"88", X"84", X"89", X"81", X"79", X"7a", X"60", X"1b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"14", X"4d", X"6b", X"6f", X"70", X"6c", X"65", X"6b", X"6a", X"67", X"60", X"6a", X"6a", X"60", X"6a", X"65", X"6a", X"6b", X"63", X"64", X"5e", X"68", X"6a", X"63", X"68", X"68", X"62", X"5d", X"61", X"63", X"63", X"66", X"5a", X"55", X"61", X"60", X"5f", X"59", X"61", X"60", X"61", X"51", X"5b", X"56", X"4e", X"53", X"52", X"49", X"46", X"49", X"37", X"36", X"31", X"2b", X"20", X"27", X"1a", X"21", X"17", X"0f", X"12", X"0d", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"01", X"06", X"05", X"03", X"00", X"07", X"05", X"03", X"09", X"0d", X"0e", X"10", X"23", X"25", X"22", X"31", X"35", X"36", X"37", X"3d", X"41", X"45", X"42", X"3d", X"4a", X"44", X"46", X"48", X"3f", X"47", X"48", X"3a", X"3d", X"45", X"3c", X"40", X"39", X"3b", X"3c", X"39", X"35", X"42", X"40", X"37", X"37", X"3b", X"35", X"3b", X"39", X"36", X"3c", X"35", X"3b", X"3d", X"36", X"3e", X"46", X"43", X"51", X"61", X"70", X"7b", X"8a", X"89", X"89", X"8e", X"86", X"8c", X"89", X"85", X"80", X"7c", X"82", X"88", X"79", X"5e", X"18", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0f", X"4a", X"62", X"62", X"5f", X"6a", X"65", X"64", X"66", X"61", X"67", X"68", X"6d", X"6e", X"62", X"6a", X"68", X"65", X"67", X"64", X"65", X"6b", X"63", X"67", X"64", X"6a", X"63", X"61", X"63", X"68", X"65", X"5e", X"56", X"61", X"5d", X"58", X"62", X"5c", X"66", X"63", X"5e", X"5f", X"50", X"53", X"54", X"4c", X"4e", X"4d", X"45", X"40", X"3a", X"30", X"30", X"30", X"27", X"27", X"1b", X"11", X"1d", X"16", X"10", X"05", X"06", X"05", X"0e", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"07", X"03", X"0d", X"07", X"0f", X"0f", X"1f", X"22", X"24", X"2e", X"34", X"30", X"40", X"37", X"39", X"40", X"4c", X"3a", X"3a", X"4b", X"41", X"48", X"52", X"41", X"4d", X"43", X"3f", X"37", X"3c", X"45", X"39", X"44", X"3d", X"35", X"38", X"36", X"3b", X"3e", X"3a", X"3c", X"38", X"33", X"37", X"34", X"41", X"36", X"3a", X"3f", X"35", X"41", X"47", X"4b", X"53", X"6a", X"76", X"82", X"8e", X"85", X"94", X"8d", X"87", X"85", X"83", X"83", X"7b", X"7d", X"77", X"83", X"75", X"61", X"19", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"0c", X"49", X"60", X"65", X"63", X"64", X"6b", X"64", X"66", X"61", X"65", X"64", X"63", X"65", X"66", X"6b", X"65", X"62", X"60", X"65", X"5d", X"68", X"63", X"65", X"63", X"64", X"64", X"62", X"69", X"67", X"65", X"65", X"5b", X"5d", X"61", X"5e", X"57", X"53", X"5c", X"57", X"55", X"56", X"51", X"4b", X"58", X"52", X"4c", X"47", X"3e", X"34", X"39", X"33", X"1e", X"31", X"24", X"22", X"20", X"13", X"11", X"14", X"09", X"07", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"09", X"0a", X"09", X"05", X"12", X"17", X"1d", X"24", X"29", X"31", X"37", X"39", X"3a", X"3a", X"3c", X"42", X"36", X"4a", X"3e", X"40", X"3f", X"46", X"4b", X"44", X"42", X"3e", X"45", X"3e", X"34", X"3d", X"3b", X"39", X"41", X"38", X"39", X"3d", X"39", X"3d", X"3a", X"40", X"37", X"33", X"3d", X"3d", X"3c", X"34", X"39", X"40", X"3e", X"46", X"52", X"63", X"70", X"75", X"80", X"88", X"88", X"8c", X"87", X"84", X"84", X"81", X"81", X"82", X"84", X"7d", X"7f", X"73", X"5b", X"22", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0e", X"42", X"5f", X"65", X"62", X"5f", X"6d", X"5e", X"60", X"67", X"5e", X"62", X"67", X"64", X"6d", X"64", X"61", X"64", X"66", X"66", X"57", X"5f", X"65", X"69", X"5a", X"67", X"62", X"5d", X"60", X"5d", X"5e", X"5e", X"58", X"59", X"59", X"5d", X"5d", X"56", X"58", X"60", X"55", X"5e", X"56", X"50", X"4b", X"50", X"4e", X"45", X"44", X"36", X"32", X"33", X"28", X"23", X"27", X"22", X"1e", X"12", X"15", X"09", X"04", X"0b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"04", X"06", X"0b", X"0e", X"12", X"1a", X"18", X"27", X"28", X"35", X"37", X"35", X"38", X"33", X"44", X"3a", X"49", X"3d", X"38", X"3a", X"3c", X"3b", X"43", X"3e", X"42", X"38", X"3f", X"3c", X"38", X"3d", X"37", X"3e", X"3f", X"3d", X"3f", X"3d", X"32", X"41", X"35", X"3e", X"3f", X"3c", X"3b", X"3c", X"3b", X"39", X"3f", X"44", X"43", X"58", X"63", X"76", X"7b", X"83", X"84", X"85", X"87", X"87", X"81", X"81", X"7c", X"8a", X"88", X"82", X"7a", X"7c", X"71", X"62", X"1d", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"10", X"45", X"5d", X"65", X"57", X"5b", X"5d", X"61", X"63", X"60", X"5f", X"6a", X"61", X"60", X"5d", X"60", X"62", X"63", X"59", X"62", X"61", X"65", X"5f", X"64", X"5e", X"61", X"5f", X"63", X"61", X"62", X"60", X"64", X"59", X"58", X"63", X"5c", X"5e", X"56", X"5c", X"54", X"53", X"54", X"51", X"52", X"47", X"43", X"43", X"3d", X"40", X"33", X"30", X"31", X"26", X"1e", X"1d", X"1d", X"18", X"0f", X"13", X"08", X"05", X"06", X"06", X"05", X"08", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0d", X"13", X"16", X"1b", X"29", X"23", X"2b", X"34", X"3c", X"33", X"39", X"38", X"3e", X"3d", X"3f", X"3c", X"3b", X"41", X"3a", X"44", X"40", X"3f", X"3e", X"3d", X"43", X"39", X"38", X"3f", X"3f", X"39", X"3b", X"3d", X"41", X"43", X"3e", X"39", X"43", X"36", X"34", X"3f", X"3d", X"41", X"3b", X"42", X"4a", X"51", X"56", X"67", X"79", X"7b", X"84", X"88", X"83", X"8a", X"83", X"7e", X"83", X"84", X"7f", X"7b", X"75", X"7b", X"73", X"74", X"64", X"27", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0a", X"3e", X"53", X"64", X"59", X"5b", X"57", X"59", X"5f", X"64", X"5e", X"64", X"5d", X"59", X"63", X"64", X"6a", X"5f", X"67", X"66", X"5e", X"5f", X"5b", X"67", X"66", X"65", X"62", X"5c", X"5d", X"5e", X"61", X"61", X"5a", X"58", X"61", X"5e", X"53", X"5b", X"54", X"58", X"59", X"54", X"54", X"4b", X"43", X"46", X"39", X"45", X"37", X"33", X"29", X"29", X"21", X"21", X"22", X"1e", X"1c", X"1b", X"0b", X"09", X"04", X"07", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"01", X"08", X"06", X"11", X"14", X"18", X"1a", X"20", X"21", X"25", X"31", X"3b", X"35", X"34", X"3b", X"3b", X"40", X"37", X"35", X"47", X"3e", X"40", X"3d", X"38", X"43", X"3d", X"3c", X"3f", X"3f", X"37", X"3c", X"37", X"3d", X"38", X"3e", X"45", X"36", X"35", X"37", X"37", X"38", X"3a", X"40", X"35", X"41", X"3f", X"3c", X"51", X"4f", X"66", X"78", X"79", X"7f", X"7f", X"86", X"8b", X"89", X"85", X"83", X"81", X"84", X"83", X"83", X"80", X"73", X"7b", X"72", X"5d", X"28", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"2f", X"54", X"5e", X"63", X"5f", X"65", X"60", X"59", X"62", X"5e", X"63", X"59", X"5f", X"60", X"62", X"64", X"5f", X"66", X"5e", X"62", X"66", X"5f", X"62", X"60", X"66", X"62", X"5a", X"61", X"5b", X"5d", X"5d", X"55", X"53", X"51", X"54", X"5b", X"5e", X"54", X"58", X"53", X"4d", X"4d", X"46", X"47", X"41", X"3c", X"3c", X"30", X"33", X"2a", X"24", X"1e", X"21", X"15", X"1c", X"12", X"0b", X"0a", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"07", X"06", X"0f", X"11", X"1d", X"16", X"25", X"2b", X"32", X"2d", X"35", X"3b", X"34", X"38", X"3a", X"40", X"3c", X"40", X"3d", X"34", X"3d", X"3a", X"3f", X"3d", X"3e", X"3d", X"3a", X"3e", X"3c", X"3a", X"3b", X"3b", X"3c", X"3e", X"38", X"45", X"40", X"3e", X"47", X"3c", X"3f", X"37", X"38", X"37", X"40", X"4c", X"5a", X"66", X"6f", X"7a", X"7a", X"85", X"89", X"82", X"81", X"86", X"7f", X"86", X"79", X"7f", X"75", X"78", X"75", X"73", X"6c", X"57", X"2f", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"2d", X"4f", X"54", X"5b", X"5b", X"60", X"60", X"5b", X"5d", X"64", X"5b", X"62", X"60", X"69", X"60", X"5d", X"5f", X"5c", X"61", X"65", X"66", X"5a", X"5c", X"5e", X"5f", X"5d", X"59", X"5c", X"65", X"5a", X"54", X"5a", X"56", X"5f", X"59", X"56", X"50", X"56", X"58", X"53", X"4f", X"53", X"4a", X"43", X"35", X"38", X"32", X"29", X"31", X"2d", X"28", X"24", X"1f", X"18", X"21", X"0e", X"10", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"02", X"06", X"05", X"08", X"0f", X"16", X"19", X"15", X"29", X"26", X"32", X"31", X"2d", X"3c", X"3a", X"31", X"3a", X"39", X"39", X"45", X"3b", X"3e", X"46", X"34", X"3e", X"41", X"3d", X"41", X"43", X"3e", X"38", X"3a", X"32", X"44", X"3e", X"3f", X"3f", X"41", X"3d", X"36", X"47", X"44", X"40", X"45", X"42", X"3c", X"48", X"42", X"5a", X"68", X"69", X"75", X"81", X"89", X"83", X"83", X"8a", X"86", X"84", X"84", X"85", X"85", X"82", X"7d", X"73", X"75", X"73", X"60", X"34", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"08", X"31", X"59", X"5d", X"54", X"5f", X"5d", X"5b", X"60", X"5c", X"69", X"65", X"63", X"60", X"56", X"58", X"63", X"5b", X"63", X"64", X"5c", X"5d", X"56", X"5a", X"5e", X"61", X"64", X"5c", X"5c", X"5b", X"59", X"57", X"5a", X"54", X"55", X"52", X"52", X"54", X"5c", X"56", X"59", X"4a", X"43", X"43", X"3c", X"3a", X"3b", X"33", X"2c", X"2c", X"2c", X"1e", X"22", X"1a", X"17", X"14", X"0d", X"0b", X"08", X"0a", X"03", X"06", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"08", X"07", X"0f", X"11", X"1c", X"22", X"25", X"21", X"28", X"30", X"2c", X"30", X"38", X"37", X"3b", X"38", X"3b", X"3a", X"37", X"3f", X"3e", X"3e", X"41", X"42", X"37", X"42", X"3f", X"40", X"38", X"3e", X"42", X"3d", X"3f", X"36", X"43", X"3a", X"3f", X"44", X"40", X"3d", X"40", X"3d", X"3f", X"48", X"4c", X"59", X"66", X"6a", X"78", X"75", X"83", X"7d", X"7b", X"84", X"84", X"82", X"83", X"7e", X"79", X"7f", X"76", X"72", X"77", X"6e", X"61", X"2e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"25", X"51", X"61", X"5b", X"5f", X"5b", X"5c", X"63", X"5e", X"61", X"57", X"5f", X"5e", X"59", X"5e", X"5f", X"62", X"59", X"56", X"57", X"5f", X"5a", X"60", X"66", X"53", X"5c", X"5a", X"62", X"59", X"56", X"5b", X"4e", X"5a", X"56", X"4d", X"51", X"5b", X"52", X"56", X"4c", X"46", X"42", X"47", X"3b", X"36", X"33", X"34", X"2c", X"2b", X"20", X"24", X"19", X"10", X"13", X"10", X"13", X"0b", X"09", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"06", X"06", X"08", X"0d", X"16", X"1f", X"1b", X"1c", X"20", X"24", X"28", X"34", X"35", X"35", X"39", X"2b", X"39", X"3a", X"40", X"3e", X"3d", X"3c", X"3a", X"40", X"3f", X"3d", X"45", X"43", X"3d", X"42", X"48", X"41", X"44", X"4a", X"50", X"48", X"45", X"45", X"47", X"46", X"3c", X"3e", X"42", X"49", X"4f", X"5d", X"66", X"67", X"77", X"76", X"7e", X"83", X"87", X"7b", X"80", X"7f", X"81", X"7d", X"7b", X"70", X"78", X"6d", X"70", X"71", X"68", X"35", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"2c", X"4f", X"5b", X"5c", X"62", X"60", X"5c", X"55", X"5c", X"64", X"5d", X"61", X"5a", X"56", X"5d", X"55", X"64", X"57", X"5c", X"59", X"58", X"61", X"5f", X"5e", X"60", X"51", X"58", X"57", X"54", X"4e", X"59", X"5a", X"58", X"53", X"50", X"56", X"53", X"51", X"48", X"48", X"47", X"3c", X"40", X"37", X"30", X"30", X"29", X"2a", X"24", X"24", X"23", X"15", X"11", X"0b", X"0f", X"0f", X"0c", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"08", X"07", X"0e", X"10", X"1f", X"1a", X"19", X"26", X"22", X"30", X"31", X"2f", X"34", X"34", X"34", X"3b", X"47", X"38", X"43", X"44", X"3c", X"41", X"3f", X"3c", X"3b", X"3e", X"47", X"41", X"41", X"44", X"47", X"4c", X"4c", X"48", X"4a", X"58", X"50", X"54", X"54", X"53", X"47", X"47", X"49", X"51", X"58", X"61", X"62", X"6f", X"70", X"86", X"83", X"85", X"7e", X"7c", X"7e", X"78", X"7d", X"7a", X"76", X"6e", X"73", X"75", X"69", X"5f", X"37", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"1f", X"4e", X"58", X"58", X"5d", X"59", X"52", X"58", X"5c", X"58", X"60", X"5a", X"5e", X"65", X"59", X"5c", X"5d", X"55", X"5c", X"5a", X"59", X"62", X"59", X"61", X"5e", X"58", X"5b", X"61", X"5e", X"62", X"62", X"5c", X"50", X"5b", X"59", X"53", X"4d", X"4b", X"46", X"48", X"44", X"3b", X"3b", X"36", X"2f", X"36", X"2a", X"29", X"20", X"24", X"1b", X"19", X"10", X"0d", X"0f", X"10", X"04", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"07", X"06", X"07", X"03", X"0c", X"06", X"0b", X"09", X"16", X"1d", X"16", X"22", X"27", X"27", X"37", X"35", X"2d", X"33", X"35", X"3a", X"36", X"3f", X"42", X"3e", X"47", X"41", X"49", X"4d", X"41", X"49", X"48", X"41", X"52", X"4b", X"4e", X"54", X"59", X"54", X"60", X"65", X"5e", X"54", X"56", X"57", X"51", X"53", X"51", X"50", X"53", X"59", X"55", X"6e", X"67", X"74", X"7b", X"7e", X"84", X"82", X"7b", X"74", X"7d", X"79", X"78", X"75", X"70", X"6c", X"65", X"65", X"3c", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"1b", X"4e", X"5f", X"57", X"5f", X"5a", X"5f", X"5f", X"5a", X"5e", X"60", X"59", X"5a", X"59", X"58", X"5c", X"5f", X"5c", X"66", X"57", X"62", X"58", X"57", X"52", X"5f", X"51", X"52", X"58", X"56", X"5b", X"54", X"57", X"57", X"5d", X"59", X"52", X"4f", X"4a", X"49", X"3b", X"3a", X"3e", X"25", X"3d", X"32", X"27", X"2e", X"21", X"1f", X"19", X"1f", X"15", X"14", X"10", X"0e", X"06", X"04", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"05", X"07", X"10", X"0d", X"0b", X"15", X"16", X"26", X"27", X"25", X"2c", X"34", X"2f", X"32", X"27", X"35", X"37", X"42", X"46", X"41", X"44", X"46", X"40", X"44", X"42", X"44", X"4a", X"49", X"42", X"42", X"4e", X"56", X"60", X"60", X"64", X"68", X"62", X"61", X"68", X"66", X"60", X"52", X"59", X"51", X"54", X"55", X"50", X"5f", X"6f", X"73", X"79", X"76", X"72", X"79", X"79", X"79", X"73", X"78", X"76", X"75", X"6e", X"6b", X"65", X"5d", X"3e", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"19", X"50", X"51", X"52", X"59", X"59", X"4f", X"56", X"54", X"5b", X"5d", X"58", X"5b", X"5a", X"5e", X"5e", X"5b", X"5c", X"53", X"54", X"5a", X"59", X"56", X"58", X"5a", X"57", X"5c", X"4e", X"5a", X"57", X"5d", X"50", X"54", X"59", X"4c", X"4e", X"54", X"44", X"41", X"43", X"39", X"3b", X"3a", X"28", X"29", X"28", X"25", X"18", X"20", X"13", X"18", X"16", X"10", X"09", X"0f", X"0a", X"05", X"09", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"06", X"06", X"05", X"03", X"09", X"08", X"09", X"05", X"11", X"0f", X"19", X"22", X"28", X"23", X"25", X"2b", X"34", X"33", X"32", X"30", X"37", X"3e", X"3b", X"4a", X"4f", X"52", X"47", X"48", X"4a", X"49", X"4d", X"48", X"48", X"4f", X"4e", X"55", X"62", X"5b", X"70", X"6f", X"66", X"65", X"66", X"6b", X"63", X"63", X"61", X"61", X"5e", X"55", X"5b", X"54", X"5e", X"65", X"6a", X"6a", X"77", X"76", X"75", X"73", X"6e", X"70", X"78", X"6d", X"6d", X"75", X"70", X"65", X"3b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"18", X"4a", X"58", X"56", X"50", X"5b", X"4f", X"5e", X"55", X"50", X"5b", X"55", X"5b", X"59", X"58", X"5b", X"56", X"5e", X"5c", X"57", X"5e", X"54", X"5d", X"53", X"5c", X"50", X"55", X"55", X"5a", X"55", X"5b", X"5d", X"58", X"59", X"51", X"48", X"4b", X"49", X"3c", X"3b", X"30", X"36", X"2f", X"26", X"2c", X"25", X"2d", X"26", X"1a", X"1f", X"14", X"12", X"19", X"0b", X"09", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"0c", X"0f", X"0c", X"0d", X"13", X"1c", X"1d", X"1f", X"27", X"23", X"2b", X"33", X"30", X"3b", X"31", X"39", X"3f", X"49", X"54", X"5b", X"5a", X"54", X"57", X"53", X"58", X"4a", X"4a", X"45", X"53", X"53", X"59", X"63", X"6b", X"6f", X"70", X"65", X"6a", X"6a", X"6b", X"63", X"6c", X"69", X"5f", X"5f", X"5f", X"55", X"54", X"65", X"5c", X"6a", X"6f", X"71", X"6d", X"70", X"71", X"6a", X"6f", X"66", X"74", X"6c", X"6b", X"55", X"44", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"10", X"40", X"5f", X"58", X"55", X"56", X"4c", X"52", X"56", X"50", X"50", X"53", X"56", X"50", X"54", X"55", X"55", X"59", X"5c", X"57", X"5a", X"56", X"5a", X"55", X"57", X"5d", X"4a", X"59", X"60", X"5b", X"57", X"55", X"56", X"55", X"49", X"51", X"49", X"3e", X"3a", X"31", X"35", X"2e", X"36", X"2d", X"2f", X"29", X"1d", X"21", X"1e", X"16", X"12", X"11", X"10", X"0b", X"05", X"0c", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"04", X"06", X"0c", X"04", X"06", X"0d", X"11", X"11", X"17", X"1d", X"2b", X"20", X"27", X"2f", X"25", X"31", X"30", X"37", X"38", X"46", X"49", X"51", X"5e", X"64", X"59", X"57", X"5a", X"51", X"4c", X"50", X"4d", X"54", X"51", X"65", X"63", X"64", X"6c", X"63", X"6f", X"6b", X"6b", X"61", X"62", X"66", X"68", X"62", X"5d", X"5c", X"50", X"53", X"57", X"5d", X"61", X"65", X"73", X"6b", X"6d", X"65", X"6c", X"6d", X"69", X"6c", X"6b", X"5e", X"3f", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"10", X"43", X"53", X"52", X"57", X"57", X"51", X"45", X"48", X"3b", X"3c", X"3c", X"41", X"44", X"49", X"58", X"53", X"52", X"59", X"5c", X"5a", X"58", X"58", X"57", X"56", X"4e", X"56", X"51", X"53", X"55", X"4c", X"57", X"51", X"4c", X"4b", X"3e", X"3d", X"40", X"3d", X"37", X"2e", X"2c", X"2d", X"2b", X"22", X"24", X"1c", X"23", X"18", X"14", X"0a", X"0c", X"06", X"06", X"05", X"03", X"01", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"10", X"08", X"0a", X"0b", X"0b", X"10", X"12", X"14", X"16", X"1f", X"1e", X"28", X"19", X"26", X"29", X"32", X"2d", X"3e", X"44", X"4a", X"47", X"54", X"5a", X"5f", X"5f", X"62", X"65", X"54", X"59", X"51", X"4b", X"4e", X"56", X"57", X"64", X"5d", X"69", X"62", X"6d", X"63", X"64", X"6f", X"67", X"64", X"6d", X"6a", X"63", X"59", X"4f", X"54", X"52", X"56", X"58", X"58", X"60", X"5e", X"5e", X"67", X"6a", X"66", X"69", X"6e", X"63", X"5f", X"4a", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0c", X"3c", X"54", X"52", X"5a", X"4f", X"4a", X"34", X"29", X"1d", X"24", X"18", X"25", X"1f", X"3c", X"57", X"53", X"5e", X"54", X"59", X"53", X"52", X"5e", X"5c", X"60", X"52", X"59", X"5a", X"50", X"56", X"59", X"4f", X"54", X"43", X"4d", X"40", X"3b", X"3e", X"3b", X"39", X"22", X"2e", X"26", X"2a", X"27", X"29", X"1f", X"1a", X"1f", X"15", X"18", X"0d", X"08", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"0e", X"13", X"13", X"15", X"1e", X"23", X"1e", X"26", X"27", X"2d", X"28", X"36", X"31", X"37", X"3c", X"3d", X"53", X"53", X"5f", X"63", X"6a", X"67", X"64", X"64", X"5e", X"5e", X"62", X"5e", X"5e", X"59", X"60", X"67", X"59", X"64", X"66", X"67", X"65", X"6b", X"65", X"69", X"6b", X"61", X"60", X"56", X"45", X"49", X"47", X"4a", X"53", X"5a", X"5a", X"56", X"5e", X"57", X"5f", X"64", X"62", X"62", X"57", X"42", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"11", X"3b", X"56", X"51", X"5b", X"3f", X"2e", X"17", X"09", X"06", X"05", X"03", X"09", X"11", X"1f", X"4a", X"52", X"5d", X"62", X"57", X"5e", X"5a", X"56", X"58", X"5c", X"4d", X"59", X"5a", X"51", X"58", X"50", X"4d", X"4d", X"49", X"4a", X"41", X"3a", X"34", X"2d", X"2c", X"25", X"2b", X"26", X"26", X"2a", X"1a", X"18", X"1d", X"0f", X"12", X"17", X"0b", X"00", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0c", X"0e", X"08", X"12", X"17", X"15", X"17", X"21", X"15", X"25", X"2c", X"33", X"34", X"35", X"3e", X"3a", X"43", X"4a", X"50", X"58", X"66", X"68", X"64", X"62", X"67", X"65", X"66", X"66", X"59", X"54", X"54", X"5a", X"5c", X"60", X"5f", X"5d", X"5e", X"5e", X"66", X"68", X"65", X"67", X"60", X"57", X"5b", X"42", X"48", X"3e", X"42", X"45", X"48", X"4a", X"4e", X"54", X"54", X"51", X"57", X"63", X"52", X"52", X"3b", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0e", X"3d", X"4b", X"3f", X"52", X"35", X"0a", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"2e", X"50", X"58", X"60", X"60", X"5f", X"5d", X"60", X"54", X"52", X"55", X"51", X"50", X"4a", X"52", X"58", X"4a", X"49", X"43", X"40", X"3a", X"38", X"29", X"2f", X"32", X"31", X"2d", X"25", X"24", X"1f", X"22", X"18", X"12", X"10", X"11", X"12", X"04", X"02", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"09", X"03", X"04", X"07", X"0a", X"0d", X"11", X"1e", X"11", X"19", X"1d", X"14", X"25", X"27", X"2b", X"2d", X"31", X"38", X"3f", X"46", X"51", X"52", X"5e", X"5e", X"63", X"66", X"6f", X"67", X"67", X"69", X"5f", X"5e", X"5e", X"50", X"54", X"5b", X"56", X"5a", X"57", X"58", X"5e", X"5d", X"60", X"5e", X"5c", X"5e", X"56", X"51", X"4c", X"37", X"41", X"3a", X"42", X"45", X"3e", X"40", X"49", X"51", X"4a", X"54", X"51", X"55", X"3d", X"10", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0e", X"39", X"46", X"4b", X"38", X"15", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"12", X"42", X"54", X"5c", X"59", X"5f", X"5a", X"61", X"5b", X"54", X"56", X"46", X"4d", X"50", X"55", X"4e", X"49", X"49", X"3e", X"37", X"34", X"35", X"3a", X"35", X"37", X"27", X"25", X"29", X"1a", X"18", X"16", X"1f", X"0c", X"0c", X"14", X"0c", X"0a", X"08", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0c", X"0a", X"09", X"15", X"13", X"11", X"16", X"21", X"18", X"1b", X"22", X"22", X"28", X"34", X"30", X"35", X"3a", X"3c", X"3d", X"4a", X"50", X"5a", X"63", X"60", X"66", X"65", X"64", X"6a", X"64", X"61", X"5f", X"4e", X"59", X"48", X"52", X"5c", X"56", X"58", X"61", X"62", X"59", X"54", X"5b", X"50", X"54", X"45", X"3b", X"36", X"36", X"3d", X"3d", X"47", X"3e", X"42", X"3f", X"3f", X"44", X"44", X"45", X"48", X"39", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0f", X"32", X"49", X"38", X"1c", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0d", X"40", X"54", X"5f", X"57", X"51", X"4d", X"52", X"56", X"50", X"55", X"4c", X"4c", X"59", X"4c", X"47", X"4e", X"3b", X"3f", X"38", X"2f", X"38", X"2b", X"2a", X"30", X"2c", X"24", X"28", X"1e", X"1d", X"15", X"17", X"11", X"14", X"12", X"05", X"06", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0a", X"06", X"05", X"0d", X"0e", X"15", X"14", X"0f", X"19", X"1a", X"1e", X"1f", X"2a", X"23", X"2b", X"34", X"3d", X"39", X"39", X"3f", X"4c", X"4d", X"4e", X"57", X"5b", X"61", X"62", X"6a", X"61", X"62", X"5b", X"54", X"55", X"44", X"47", X"4f", X"4e", X"4d", X"58", X"49", X"51", X"5a", X"4c", X"4c", X"49", X"42", X"3e", X"31", X"3b", X"37", X"36", X"3b", X"36", X"33", X"3c", X"36", X"36", X"3e", X"3f", X"3a", X"30", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"1b", X"2f", X"13", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0d", X"3e", X"53", X"54", X"5d", X"5e", X"52", X"61", X"53", X"54", X"4f", X"4c", X"53", X"4f", X"4c", X"45", X"40", X"39", X"2d", X"30", X"34", X"36", X"35", X"25", X"24", X"22", X"27", X"21", X"1b", X"17", X"19", X"0e", X"10", X"0c", X"0b", X"05", X"03", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"06", X"0d", X"0c", X"13", X"16", X"14", X"11", X"1e", X"1f", X"20", X"19", X"21", X"28", X"2b", X"30", X"33", X"31", X"3a", X"3a", X"3f", X"4c", X"4c", X"51", X"54", X"58", X"5f", X"5b", X"5c", X"5b", X"57", X"55", X"42", X"47", X"41", X"44", X"46", X"45", X"4b", X"4a", X"48", X"46", X"48", X"39", X"3f", X"41", X"34", X"35", X"39", X"2f", X"31", X"30", X"36", X"35", X"32", X"3c", X"38", X"34", X"33", X"2f", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"10", X"06", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"24", X"45", X"4f", X"5c", X"5b", X"54", X"55", X"52", X"49", X"4d", X"4f", X"46", X"45", X"4c", X"42", X"35", X"36", X"34", X"35", X"2b", X"2f", X"31", X"25", X"2b", X"2c", X"27", X"1e", X"18", X"18", X"18", X"13", X"0e", X"0b", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"07", X"06", X"05", X"12", X"0f", X"13", X"14", X"13", X"1a", X"15", X"14", X"24", X"24", X"2a", X"28", X"2a", X"28", X"2f", X"3a", X"40", X"3f", X"47", X"41", X"4a", X"49", X"4c", X"55", X"50", X"56", X"5d", X"55", X"5a", X"4f", X"45", X"48", X"4d", X"4d", X"4d", X"4e", X"48", X"46", X"3f", X"45", X"36", X"3d", X"3e", X"3b", X"32", X"38", X"39", X"38", X"30", X"32", X"3a", X"31", X"31", X"33", X"39", X"3b", X"32", X"26", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"0b", X"0b", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"1a", X"37", X"51", X"5b", X"57", X"52", X"51", X"4c", X"57", X"4e", X"46", X"40", X"3d", X"46", X"39", X"39", X"37", X"37", X"32", X"2b", X"2b", X"37", X"28", X"2e", X"2b", X"20", X"1a", X"1f", X"1e", X"16", X"16", X"0c", X"08", X"0f", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"08", X"03", X"05", X"09", X"12", X"0d", X"11", X"1f", X"14", X"21", X"1f", X"20", X"1f", X"22", X"2f", X"2e", X"30", X"39", X"30", X"33", X"40", X"38", X"3e", X"44", X"46", X"4c", X"4b", X"57", X"53", X"50", X"4f", X"4e", X"4f", X"48", X"4f", X"4d", X"45", X"4c", X"4a", X"4c", X"3c", X"3c", X"3b", X"37", X"3f", X"35", X"3c", X"35", X"32", X"35", X"32", X"36", X"2f", X"35", X"2b", X"3c", X"36", X"2f", X"20", X"0c", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0f", X"1c", X"2a", X"1f", X"0d", X"07", X"03", X"06", X"05", X"05", X"06", X"17", X"39", X"3a", X"4b", X"52", X"4f", X"51", X"45", X"4e", X"51", X"4b", X"4b", X"48", X"3b", X"41", X"38", X"36", X"34", X"31", X"2e", X"2d", X"35", X"2c", X"1e", X"2f", X"25", X"2a", X"1e", X"15", X"16", X"19", X"08", X"16", X"06", X"0a", X"0c", X"06", X"05", X"03", X"01", X"06", X"05", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"0e", X"07", X"07", X"06", X"0c", X"13", X"16", X"17", X"11", X"15", X"15", X"16", X"22", X"26", X"21", X"28", X"2a", X"2f", X"31", X"35", X"35", X"33", X"30", X"3c", X"40", X"40", X"48", X"4c", X"4a", X"51", X"49", X"45", X"45", X"4c", X"45", X"44", X"41", X"3c", X"40", X"42", X"44", X"41", X"37", X"36", X"35", X"33", X"3b", X"34", X"3d", X"35", X"2f", X"2c", X"31", X"30", X"28", X"31", X"34", X"2b", X"2d", X"0c", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"09", X"2c", X"39", X"49", X"3a", X"2b", X"24", X"19", X"09", X"17", X"1c", X"2b", X"3a", X"48", X"49", X"49", X"4d", X"48", X"42", X"46", X"47", X"49", X"4c", X"45", X"36", X"3e", X"2e", X"36", X"2e", X"29", X"34", X"2b", X"30", X"25", X"28", X"26", X"23", X"1f", X"1d", X"1f", X"1e", X"16", X"06", X"0c", X"07", X"05", X"04", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"09", X"0a", X"0a", X"10", X"14", X"0e", X"15", X"14", X"15", X"1e", X"1f", X"1e", X"25", X"25", X"2c", X"2f", X"2b", X"33", X"37", X"30", X"35", X"39", X"34", X"43", X"37", X"47", X"45", X"41", X"44", X"40", X"47", X"4f", X"4a", X"4a", X"42", X"42", X"44", X"43", X"46", X"40", X"37", X"3a", X"38", X"33", X"3f", X"34", X"36", X"2e", X"29", X"33", X"31", X"32", X"33", X"37", X"32", X"38", X"28", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"13", X"41", X"38", X"3d", X"45", X"41", X"38", X"34", X"35", X"33", X"3c", X"3a", X"3b", X"44", X"43", X"4f", X"45", X"48", X"46", X"41", X"4a", X"43", X"43", X"42", X"36", X"37", X"35", X"33", X"30", X"33", X"35", X"30", X"2d", X"29", X"28", X"25", X"24", X"1d", X"21", X"1a", X"1a", X"12", X"10", X"0f", X"07", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"08", X"05", X"03", X"0a", X"06", X"09", X"08", X"14", X"13", X"10", X"10", X"18", X"1c", X"20", X"1a", X"23", X"22", X"24", X"30", X"2f", X"29", X"32", X"35", X"32", X"33", X"39", X"35", X"36", X"3f", X"35", X"3c", X"43", X"42", X"44", X"43", X"44", X"47", X"46", X"3f", X"46", X"3e", X"3f", X"44", X"44", X"35", X"35", X"39", X"39", X"2d", X"30", X"32", X"31", X"2d", X"29", X"30", X"30", X"2e", X"35", X"2b", X"26", X"07", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"1c", X"3c", X"36", X"37", X"45", X"3d", X"3f", X"45", X"3c", X"42", X"36", X"3e", X"3f", X"44", X"46", X"47", X"46", X"3a", X"3f", X"41", X"40", X"3f", X"38", X"3d", X"37", X"32", X"31", X"26", X"2d", X"29", X"33", X"2a", X"2c", X"2d", X"2d", X"2b", X"28", X"19", X"1c", X"18", X"10", X"13", X"07", X"04", X"09", X"07", X"03", X"01", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"0b", X"0a", X"0c", X"09", X"06", X"0e", X"13", X"1a", X"15", X"11", X"1f", X"1d", X"21", X"22", X"27", X"29", X"2a", X"26", X"34", X"2f", X"2b", X"31", X"33", X"39", X"36", X"3e", X"3d", X"35", X"3b", X"3e", X"45", X"3e", X"40", X"40", X"3d", X"3f", X"44", X"3f", X"33", X"39", X"3e", X"3e", X"2f", X"37", X"38", X"2e", X"30", X"31", X"30", X"32", X"2c", X"2f", X"2c", X"2f", X"2b", X"21", X"0c", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"11", X"33", X"37", X"42", X"3e", X"3b", X"30", X"3c", X"3f", X"3e", X"3d", X"3b", X"3e", X"3c", X"38", X"42", X"40", X"42", X"3e", X"3f", X"41", X"42", X"39", X"38", X"32", X"30", X"29", X"31", X"2c", X"2d", X"2e", X"2b", X"31", X"2d", X"2a", X"1e", X"16", X"16", X"17", X"16", X"15", X"14", X"0c", X"0e", X"06", X"05", X"0a", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"03", X"0a", X"05", X"05", X"09", X"09", X"0e", X"17", X"12", X"15", X"12", X"0f", X"1d", X"1e", X"25", X"2a", X"24", X"29", X"2c", X"2f", X"2d", X"2c", X"38", X"27", X"30", X"32", X"33", X"2f", X"30", X"31", X"37", X"43", X"42", X"47", X"3f", X"44", X"43", X"40", X"44", X"3c", X"38", X"3f", X"38", X"35", X"39", X"33", X"35", X"30", X"33", X"2f", X"29", X"30", X"29", X"2d", X"2f", X"29", X"28", X"10", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"36", X"37", X"41", X"3f", X"3d", X"3b", X"39", X"43", X"3d", X"41", X"3e", X"3c", X"41", X"43", X"44", X"40", X"3b", X"3f", X"3d", X"36", X"3e", X"39", X"35", X"2f", X"32", X"2c", X"30", X"2d", X"2f", X"32", X"27", X"29", X"1d", X"1c", X"1e", X"18", X"1b", X"17", X"0e", X"13", X"06", X"0c", X"01", X"06", X"05", X"08", X"01", X"06", X"08", X"03", X"09", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"07", X"06", X"05", X"03", X"07", X"0a", X"0f", X"11", X"0d", X"18", X"11", X"1a", X"1a", X"1e", X"22", X"23", X"22", X"29", X"30", X"21", X"2e", X"2e", X"26", X"28", X"30", X"31", X"33", X"2e", X"3b", X"30", X"39", X"37", X"39", X"44", X"43", X"3b", X"46", X"3c", X"40", X"41", X"3b", X"3b", X"3a", X"38", X"2f", X"2c", X"3a", X"28", X"33", X"32", X"35", X"2b", X"31", X"32", X"28", X"21", X"25", X"0f", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"07", X"2c", X"34", X"36", X"3e", X"36", X"3b", X"41", X"3b", X"40", X"3c", X"41", X"41", X"43", X"42", X"41", X"3f", X"42", X"40", X"38", X"34", X"33", X"32", X"38", X"30", X"2b", X"28", X"29", X"29", X"35", X"29", X"23", X"20", X"21", X"22", X"1c", X"1b", X"14", X"0e", X"10", X"08", X"06", X"03", X"03", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"04", X"0e", X"0a", X"05", X"14", X"14", X"17", X"12", X"16", X"18", X"12", X"20", X"1f", X"2a", X"20", X"27", X"2f", X"24", X"25", X"2c", X"26", X"2b", X"2e", X"2d", X"32", X"32", X"30", X"35", X"37", X"36", X"3b", X"3b", X"42", X"3a", X"40", X"3d", X"3c", X"37", X"42", X"3e", X"35", X"38", X"2e", X"2f", X"2f", X"2e", X"34", X"2d", X"2e", X"2a", X"2a", X"2b", X"26", X"2b", X"0e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"30", X"36", X"3f", X"3a", X"3c", X"44", X"43", X"3c", X"3e", X"3c", X"3f", X"3c", X"3b", X"3f", X"3a", X"3b", X"3e", X"37", X"3c", X"32", X"31", X"31", X"2c", X"2b", X"24", X"28", X"2a", X"21", X"2a", X"27", X"1f", X"1c", X"17", X"18", X"12", X"0f", X"12", X"10", X"09", X"08", X"06", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"07", X"06", X"09", X"0f", X"16", X"12", X"10", X"11", X"18", X"17", X"1e", X"16", X"1c", X"24", X"2b", X"22", X"26", X"2a", X"2a", X"32", X"29", X"2d", X"2c", X"27", X"31", X"2e", X"33", X"39", X"30", X"3c", X"3a", X"36", X"3b", X"3f", X"44", X"3e", X"36", X"40", X"43", X"46", X"34", X"31", X"2d", X"2b", X"32", X"2d", X"2f", X"28", X"2f", X"28", X"35", X"2c", X"22", X"0c", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"08", X"31", X"31", X"3b", X"43", X"3f", X"38", X"3e", X"38", X"3a", X"39", X"41", X"41", X"45", X"3a", X"41", X"37", X"36", X"3d", X"3a", X"2a", X"2e", X"24", X"2e", X"27", X"29", X"28", X"24", X"26", X"2a", X"24", X"22", X"20", X"18", X"13", X"18", X"0e", X"09", X"11", X"0b", X"06", X"05", X"03", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"09", X"09", X"14", X"0e", X"11", X"0b", X"11", X"18", X"14", X"1b", X"21", X"22", X"24", X"1f", X"25", X"26", X"28", X"22", X"28", X"27", X"2a", X"2b", X"2e", X"2e", X"29", X"28", X"31", X"32", X"2e", X"36", X"3f", X"34", X"3f", X"37", X"40", X"3d", X"3a", X"41", X"3e", X"40", X"33", X"2e", X"2f", X"2f", X"28", X"2d", X"30", X"2e", X"33", X"2d", X"28", X"1f", X"15", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"32", X"34", X"34", X"37", X"3a", X"39", X"33", X"43", X"3d", X"30", X"37", X"40", X"38", X"3c", X"3c", X"38", X"3d", X"39", X"2f", X"2c", X"2e", X"2a", X"26", X"29", X"20", X"26", X"2e", X"1d", X"20", X"1d", X"21", X"13", X"17", X"15", X"10", X"13", X"15", X"0d", X"08", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"0b", X"12", X"06", X"0d", X"0f", X"0b", X"10", X"16", X"18", X"19", X"18", X"1d", X"24", X"24", X"1f", X"28", X"26", X"20", X"1e", X"29", X"24", X"29", X"2b", X"2e", X"2a", X"29", X"26", X"2d", X"33", X"3e", X"35", X"32", X"41", X"34", X"35", X"33", X"3a", X"39", X"35", X"31", X"2d", X"2a", X"27", X"2e", X"2d", X"21", X"2d", X"28", X"22", X"25", X"10", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"30", X"30", X"36", X"34", X"32", X"33", X"36", X"39", X"3a", X"33", X"2f", X"34", X"38", X"36", X"36", X"2b", X"32", X"2f", X"2c", X"25", X"27", X"28", X"29", X"1f", X"1d", X"1c", X"24", X"22", X"21", X"1c", X"1d", X"10", X"19", X"0c", X"08", X"09", X"08", X"07", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"07", X"05", X"04", X"06", X"06", X"05", X"0d", X"0b", X"06", X"05", X"06", X"11", X"17", X"14", X"16", X"15", X"16", X"1b", X"26", X"27", X"1f", X"1e", X"24", X"24", X"26", X"2e", X"29", X"28", X"1a", X"26", X"2e", X"2c", X"32", X"36", X"2c", X"35", X"30", X"35", X"3a", X"39", X"33", X"31", X"34", X"34", X"36", X"36", X"31", X"2e", X"2c", X"38", X"26", X"26", X"32", X"23", X"21", X"1e", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"30", X"37", X"35", X"3b", X"34", X"33", X"2d", X"32", X"2b", X"36", X"36", X"33", X"2f", X"35", X"2b", X"24", X"24", X"2f", X"2f", X"25", X"24", X"1f", X"29", X"23", X"1e", X"20", X"25", X"23", X"21", X"1e", X"1b", X"1d", X"15", X"07", X"06", X"0c", X"0b", X"03", X"00", X"0f", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"04", X"06", X"07", X"09", X"04", X"06", X"09", X"11", X"12", X"11", X"10", X"12", X"1d", X"1a", X"20", X"1a", X"25", X"22", X"22", X"2d", X"27", X"2a", X"25", X"26", X"2e", X"2e", X"26", X"30", X"28", X"28", X"2d", X"2b", X"2d", X"32", X"31", X"31", X"39", X"3b", X"3d", X"3a", X"39", X"37", X"2c", X"34", X"2f", X"31", X"31", X"2f", X"2b", X"34", X"35", X"23", X"2a", X"1b", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"28", X"2f", X"2f", X"36", X"35", X"29", X"3a", X"2f", X"33", X"32", X"2e", X"2f", X"32", X"2c", X"2b", X"2c", X"25", X"25", X"23", X"29", X"29", X"20", X"1f", X"1f", X"25", X"21", X"21", X"22", X"1b", X"10", X"10", X"0d", X"05", X"13", X"0e", X"07", X"08", X"03", X"00", X"0a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"0f", X"07", X"0c", X"05", X"0b", X"09", X"10", X"0d", X"16", X"16", X"12", X"0a", X"20", X"17", X"22", X"20", X"1f", X"25", X"27", X"2b", X"25", X"2a", X"23", X"25", X"25", X"27", X"2f", X"29", X"2d", X"2f", X"25", X"2d", X"2a", X"2b", X"34", X"34", X"30", X"24", X"2a", X"32", X"2f", X"39", X"2e", X"30", X"27", X"32", X"34", X"21", X"27", X"1b", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"24", X"20", X"3a", X"36", X"26", X"2b", X"2b", X"2d", X"37", X"38", X"2f", X"2b", X"2b", X"29", X"26", X"24", X"27", X"2b", X"22", X"23", X"29", X"1e", X"23", X"28", X"1d", X"24", X"20", X"17", X"16", X"11", X"0b", X"14", X"05", X"07", X"03", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"03", X"06", X"05", X"03", X"00", X"06", X"09", X"09", X"0d", X"07", X"0d", X"0c", X"13", X"17", X"1a", X"15", X"10", X"13", X"1b", X"20", X"29", X"20", X"19", X"21", X"1e", X"28", X"28", X"24", X"21", X"28", X"24", X"29", X"2c", X"29", X"22", X"28", X"2e", X"33", X"38", X"2d", X"2a", X"31", X"2b", X"2d", X"2f", X"2d", X"2a", X"25", X"2d", X"2f", X"25", X"27", X"1d", X"11", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"14", X"2b", X"27", X"23", X"2b", X"24", X"25", X"2e", X"24", X"28", X"30", X"23", X"23", X"29", X"20", X"29", X"2c", X"24", X"23", X"1c", X"24", X"1a", X"24", X"1d", X"19", X"19", X"1b", X"14", X"11", X"15", X"0a", X"10", X"10", X"08", X"09", X"06", X"06", X"08", X"05", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"06", X"07", X"0a", X"05", X"03", X"07", X"09", X"14", X"11", X"10", X"14", X"14", X"14", X"14", X"1a", X"19", X"1d", X"15", X"21", X"22", X"20", X"27", X"27", X"22", X"23", X"20", X"23", X"23", X"26", X"29", X"26", X"1b", X"27", X"29", X"32", X"30", X"27", X"2c", X"27", X"2c", X"2a", X"2d", X"29", X"2a", X"2e", X"31", X"32", X"26", X"26", X"20", X"1e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"14", X"25", X"2d", X"28", X"25", X"29", X"2b", X"28", X"29", X"28", X"21", X"2a", X"25", X"28", X"16", X"25", X"21", X"23", X"24", X"27", X"20", X"2b", X"1f", X"10", X"1f", X"16", X"1e", X"12", X"0f", X"0e", X"0c", X"0b", X"0b", X"05", X"0b", X"06", X"05", X"06", X"00", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"05", X"01", X"06", X"05", X"05", X"04", X"07", X"0b", X"10", X"11", X"18", X"13", X"0a", X"13", X"12", X"1b", X"21", X"1b", X"17", X"22", X"1e", X"1a", X"1d", X"23", X"25", X"27", X"21", X"23", X"24", X"24", X"2a", X"25", X"25", X"22", X"2b", X"28", X"22", X"30", X"27", X"25", X"2d", X"25", X"23", X"29", X"20", X"2f", X"27", X"2d", X"25", X"30", X"21", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"17", X"21", X"27", X"29", X"1d", X"25", X"29", X"24", X"25", X"23", X"22", X"1e", X"23", X"24", X"21", X"22", X"22", X"1a", X"20", X"26", X"1f", X"1f", X"1b", X"18", X"19", X"12", X"15", X"10", X"12", X"0d", X"06", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"00", X"06", X"13", X"0c", X"0d", X"0f", X"14", X"14", X"14", X"0f", X"13", X"17", X"16", X"14", X"1c", X"1e", X"25", X"18", X"22", X"1a", X"1f", X"1b", X"17", X"20", X"24", X"23", X"21", X"27", X"25", X"1f", X"26", X"28", X"2d", X"22", X"2c", X"21", X"20", X"25", X"25", X"2b", X"28", X"21", X"2b", X"1f", X"24", X"1a", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"11", X"18", X"25", X"22", X"14", X"23", X"24", X"1b", X"26", X"21", X"17", X"1a", X"1c", X"1f", X"19", X"20", X"2b", X"12", X"1c", X"20", X"1e", X"11", X"18", X"0b", X"08", X"0d", X"08", X"0e", X"0b", X"03", X"00", X"06", X"06", X"05", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"0d", X"0b", X"0d", X"05", X"05", X"07", X"13", X"0f", X"0a", X"09", X"13", X"17", X"15", X"16", X"1b", X"17", X"11", X"1c", X"1a", X"22", X"21", X"1c", X"18", X"1a", X"1f", X"21", X"21", X"1d", X"28", X"1d", X"28", X"25", X"1d", X"25", X"22", X"28", X"1f", X"22", X"21", X"25", X"27", X"20", X"26", X"22", X"21", X"1d", X"18", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"13", X"1f", X"1f", X"21", X"1d", X"1a", X"21", X"22", X"27", X"1a", X"22", X"15", X"1b", X"1b", X"1f", X"21", X"1b", X"18", X"1b", X"15", X"14", X"14", X"14", X"0f", X"0f", X"0d", X"0f", X"0b", X"05", X"03", X"05", X"06", X"05", X"0a", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"0a", X"10", X"05", X"07", X"0a", X"0c", X"12", X"10", X"0a", X"0f", X"0b", X"12", X"16", X"16", X"16", X"0d", X"12", X"1e", X"1a", X"13", X"1a", X"17", X"20", X"1d", X"1f", X"23", X"24", X"17", X"24", X"1f", X"21", X"25", X"1e", X"1f", X"1d", X"26", X"23", X"1b", X"23", X"16", X"1e", X"1c", X"1a", X"19", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"12", X"14", X"10", X"0b", X"11", X"10", X"1f", X"15", X"13", X"19", X"1d", X"13", X"0e", X"13", X"16", X"16", X"12", X"18", X"0b", X"14", X"10", X"0e", X"09", X"05", X"03", X"06", X"0d", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"04", X"00", X"06", X"05", X"0d", X"00", X"06", X"09", X"03", X"05", X"06", X"06", X"0f", X"0c", X"0c", X"0f", X"08", X"0c", X"06", X"10", X"0b", X"0c", X"0f", X"13", X"16", X"1a", X"1b", X"16", X"1b", X"12", X"18", X"1e", X"11", X"1e", X"1f", X"1f", X"1c", X"16", X"17", X"1d", X"16", X"16", X"1b", X"15", X"16", X"10", X"0e", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"0c", X"0a", X"0c", X"07", X"0a", X"0e", X"0a", X"09", X"0c", X"0a", X"09", X"05", X"17", X"11", X"09", X"0f", X"0b", X"0a", X"06", X"0a", X"09", X"02", X"06", X"05", X"04", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"08", X"03", X"00", X"09", X"05", X"10", X"09", X"06", X"08", X"0b", X"07", X"07", X"09", X"03", X"03", X"06", X"09", X"0b", X"09", X"09", X"11", X"16", X"0f", X"13", X"14", X"0f", X"19", X"15", X"19", X"17", X"1c", X"20", X"1a", X"14", X"13", X"13", X"10", X"14", X"13", X"12", X"14", X"11", X"08", X"09", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"05", X"06", X"05", X"03", X"03", X"0d", X"05", X"0c", X"07", X"0a", X"05", X"06", X"04", X"06", X"06", X"03", X"01", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"01", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"07", X"05", X"06", X"05", X"05", X"04", X"06", X"05", X"03", X"00", X"06", X"05", X"05", X"00", X"06", X"05", X"07", X"0a", X"0a", X"08", X"05", X"08", X"0f", X"0c", X"06", X"12", X"0a", X"07", X"12", X"0d", X"0c", X"0b", X"0c", X"04", X"08", X"0b", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"06", X"03", X"0b", X"06", X"05", X"06", X"00", X"08", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"02", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"),
(X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05", X"03", X"00", X"06", X"05"));