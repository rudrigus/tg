 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 07 07 07 07 07 07 18 18 18 26 26 26 19 19 19 15 15 15 22 22 22 1a 1a 1a 0b 0b 0b 09 09 09 08 08 08 0a 0a 0a 09 09 09 05 05 05 05 05 05 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 0c 0c 0c 10 10 10 26 26 26 42 42 42 5f 5f 5f 6c 6c 6c 5d 5d 5d 5d 5d 5d 47 47 47 48 48 48 3d 3d 3d 38 38 38 3d 3d 3d 43 43 43 46 46 46 3f 3f 3f 2c 2c 2c 22 22 22 15 15 15 0d 0d 0d 08 08 08 07 07 07 05 05 05 05 05 05 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 04 04 04 05 05 05 08 08 08 0e 0e 0e 24 24 24 45 45 45 4a 4a 4a 78 78 78 83 83 83 79 79 79 7b 7b 7b 7d 7d 7d 84 84 84 88 88 88 70 70 70 5e 5e 5e 70 70 70 7b 7b 7b 8a 8a 8a 93 93 93 90 90 90 7e 7e 7e 6b 6b 6b 68 68 68 6d 6d 6d 52 52 52 30 30 30 17 17 17 0b 0b 0b 07 07 07 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 0a 0a 0a 16 16 16 31 31 31 4f 4f 4f 48 48 48 5f 5f 5f 6d 6d 6d 78 78 78 7e 7e 7e 89 89 89 8e 8e 8e 8b 8b 8b 84 84 84 8e 8e 8e 89 89 89 98 98 98 d1 d1 d1 bb bb bb b5 b5 b5 be be be bc bc bc b5 b5 b5 ac ac ac ad ad ad ab ab ab ad ad ad b6 b6 b6 c8 c8 c8 a0 a0 a0 5d 5d 5d 39 39 39 1d 1d 1d 0c 0c 0c 06 06 06 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 05 05 05 0d 0d 0d 2f 2f 2f 60 60 60 8d 8d 8d 9f 9f 9f a8 a8 a8 a0 a0 a0 7a 7a 7a 74 74 74 87 87 87 8c 8c 8c 97 97 97 a7 a7 a7 a5 a5 a5 ae ae ae b3 b3 b3 cd cd cd f8 f8 f8 f8 f8 f8 e3 e3 e3 f1 f1 f1 ec ec ec e4 e4 e4 e3 e3 e3 e2 e2 e2 da da da d3 d3 d3 c9 c9 c9 b8 b8 b8 b2 b2 b2 ab ab ab a0 a0 a0 a0 a0 a0 7e 7e 7e 48 48 48 24 24 24 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 13 13 13 14 14 14 16 16 16 5d 5d 5d 9c 9c 9c bb bb bb d0 d0 d0 d4 d4 d4 cf cf cf df df df e8 e8 e8 e4 e4 e4 ec ec ec e6 e6 e6 eb eb eb ef ef ef e6 e6 e6 e8 e8 e8 f1 f1 f1 f9 f9 f9 f4 f4 f4 f6 f6 f6 fb fb fb ff ff ff fd fd fd fc fc fc fc fc fc f8 f8 f8 ec ec ec df df df cd cd cd bc bc bc b0 b0 b0 a0 a0 a0 96 96 96 8f 8f 8f 96 96 96 97 97 97 5a 5a 5a 1f 1f 1f 0f 0f 0f 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0e 0e 0e 1d 1d 1d 54 54 54 99 99 99 a4 a4 a4 c1 c1 c1 ee ee ee fe fe fe fc fc fc fe fe fe ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe ff ff ff fa fa fa ee ee ee d9 d9 d9 c0 c0 c0 a8 a8 a8 96 96 96 8d 8d 8d 85 85 85 79 79 79 6c 6c 6c 6e 6e 6e 5b 5b 5b 28 28 28 21 21 21 07 07 07 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0e 0e 0e 1c 1c 1c 58 58 58 a2 a2 a2 98 98 98 a8 a8 a8 be be be db db db f5 f5 f5 fc fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 d6 d6 d6 be be be b4 b4 b4 a9 a9 a9 9c 9c 9c 87 87 87 73 73 73 66 66 66 5c 5c 5c 63 63 63 68 68 68 4c 4c 4c 1c 1c 1c 07 07 07 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 12 12 12 29 29 29 5f 5f 5f 8d 8d 8d 93 93 93 a4 a4 a4 bd bd bd d4 d4 d4 e3 e3 e3 ee ee ee f9 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f3 f3 dd dd dd df df df d7 d7 d7 c6 c6 c6 aa aa aa 8e 8e 8e 7f 7f 7f 77 77 77 72 72 72 6a 6a 6a 62 62 62 6d 6d 6d 4b 4b 4b 24 24 24 06 06 06 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 20 20 20 49 49 49 77 77 77 84 84 84 8f 8f 8f a0 a0 a0 bb bb bb dc dc dc f8 f8 f8 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fb fb fb f1 f1 f1 db db db c3 c3 c3 ab ab ab 9d 9d 9d 93 93 93 8f 8f 8f 85 85 85 79 79 79 6a 6a 6a 66 66 66 81 81 81 57 57 57 1c 1c 1c 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 1d 1d 1d 41 41 41 65 65 65 71 71 71 80 80 80 9e 9e 9e b3 b3 b3 c6 c6 c6 df df df f3 f3 f3 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f9 f9 e2 e2 e2 c8 c8 c8 b6 b6 b6 aa aa aa a4 a4 a4 98 98 98 8f 8f 8f 88 88 88 7f 7f 7f 75 75 75 6f 6f 6f 7a 7a 7a 7d 7d 7d 32 32 32 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0f 0f 0f 3a 3a 3a 62 62 62 77 77 77 7a 7a 7a 9f 9f 9f aa aa aa b0 b0 b0 bb bb bb c9 c9 c9 da da da ed ed ed f7 f7 f7 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fa fa e5 e5 e5 d0 d0 d0 bc bc bc ad ad ad a4 a4 a4 9c 9c 9c 94 94 94 91 91 91 8b 8b 8b 82 82 82 78 78 78 6c 6c 6c 6c 6c 6c 90 90 90 46 46 46 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 2d 2d 2d 5f 5f 5f 73 73 73 69 69 69 85 85 85 8f 8f 8f 8b 8b 8b 99 99 99 ab ab ab be be be cd cd cd d7 d7 d7 de de de ec ec ec f9 f9 f9 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 e8 e8 e8 d3 d3 d3 bd bd bd af af af a5 a5 a5 9f 9f 9f a0 a0 a0 9a 9a 9a 8c 8c 8c 80 80 80 78 78 78 6f 6f 6f 6f 6f 6f 73 73 73 91 91 91 58 58 58 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 47 47 47 7a 7a 7a 7c 7c 7c 69 69 69 75 75 75 73 73 73 7d 7d 7d 90 90 90 a5 a5 a5 b0 b0 b0 b7 b7 b7 bd bd bd c6 c6 c6 d6 d6 d6 e0 e0 e0 e7 e7 e7 ee ee ee f6 f6 f6 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb ea ea ea d9 d9 d9 c8 c8 c8 ba ba ba b0 b0 b0 aa aa aa a5 a5 a5 a1 a1 a1 8e 8e 8e 7d 7d 7d 74 74 74 76 76 76 78 78 78 7a 7a 7a 7a 7a 7a 92 92 92 56 56 56 07 07 07 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0e 0e 0e 4d 4d 4d 6b 6b 6b 6f 6f 6f 5f 5f 5f 69 69 69 73 73 73 7f 7f 7f 8e 8e 8e 9b 9b 9b 99 99 99 a0 a0 a0 a9 a9 a9 b3 b3 b3 c3 c3 c3 d0 d0 d0 d0 d0 d0 c9 c9 c9 d5 d5 d5 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fd fd fd fb fb fb ee ee ee dc dc dc cf cf cf c1 c1 c1 b6 b6 b6 ab ab ab a1 a1 a1 9d 9d 9d 8d 8d 8d 82 82 82 7b 7b 7b 7b 7b 7b 81 81 81 84 84 84 86 86 86 84 84 84 99 99 99 4f 4f 4f 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 56 56 56 67 67 67 58 58 58 62 62 62 6a 6a 6a 74 74 74 81 81 81 8e 8e 8e 8c 8c 8c 8d 8d 8d 97 97 97 a0 a0 a0 ab ab ab b9 b9 b9 c6 c6 c6 c4 c4 c4 bd bd bd d1 d1 d1 ff ff ff f4 f4 f4 dc dc dc be be be c1 c1 c1 d9 d9 d9 f5 f5 f5 fe fe fe f5 f5 f5 ed ed ed e6 e6 e6 e1 e1 e1 dc dc dc d6 d6 d6 ce ce ce c5 c5 c5 bb bb bb b0 b0 b0 aa aa aa a1 a1 a1 99 99 99 92 92 92 87 87 87 84 84 84 86 86 86 87 87 87 8c 8c 8c 8b 8b 8b 88 88 88 98 98 98 3a 3a 3a 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 58 58 58 87 87 87 62 62 62 66 66 66 6d 6d 6d 72 72 72 78 78 78 89 89 89 78 78 78 83 83 83 91 91 91 9f 9f 9f a9 a9 a9 b6 b6 b6 bf bf bf bf bf bf ba ba ba dd dd dd fb fb fb 98 98 98 5a 5a 5a 49 49 49 46 46 46 52 52 52 7f 7f 7f e2 e2 e2 d6 d6 d6 cb cb cb c4 c4 c4 c3 c3 c3 c1 c1 c1 bf bf bf b8 b8 b8 b2 b2 b2 af af af a9 a9 a9 a4 a4 a4 99 99 99 8f 8f 8f 89 89 89 80 80 80 7e 7e 7e 7c 7c 7c 80 80 80 86 86 86 8c 8c 8c 86 86 86 97 97 97 34 34 34 05 05 05 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 11 11 11 5f 5f 5f 9c 9c 9c 72 72 72 63 63 63 65 65 65 6c 6c 6c 74 74 74 78 78 78 73 73 73 78 78 78 86 86 86 93 93 93 9f 9f 9f ad ad ad b5 b5 b5 b7 b7 b7 b5 b5 b5 dd dd dd d7 d7 d7 4c 4c 4c 2a 2a 2a 20 20 20 1e 1e 1e 26 26 26 3a 3a 3a 99 99 99 c7 c7 c7 bb bb bb b6 b6 b6 b2 b2 b2 b1 b1 b1 ae ae ae a7 a7 a7 a0 a0 a0 9e 9e 9e 9a 9a 9a 94 94 94 88 88 88 7e 7e 7e 79 79 79 71 71 71 70 70 70 71 71 71 71 71 71 7a 7a 7a 81 81 81 80 80 80 9b 9b 9b 47 47 47 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 1e 1e 1e 6f 6f 6f a5 a5 a5 6f 6f 6f 61 61 61 64 64 64 69 69 69 6c 6c 6c 6c 6c 6c 73 73 73 77 77 77 7d 7d 7d 86 86 86 8e 8e 8e 9f 9f 9f a7 a7 a7 ab ab ab b0 b0 b0 cd cd cd aa aa aa 27 27 27 10 10 10 0c 0c 0c 0b 0b 0b 0e 0e 0e 1e 1e 1e 7b 7b 7b bb bb bb b3 b3 b3 af af af a8 a8 a8 a2 a2 a2 9b 9b 9b 95 95 95 94 94 94 91 91 91 8e 8e 8e 88 88 88 7a 7a 7a 72 72 72 6f 6f 6f 6b 6b 6b 6b 6b 6b 6b 6b 6b 6b 6b 6b 70 70 70 76 76 76 7a 7a 7a 9a 9a 9a 5b 5b 5b 11 11 11 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 08 08 08 30 30 30 80 80 80 a2 a2 a2 64 64 64 67 67 67 61 61 61 5e 5e 5e 63 63 63 66 66 66 6a 6a 6a 74 74 74 7d 7d 7d 81 81 81 84 84 84 90 90 90 9b 9b 9b a3 a3 a3 a5 a5 a5 af af af c1 c1 c1 1d 1d 1d 07 07 07 06 06 06 05 05 05 06 06 06 11 11 11 6d 6d 6d b6 b6 b6 af af af a5 a5 a5 9e 9e 9e 97 97 97 91 91 91 8b 8b 8b 8a 8a 8a 87 87 87 84 84 84 7f 7f 7f 71 71 71 69 69 69 68 68 68 67 67 67 66 66 66 69 69 69 6a 6a 6a 69 69 69 69 69 69 72 72 72 87 87 87 6c 6c 6c 25 25 25 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0c 0c 0c 3e 3e 3e 8f 8f 8f 78 78 78 66 66 66 65 65 65 5b 5b 5b 5f 5f 5f 64 64 64 68 68 68 6b 6b 6b 6e 6e 6e 75 75 75 7c 7c 7c 7e 7e 7e 84 84 84 91 91 91 91 91 91 96 96 96 9d 9d 9d aa aa aa 27 27 27 04 04 04 04 04 04 03 03 03 04 04 04 0b 0b 0b 62 62 62 b4 b4 b4 a4 a4 a4 9e 9e 9e 99 99 99 90 90 90 8b 8b 8b 85 85 85 84 84 84 82 82 82 7c 7c 7c 77 77 77 68 68 68 65 65 65 64 64 64 62 62 62 65 65 65 66 66 66 65 65 65 63 63 63 62 62 62 69 69 69 6f 6f 6f 71 71 71 38 38 38 06 06 06 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0d 0d 0d 4b 4b 4b 92 92 92 73 73 73 6b 6b 6b 62 62 62 5f 5f 5f 64 64 64 67 67 67 68 68 68 68 68 68 6a 6a 6a 6c 6c 6c 74 74 74 77 77 77 7f 7f 7f 85 85 85 81 81 81 89 89 89 8b 8b 8b 88 88 88 26 26 26 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 4f 4f 4f a3 a3 a3 98 98 98 92 92 92 91 91 91 89 89 89 84 84 84 80 80 80 7f 7f 7f 7e 7e 7e 77 77 77 6f 6f 6f 63 63 63 62 62 62 61 61 61 5d 5d 5d 5f 5f 5f 5f 5f 5f 5e 5e 5e 5d 5d 5d 5a 5a 5a 5f 5f 5f 64 64 64 6e 6e 6e 45 45 45 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 12 12 12 58 58 58 95 95 95 7c 7c 7c 6d 6d 6d 63 63 63 63 63 63 66 66 66 65 65 65 66 66 66 65 65 65 66 66 66 67 67 67 68 68 68 76 76 76 7d 7d 7d 76 76 76 78 78 78 7b 7b 7b 83 83 83 81 81 81 2b 2b 2b 03 03 03 04 04 04 03 03 03 03 03 03 06 06 06 39 39 39 94 94 94 8a 8a 8a 88 88 88 87 87 87 86 86 86 7f 7f 7f 7d 7d 7d 7f 7f 7f 7b 7b 7b 78 78 78 6c 6c 6c 60 60 60 5d 5d 5d 5c 5c 5c 5a 5a 5a 59 59 59 5b 5b 5b 59 59 59 59 59 59 5a 5a 5a 5b 5b 5b 62 62 62 6d 6d 6d 4f 4f 4f 0b 0b 0b 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 13 13 13 61 61 61 90 90 90 79 79 79 6e 6e 6e 63 63 63 61 61 61 61 61 61 62 62 62 5e 5e 5e 60 60 60 63 63 63 62 62 62 61 61 61 70 70 70 76 76 76 6e 6e 6e 6f 6f 6f 76 76 76 73 73 73 76 76 76 32 32 32 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 2a 2a 2a 89 89 89 7f 7f 7f 7e 7e 7e 7e 7e 7e 7f 7f 7f 7b 7b 7b 7a 7a 7a 7c 7c 7c 7a 7a 7a 75 75 75 64 64 64 5d 5d 5d 59 59 59 58 58 58 59 59 59 56 56 56 57 57 57 58 58 58 5a 5a 5a 59 59 59 58 58 58 5d 5d 5d 69 69 69 53 53 53 0b 0b 0b 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 13 13 13 62 62 62 92 92 92 79 79 79 6a 6a 6a 61 61 61 61 61 61 61 61 61 5d 5d 5d 5c 5c 5c 5e 5e 5e 5f 5f 5f 61 61 61 5d 5d 5d 64 64 64 6f 6f 6f 70 70 70 6a 6a 6a 70 70 70 68 68 68 6e 6e 6e 35 35 35 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1e 1e 1e 80 80 80 73 73 73 75 75 75 79 79 79 77 77 77 78 78 78 79 79 79 78 78 78 75 75 75 6e 6e 6e 5e 5e 5e 5a 5a 5a 57 57 57 57 57 57 56 56 56 54 54 54 56 56 56 59 59 59 59 59 59 59 59 59 59 59 59 55 55 55 62 62 62 5b 5b 5b 0e 0e 0e 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0f 0f 0f 5e 5e 5e 8e 8e 8e 90 90 90 86 86 86 61 61 61 5f 5f 5f 5e 5e 5e 5d 5d 5d 5c 5c 5c 5d 5d 5d 5c 5c 5c 5d 5d 5d 5a 5a 5a 5a 5a 5a 5c 5c 5c 64 64 64 66 66 66 6d 6d 6d 66 66 66 6a 6a 6a 3a 3a 3a 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 16 16 16 83 83 83 70 70 70 70 70 70 74 74 74 73 73 73 76 76 76 74 74 74 76 76 76 70 70 70 62 62 62 5b 5b 5b 5a 5a 5a 53 53 53 54 54 54 54 54 54 57 57 57 58 58 58 5a 5a 5a 58 58 58 56 56 56 58 58 58 55 55 55 63 63 63 58 58 58 0c 0c 0c 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 08 08 08 51 51 51 83 83 83 75 75 75 81 81 81 7a 7a 7a 60 60 60 5a 5a 5a 5c 5c 5c 5c 5c 5c 59 59 59 57 57 57 59 59 59 57 57 57 54 54 54 54 54 54 5a 5a 5a 63 63 63 74 74 74 64 64 64 63 63 63 3b 3b 3b 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 0e 0e 0e 79 79 79 7d 7d 7d 75 75 75 74 74 74 70 70 70 70 70 70 6e 6e 6e 6d 6d 6d 63 63 63 5b 5b 5b 59 59 59 56 56 56 53 53 53 53 53 53 53 53 53 54 54 54 58 58 58 57 57 57 56 56 56 55 55 55 55 55 55 54 54 54 65 65 65 48 48 48 07 07 07 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 06 06 06 3a 3a 3a 81 81 81 69 69 69 6d 6d 6d 7f 7f 7f 62 62 62 56 56 56 5a 5a 5a 56 56 56 54 54 54 54 54 54 54 54 54 56 56 56 52 52 52 51 51 51 55 55 55 5a 5a 5a 61 61 61 64 64 64 60 60 60 3f 3f 3f 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 09 09 09 77 77 77 7f 7f 7f 74 74 74 75 75 75 76 76 76 74 74 74 6b 6b 6b 61 61 61 59 59 59 58 58 58 59 59 59 54 54 54 52 52 52 50 50 50 51 51 51 54 54 54 56 56 56 58 58 58 56 56 56 55 55 55 55 55 55 58 58 58 54 54 54 27 27 27 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 05 05 05 1c 1c 1c 72 72 72 61 61 61 66 66 66 6a 6a 6a 5f 5f 5f 54 54 54 57 57 57 55 55 55 52 52 52 52 52 52 54 54 54 53 53 53 4f 4f 4f 51 51 51 52 52 52 59 59 59 5b 5b 5b 61 61 61 60 60 60 45 45 45 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 73 73 73 7a 7a 7a 70 70 70 6d 6d 6d 6e 6e 6e 73 73 73 6a 6a 6a 5d 5d 5d 58 58 58 57 57 57 57 57 57 55 55 55 53 53 53 50 50 50 4e 4e 4e 51 51 51 55 55 55 57 57 57 57 57 57 57 57 57 5c 5c 5c 5c 5c 5c 43 43 43 12 12 12 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 0d 0d 0d 4d 4d 4d 62 62 62 67 67 67 5a 5a 5a 4f 4f 4f 50 50 50 4f 4f 4f 4d 4d 4d 4a 4a 4a 49 49 49 4b 4b 4b 4b 4b 4b 49 49 49 4c 4c 4c 4f 4f 4f 54 54 54 55 55 55 59 59 59 56 56 56 42 42 42 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 5e 5e 5e 72 72 72 69 69 69 66 66 66 63 63 63 63 63 63 62 62 62 5c 5c 5c 53 53 53 4e 4e 4e 50 50 50 50 50 50 4e 4e 4e 4b 4b 4b 4b 4b 4b 4d 4d 4d 52 52 52 54 54 54 56 56 56 56 56 56 56 56 56 54 54 54 3b 3b 3b 08 08 08 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 31 31 31 5b 5b 5b 5e 5e 5e 4e 4e 4e 4b 4b 4b 4a 4a 4a 48 48 48 48 48 48 47 47 47 47 47 47 47 47 47 48 48 48 49 49 49 4b 4b 4b 4d 4d 4d 4f 4f 4f 52 52 52 56 56 56 50 50 50 3e 3e 3e 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 49 49 49 6b 6b 6b 63 63 63 5e 5e 5e 5c 5c 5c 5b 5b 5b 5c 5c 5c 60 60 60 50 50 50 4d 4d 4d 4d 4d 4d 4b 4b 4b 47 47 47 49 49 49 49 49 49 4c 4c 4c 51 51 51 54 54 54 57 57 57 56 56 56 53 53 53 54 54 54 30 30 30 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 21 21 21 50 50 50 4d 4d 4d 4a 4a 4a 49 49 49 4c 4c 4c 49 49 49 47 47 47 47 47 47 48 48 48 49 49 49 4d 4d 4d 4c 4c 4c 4c 4c 4c 4e 4e 4e 51 51 51 50 50 50 56 56 56 55 55 55 41 41 41 04 04 04 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 3c 3c 3c 5f 5f 5f 5d 5d 5d 5a 5a 5a 58 58 58 54 54 54 57 57 57 54 54 54 4d 4d 4d 4a 4a 4a 4b 4b 4b 4c 4c 4c 49 49 49 4c 4c 4c 49 49 49 4c 4c 4c 52 52 52 55 55 55 57 57 57 59 59 59 53 53 53 4f 4f 4f 1e 1e 1e 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 19 19 19 42 42 42 48 48 48 46 46 46 47 47 47 49 49 49 47 47 47 4d 4d 4d 49 49 49 49 49 49 48 48 48 49 49 49 4b 4b 4b 4e 4e 4e 50 50 50 51 51 51 51 51 51 54 54 54 5b 5b 5b 49 49 49 06 06 06 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 2f 2f 2f 52 52 52 55 55 55 56 56 56 54 54 54 52 52 52 52 52 52 51 51 51 4a 4a 4a 47 47 47 49 49 49 4b 4b 4b 4a 4a 4a 49 49 49 48 48 48 4e 4e 4e 52 52 52 57 57 57 59 59 59 52 52 52 4f 4f 4f 48 48 48 0f 0f 0f 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 3b 3b 3b 47 47 47 47 47 47 46 46 46 4a 4a 4a 45 45 45 4b 4b 4b 47 47 47 45 45 45 43 43 43 46 46 46 46 46 46 49 49 49 4b 4b 4b 4d 4d 4d 4a 4a 4a 4a 4a 4a 4b 4b 4b 46 46 46 08 08 08 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 24 24 24 4a 4a 4a 4e 4e 4e 51 51 51 52 52 52 52 52 52 4e 4e 4e 4a 4a 4a 4a 4a 4a 48 48 48 49 49 49 4b 4b 4b 48 48 48 49 49 49 49 49 49 4e 4e 4e 52 52 52 57 57 57 53 53 53 50 50 50 4b 4b 4b 39 39 39 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 31 31 31 46 46 46 46 46 46 43 43 43 45 45 45 44 44 44 3f 3f 3f 40 40 40 42 42 42 43 43 43 40 40 40 41 41 41 43 43 43 43 43 43 46 46 46 44 44 44 41 41 41 40 40 40 39 39 39 08 08 08 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 1e 1e 1e 45 45 45 4c 4c 4c 58 58 58 51 51 51 50 50 50 4a 4a 4a 48 48 48 46 46 46 47 47 47 4a 4a 4a 4a 4a 4a 49 49 49 49 49 49 4a 4a 4a 4e 4e 4e 51 51 51 51 51 51 4e 4e 4e 4a 4a 4a 46 46 46 1f 1f 1f 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 23 23 23 48 48 48 45 45 45 43 43 43 42 42 42 40 40 40 3d 3d 3d 3b 3b 3b 3e 3e 3e 3f 3f 3f 40 40 40 3e 3e 3e 3f 3f 3f 40 40 40 40 40 40 40 40 40 3c 3c 3c 3c 3c 3c 36 36 36 0a 0a 0a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 18 18 18 44 44 44 52 52 52 5b 5b 5b 50 50 50 4c 4c 4c 4a 4a 4a 4a 4a 4a 47 47 47 49 49 49 49 49 49 4b 4b 4b 49 49 49 4b 4b 4b 4c 4c 4c 4e 4e 4e 4f 4f 4f 4d 4d 4d 49 49 49 47 47 47 3a 3a 3a 0d 0d 0d 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 15 15 15 3f 3f 3f 45 45 45 42 42 42 44 44 44 3f 3f 3f 3d 3d 3d 3b 3b 3b 3d 3d 3d 3e 3e 3e 3c 3c 3c 3a 3a 3a 3c 3c 3c 3a 3a 3a 39 39 39 3a 3a 3a 38 38 38 3a 3a 3a 35 35 35 0e 0e 0e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 14 14 14 43 43 43 46 46 46 4a 4a 4a 4d 4d 4d 4d 4d 4d 4a 4a 4a 4a 4a 4a 47 47 47 49 49 49 4b 4b 4b 4b 4b 4b 4a 4a 4a 4b 4b 4b 4c 4c 4c 4c 4c 4c 4c 4c 4c 4a 4a 4a 47 47 47 47 47 47 2b 2b 2b 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 35 35 35 45 45 45 41 41 41 42 42 42 40 40 40 3e 3e 3e 3a 3a 3a 39 39 39 3a 3a 3a 39 39 39 39 39 39 3b 3b 3b 38 38 38 38 38 38 35 35 35 35 35 35 36 36 36 33 33 33 0f 0f 0f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 10 10 10 44 44 44 41 41 41 45 45 45 47 47 47 49 49 49 4a 4a 4a 48 48 48 4a 4a 4a 49 49 49 4b 4b 4b 4b 4b 4b 4c 4c 4c 4f 4f 4f 4b 4b 4b 4a 4a 4a 4a 4a 4a 4a 4a 4a 45 45 45 46 46 46 16 16 16 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 2a 2a 2a 44 44 44 42 42 42 45 45 45 41 41 41 3f 3f 3f 3c 3c 3c 38 38 38 38 38 38 37 37 37 38 38 38 3a 3a 3a 37 37 37 37 37 37 35 35 35 35 35 35 34 34 34 32 32 32 10 10 10 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 0b 0b 0b 3b 3b 3b 3c 3c 3c 3c 3c 3c 3f 3f 3f 41 41 41 44 44 44 48 48 48 4e 4e 4e 4b 4b 4b 49 49 49 4d 4d 4d 5e 5e 5e 57 57 57 51 51 51 55 55 55 4f 4f 4f 4b 4b 4b 48 48 48 35 35 35 07 07 07 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1b 1b 1b 3d 3d 3d 43 43 43 45 45 45 40 40 40 3e 3e 3e 3d 3d 3d 39 39 39 38 38 38 36 36 36 38 38 38 38 38 38 39 39 39 3a 3a 3a 38 38 38 39 39 39 34 34 34 32 32 32 15 15 15 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 08 08 08 37 37 37 3a 3a 3a 3e 3e 3e 41 41 41 44 44 44 46 46 46 46 46 46 4a 4a 4a 4b 4b 4b 4d 4d 4d 4f 4f 4f 58 58 58 47 47 47 47 47 47 46 46 46 51 51 51 4d 4d 4d 48 48 48 1c 1c 1c 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 31 31 31 42 42 42 44 44 44 43 43 43 3f 3f 3f 40 40 40 3d 3d 3d 39 39 39 36 36 36 36 36 36 38 38 38 37 37 37 3a 3a 3a 38 38 38 38 38 38 3c 3c 3c 38 38 38 17 17 17 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 05 05 05 34 34 34 3e 3e 3e 3f 3f 3f 46 46 46 46 46 46 4a 4a 4a 48 48 48 49 49 49 4c 4c 4c 4a 4a 4a 48 48 48 44 44 44 42 42 42 41 41 41 43 43 43 52 52 52 60 60 60 4d 4d 4d 09 09 09 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 20 20 20 3c 3c 3c 42 42 42 43 43 43 42 42 42 42 42 42 47 47 47 3d 3d 3d 35 35 35 34 34 34 38 38 38 39 39 39 39 39 39 39 39 39 3d 3d 3d 3b 3b 3b 30 30 30 16 16 16 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 32 32 32 36 36 36 38 38 38 3a 3a 3a 3d 3d 3d 3f 3f 3f 42 42 42 44 44 44 43 43 43 44 44 44 43 43 43 47 47 47 50 50 50 5e 5e 5e 6d 6d 6d 77 77 77 60 60 60 24 24 24 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 33 33 33 3c 3c 3c 41 41 41 44 44 44 45 45 45 51 51 51 52 52 52 43 43 43 3f 3f 3f 3c 3c 3c 36 36 36 37 37 37 3b 3b 3b 3a 3a 3a 32 32 32 2d 2d 2d 19 19 19 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 2a 2a 2a 31 31 31 34 34 34 35 35 35 39 39 39 3a 3a 3a 3e 3e 3e 48 48 48 54 54 54 5c 5c 5c 66 66 66 71 71 71 78 78 78 77 77 77 71 71 71 64 64 64 36 36 36 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1b 1b 1b 3c 3c 3c 3e 3e 3e 41 41 41 40 40 40 42 42 42 46 46 46 42 42 42 3e 3e 3e 3a 3a 3a 34 34 34 35 35 35 35 35 35 33 33 33 2e 2e 2e 2a 2a 2a 1b 1b 1b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 21 21 21 2d 2d 2d 2f 2f 2f 31 31 31 34 34 34 41 41 41 5e 5e 5e 72 72 72 78 78 78 78 78 78 74 74 74 6e 6e 6e 66 66 66 5e 5e 5e 55 55 55 3b 3b 3b 0a 0a 0a 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 2b 2b 2b 3c 3c 3c 3d 3d 3d 3e 3e 3e 3e 3e 3e 40 40 40 41 41 41 35 35 35 37 37 37 2e 2e 2e 2a 2a 2a 26 26 26 29 29 29 2c 2c 2c 29 29 29 1a 1a 1a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 18 18 18 27 27 27 27 27 27 2b 2b 2b 41 41 41 61 61 61 68 68 68 66 66 66 62 62 62 5f 5f 5f 5b 5b 5b 54 54 54 4f 4f 4f 49 49 49 35 35 35 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 2d 2d 2d 38 38 38 37 37 37 39 39 39 3f 3f 3f 3f 3f 3f 2d 2d 2d 2a 2a 2a 24 24 24 17 17 17 0a 0a 0a 16 16 16 16 16 16 13 13 13 0b 0b 0b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 06 06 06 09 09 09 0c 0c 0c 16 16 16 24 24 24 25 25 25 1f 1f 1f 20 20 20 1f 1f 1f 22 22 22 1f 1f 1f 1f 1f 1f 1e 1e 1e 15 15 15 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 1e 1e 1e 25 25 25 27 27 27 26 26 26 1e 1e 1e 0d 0d 0d 0b 0b 0b 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
