 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 05 05 05 07 07 07 0d 0d 0d 10 10 10 0d 0d 0d 0e 0e 0e 0c 0c 0c 0a 0a 0a 06 06 06 04 04 04 06 06 06 03 03 03 03 03 03 03 03 03 05 05 05 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 0a 0a 0a 0c 0c 0c 12 12 12 21 21 21 30 30 30 2b 2b 2b 37 37 37 42 42 42 39 39 39 2c 2c 2c 27 27 27 1f 1f 1f 1c 1c 1c 16 16 16 14 14 14 0f 0f 0f 0e 0e 0e 0b 0b 0b 07 07 07 07 07 07 07 07 07 05 05 05 05 05 05 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 06 06 06 05 05 05 0a 0a 0a 13 13 13 16 16 16 1f 1f 1f 2c 2c 2c 3b 3b 3b 48 48 48 4b 4b 4b 4d 4d 4d 57 57 57 5f 5f 5f 62 62 62 64 64 64 64 64 64 5c 5c 5c 52 52 52 4a 4a 4a 43 43 43 48 48 48 3e 3e 3e 41 41 41 45 45 45 3b 3b 3b 31 31 31 23 23 23 18 18 18 0d 0d 0d 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 0f 0f 0f 23 23 23 25 25 25 23 23 23 3a 3a 3a 48 48 48 56 56 56 64 64 64 67 67 67 6d 6d 6d 6e 6e 6e 6d 6d 6d 71 71 71 79 79 79 7a 7a 7a 7c 7c 7c 83 83 83 81 81 81 78 78 78 6e 6e 6e 68 68 68 5d 5d 5d 6b 6b 6b 72 72 72 8a 8a 8a a7 a7 a7 93 93 93 a8 a8 a8 bc bc bc 9b 9b 9b 6d 6d 6d 2a 2a 2a 10 10 10 06 06 06 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 18 18 18 2a 2a 2a 46 46 46 53 53 53 6f 6f 6f 76 76 76 75 75 75 7c 7c 7c 7f 7f 7f 77 77 77 79 79 79 78 78 78 76 76 76 7d 7d 7d 8a 8a 8a 98 98 98 99 99 99 a0 a0 a0 96 96 96 8f 8f 8f 85 85 85 7a 7a 7a 78 78 78 83 83 83 87 87 87 96 96 96 a8 a8 a8 c5 c5 c5 d0 d0 d0 cb cb cb ba ba ba 87 87 87 6f 6f 6f 52 52 52 31 31 31 14 14 14 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 19 19 19 2d 2d 2d 3c 3c 3c 49 49 49 5d 5d 5d 66 66 66 7a 7a 7a 94 94 94 93 93 93 92 92 92 98 98 98 9a 9a 9a ad ad ad b3 b3 b3 9c 9c 9c 8f 8f 8f 93 93 93 a4 a4 a4 9f 9f 9f 9c 9c 9c aa aa aa a2 a2 a2 9c 9c 9c a6 a6 a6 a1 a1 a1 a2 a2 a2 9f 9f 9f a6 a6 a6 c6 c6 c6 f9 f9 f9 f6 f6 f6 ef ef ef ce ce ce a2 a2 a2 8f 8f 8f 87 87 87 69 69 69 4e 4e 4e 34 34 34 0a 0a 0a 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 14 14 14 35 35 35 57 57 57 59 59 59 5e 5e 5e 6a 6a 6a 6d 6d 6d 85 85 85 98 98 98 a8 a8 a8 a7 a7 a7 b3 b3 b3 bf bf bf c7 c7 c7 d2 d2 d2 e6 e6 e6 ca ca ca c2 c2 c2 d9 d9 d9 e7 e7 e7 de de de c0 c0 c0 b8 b8 b8 b1 b1 b1 cb cb cb e7 e7 e7 e4 e4 e4 e4 e4 e4 d1 d1 d1 c7 c7 c7 ea ea ea fe fe fe f9 f9 f9 e9 e9 e9 e9 e9 e9 cd cd cd b3 b3 b3 ae ae ae 9f 9f 9f 82 82 82 90 90 90 48 48 48 0c 0c 0c 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 22 22 22 67 67 67 7b 7b 7b 6d 6d 6d 6b 6b 6b 79 79 79 97 97 97 a0 a0 a0 a5 a5 a5 a3 a3 a3 9e 9e 9e a2 a2 a2 b6 b6 b6 ce ce ce e1 e1 e1 eb eb eb f7 f7 f7 fc fc fc fe fe fe ff ff ff ff ff ff fe fe fe f5 f5 f5 dd dd dd e0 e0 e0 f3 f3 f3 fe fe fe fe fe fe ec ec ec d5 d5 d5 cd cd cd d2 d2 d2 f5 f5 f5 fc fc fc f2 f2 f2 df df df f0 f0 f0 d8 d8 d8 d7 d7 d7 c5 c5 c5 a2 a2 a2 a2 a2 a2 ae ae ae 3f 3f 3f 0f 0f 0f 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 10 10 10 44 44 44 76 76 76 7d 7d 7d 87 87 87 8a 8a 8a 91 91 91 9d 9d 9d 9e 9e 9e 9f 9f 9f 9a 9a 9a 92 92 92 9b 9b 9b b3 b3 b3 cd cd cd df df df e7 e7 e7 ee ee ee f9 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd fc fc fc fe fe fe ff ff ff fa fa fa e8 e8 e8 d7 d7 d7 c9 c9 c9 c7 c7 c7 d0 d0 d0 e7 e7 e7 f4 f4 f4 f1 f1 f1 f7 f7 f7 ef ef ef e8 e8 e8 f0 f0 f0 d6 d6 d6 ba ba ba bf bf bf af af af 3a 3a 3a 07 07 07 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 31 31 31 58 58 58 6b 6b 6b 84 84 84 92 92 92 96 96 96 96 96 96 9a 9a 9a 92 92 92 98 98 98 8e 8e 8e 91 91 91 9d 9d 9d b2 b2 b2 ce ce ce e3 e3 e3 e3 e3 e3 e1 e1 e1 ea ea ea fc fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f7 f7 ea ea ea da da da d2 d2 d2 d5 d5 d5 db db db d9 d9 d9 df df df e3 e3 e3 ec ec ec ed ed ed ee ee ee ef ef ef e0 e0 e0 c7 c7 c7 a2 a2 a2 9e 9e 9e 70 70 70 1b 1b 1b 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1c 1c 1c 5b 5b 5b 61 61 61 77 77 77 86 86 86 8d 8d 8d 87 87 87 8e 8e 8e 94 94 94 90 90 90 90 90 90 8c 8c 8c 94 94 94 a5 a5 a5 bf bf bf d6 d6 d6 ee ee ee e8 e8 e8 dc dc dc de de de f5 f5 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd fa fa fa f5 f5 f5 ea ea ea ea ea ea ea ea ea e9 e9 e9 e5 e5 e5 e7 e7 e7 eb eb eb ee ee ee e6 e6 e6 dc dc dc ce ce ce b6 b6 b6 a3 a3 a3 95 95 95 86 86 86 84 84 84 2c 2c 2c 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 49 49 49 7d 7d 7d 72 72 72 78 78 78 7d 7d 7d 7b 7b 7b 7a 7a 7a 81 81 81 94 94 94 ab ab ab ac ac ac a0 a0 a0 a5 a5 a5 bb bb bb d2 d2 d2 e4 e4 e4 ee ee ee ea ea ea de de de db db db ea ea ea fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fc fc fc fa fa fa fa fa fa f5 f5 f5 f1 f1 f1 e8 e8 e8 e4 e4 e4 e0 e0 e0 dd dd dd de de de dc dc dc d3 d3 d3 c5 c5 c5 b4 b4 b4 9f 9f 9f 92 92 92 87 87 87 7d 7d 7d 9e 9e 9e 49 49 49 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 26 26 26 7f 7f 7f 89 89 89 76 76 76 79 79 79 7b 7b 7b 7c 7c 7c 84 84 84 92 92 92 aa aa aa ca ca ca d6 d6 d6 cf cf cf ca ca ca cf cf cf da da da de de de e3 e3 e3 e2 e2 e2 dd dd dd da da da eb eb eb fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb f7 f7 f7 f5 f5 f5 ef ef ef eb eb eb e3 e3 e3 da da da d1 d1 d1 ce ce ce cb cb cb c8 c8 c8 c4 c4 c4 b5 b5 b5 a7 a7 a7 98 98 98 8d 8d 8d 7f 7f 7f 70 70 70 72 72 72 97 97 97 60 60 60 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 47 47 47 93 93 93 6c 6c 6c 70 70 70 74 74 74 75 75 75 7d 7d 7d 84 84 84 99 99 99 b3 b3 b3 c6 c6 c6 d1 d1 d1 cd cd cd c8 c8 c8 cd cd cd d8 d8 d8 de de de de de de dc dc dc dc dc dc dd dd dd f4 f4 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fd fd fd fe fe fe fd fd fd fa fa fa f1 f1 f1 dc dc dc c9 c9 c9 c6 c6 c6 c5 c5 c5 c2 c2 c2 bd bd bd b6 b6 b6 a7 a7 a7 99 99 99 8f 8f 8f 83 83 83 73 73 73 6e 6e 6e 6a 6a 6a 7b 7b 7b 5c 5c 5c 07 07 07 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 64 64 64 88 88 88 69 69 69 68 68 68 6d 6d 6d 72 72 72 77 77 77 7b 7b 7b 88 88 88 a1 a1 a1 b5 b5 b5 bb bb bb b9 b9 b9 b7 b7 b7 c0 c0 c0 d4 d4 d4 d1 d1 d1 d5 d5 d5 dd dd dd e6 e6 e6 f1 f1 f1 fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb e7 e7 e7 e7 e7 e7 e8 e8 e8 df df df d5 d5 d5 cd cd cd c4 c4 c4 b9 b9 b9 b9 b9 b9 ba ba ba b8 b8 b8 bc bc bc b3 b3 b3 a8 a8 a8 9e 9e 9e 91 91 91 7e 7e 7e 7a 7a 7a 73 73 73 6a 6a 6a 73 73 73 52 52 52 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 5f 5f 5f 7d 7d 7d 6f 6f 6f 69 69 69 6b 6b 6b 74 74 74 79 79 79 7e 7e 7e 88 88 88 9c 9c 9c ae ae ae b2 b2 b2 b1 b1 b1 b0 b0 b0 b0 b0 b0 bf bf bf c2 c2 c2 be be be c2 c2 c2 dc dc dc f9 f9 f9 ec ec ec de de de da da da f5 f5 f5 fe fe fe fb fb fb dc dc dc bb bb bb b8 b8 b8 b2 b2 b2 b3 b3 b3 b2 b2 b2 b0 b0 b0 ad ad ad aa aa aa ad ad ad ad ad ad b1 b1 b1 b1 b1 b1 a6 a6 a6 9d 9d 9d 90 90 90 83 83 83 7c 7c 7c 70 70 70 6d 6d 6d 6a 6a 6a 3b 3b 3b 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 59 59 59 77 77 77 7b 7b 7b 78 78 78 73 73 73 7d 7d 7d 86 86 86 8b 8b 8b 92 92 92 a2 a2 a2 aa aa aa ad ad ad ac ac ac aa aa aa a8 a8 a8 b2 b2 b2 ae ae ae a8 a8 a8 ac ac ac c9 c9 c9 c3 c3 c3 8f 8f 8f 7a 7a 7a 75 75 75 9b 9b 9b d2 d2 d2 fc fc fc df df df ae ae ae 9f 9f 9f a9 a9 a9 ad ad ad a7 a7 a7 a2 a2 a2 a2 a2 a2 a1 a1 a1 a1 a1 a1 a2 a2 a2 a4 a4 a4 a3 a3 a3 99 99 99 92 92 92 87 87 87 7f 7f 7f 78 78 78 76 76 76 6f 6f 6f 63 63 63 34 34 34 05 05 05 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0f 0f 0f 62 62 62 78 78 78 7f 7f 7f 8a 8a 8a 86 86 86 8c 8c 8c 94 94 94 9a 9a 9a a0 a0 a0 a4 a4 a4 a9 a9 a9 ab ab ab a8 a8 a8 a8 a8 a8 aa aa aa b7 b7 b7 a8 a8 a8 a6 a6 a6 ab ab ab bc bc bc 71 71 71 52 52 52 41 41 41 49 49 49 6b 6b 6b 81 81 81 d5 d5 d5 ea ea ea b3 b3 b3 97 97 97 a7 a7 a7 aa aa aa a2 a2 a2 9a 9a 9a 9a 9a 9a 97 97 97 96 96 96 97 97 97 97 97 97 93 93 93 8a 8a 8a 87 87 87 82 82 82 7b 7b 7b 7b 7b 7b 77 77 77 6e 6e 6e 69 69 69 49 49 49 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 1d 1d 1d 75 75 75 7f 7f 7f 81 81 81 91 91 91 93 93 93 97 97 97 9f 9f 9f a3 a3 a3 a7 a7 a7 a8 a8 a8 ab ab ab ab ab ab a6 a6 a6 ad ad ad b1 b1 b1 b1 b1 b1 af af af ad ad ad b3 b3 b3 9d 9d 9d 3a 3a 3a 24 24 24 1f 1f 1f 23 23 23 30 30 30 58 58 58 c9 c9 c9 e1 e1 e1 a5 a5 a5 96 96 96 a7 a7 a7 a3 a3 a3 9a 9a 9a 96 96 96 91 91 91 90 90 90 8e 8e 8e 8a 8a 8a 89 89 89 85 85 85 80 80 80 7e 7e 7e 7c 7c 7c 7b 7b 7b 79 79 79 71 71 71 6d 6d 6d 70 70 70 5a 5a 5a 16 16 16 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 06 06 06 2d 2d 2d 85 85 85 81 81 81 86 86 86 8c 8c 8c 90 90 90 9a 9a 9a a0 a0 a0 a3 a3 a3 a5 a5 a5 a7 a7 a7 a8 a8 a8 ac ac ac aa aa aa b0 b0 b0 b3 b3 b3 b6 b6 b6 b3 b3 b3 b3 b3 b3 c2 c2 c2 85 85 85 17 17 17 0f 0f 0f 0a 0a 0a 0c 0c 0c 16 16 16 34 34 34 a5 a5 a5 ab ab ab 98 98 98 98 98 98 9f 9f 9f 9d 9d 9d 95 95 95 8e 8e 8e 88 88 88 87 87 87 85 85 85 81 81 81 7b 7b 7b 77 77 77 75 75 75 74 74 74 79 79 79 77 77 77 6f 6f 6f 6a 6a 6a 70 70 70 69 69 69 67 67 67 2d 2d 2d 05 05 05 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 09 09 09 3b 3b 3b 91 91 91 7b 7b 7b 83 83 83 8a 8a 8a 89 89 89 92 92 92 98 98 98 9c 9c 9c 9f 9f 9f a0 a0 a0 a3 a3 a3 a3 a3 a3 ab ab ab b6 b6 b6 b9 b9 b9 b6 b6 b6 b4 b4 b4 bc bc bc c8 c8 c8 84 84 84 0a 0a 0a 06 06 06 04 04 04 03 03 03 08 08 08 1d 1d 1d 7d 7d 7d 95 95 95 98 98 98 95 95 95 96 96 96 98 98 98 90 90 90 89 89 89 83 83 83 7f 7f 7f 7d 7d 7d 77 77 77 71 71 71 6d 6d 6d 6b 6b 6b 70 70 70 70 70 70 69 69 69 6b 6b 6b 6d 6d 6d 6b 6b 6b 61 61 61 70 70 70 3f 3f 3f 09 09 09 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0a 0a 0a 44 44 44 93 93 93 76 76 76 7d 7d 7d 89 89 89 88 88 88 8d 8d 8d 91 91 91 92 92 92 93 93 93 96 96 96 99 99 99 9f 9f 9f ac ac ac b6 b6 b6 b3 b3 b3 b0 b0 b0 ac ac ac b7 b7 b7 bf bf bf 84 84 84 06 06 06 04 04 04 03 03 03 03 03 03 06 06 06 11 11 11 7b 7b 7b 8e 8e 8e 89 89 89 8b 8b 8b 8b 8b 8b 8e 8e 8e 8b 8b 8b 83 83 83 7e 7e 7e 79 79 79 76 76 76 6f 6f 6f 6b 6b 6b 68 68 68 67 67 67 6c 6c 6c 63 63 63 65 65 65 6d 6d 6d 65 65 65 59 59 59 57 57 57 72 72 72 4a 4a 4a 0c 0c 0c 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0d 0d 0d 4b 4b 4b 95 95 95 76 76 76 72 72 72 7f 7f 7f 85 85 85 88 88 88 87 87 87 88 88 88 8a 8a 8a 8c 8c 8c 92 92 92 99 99 99 a1 a1 a1 ab ab ab a7 a7 a7 a1 a1 a1 9a 9a 9a 9f 9f 9f a2 a2 a2 80 80 80 05 05 05 04 04 04 03 03 03 03 03 03 04 04 04 0a 0a 0a 71 71 71 80 80 80 81 81 81 82 82 82 85 85 85 87 87 87 85 85 85 81 81 81 7a 7a 7a 76 76 76 72 72 72 6b 6b 6b 66 66 66 65 65 65 67 67 67 61 61 61 62 62 62 67 67 67 62 62 62 5d 5d 5d 53 53 53 50 50 50 70 70 70 52 52 52 11 11 11 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0e 0e 0e 4e 4e 4e 92 92 92 76 76 76 6b 6b 6b 70 70 70 7b 7b 7b 84 84 84 83 83 83 80 80 80 82 82 82 84 84 84 86 86 86 8d 8d 8d 92 92 92 9c 9c 9c 9d 9d 9d 96 96 96 8c 8c 8c 8b 8b 8b 89 89 89 78 78 78 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 63 63 63 78 78 78 79 79 79 7b 7b 7b 7e 7e 7e 7f 7f 7f 7e 7e 7e 7c 7c 7c 76 76 76 6d 6d 6d 6a 6a 6a 66 66 66 61 61 61 63 63 63 60 60 60 5c 5c 5c 63 63 63 64 64 64 5b 5b 5b 58 58 58 50 50 50 4a 4a 4a 6c 6c 6c 53 53 53 11 11 11 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0e 0e 0e 4f 4f 4f 87 87 87 65 65 65 66 66 66 67 67 67 6c 6c 6c 84 84 84 8b 8b 8b 84 84 84 83 83 83 83 83 83 88 88 88 8a 8a 8a 8d 8d 8d 95 95 95 95 95 95 8f 8f 8f 8a 8a 8a 86 86 86 83 83 83 72 72 72 08 08 08 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 57 57 57 73 73 73 73 73 73 76 76 76 75 75 75 77 77 77 76 76 76 72 72 72 6d 6d 6d 68 68 68 64 64 64 60 60 60 5e 5e 5e 5d 5d 5d 57 57 57 5a 5a 5a 65 65 65 62 62 62 59 59 59 59 59 59 51 51 51 44 44 44 5a 5a 5a 56 56 56 14 14 14 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0b 0b 0b 4f 4f 4f 7f 7f 7f 58 58 58 5a 5a 5a 68 68 68 65 65 65 6a 6a 6a 79 79 79 84 84 84 86 86 86 86 86 86 8a 8a 8a 8f 8f 8f 91 91 91 8e 8e 8e 8e 8e 8e 8c 8c 8c 8c 8c 8c 8f 8f 8f 8c 8c 8c 7e 7e 7e 0b 0b 0b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 56 56 56 84 84 84 7b 7b 7b 7d 7d 7d 7b 7b 7b 7b 7b 7b 72 72 72 6d 6d 6d 66 66 66 62 62 62 5f 5f 5f 5d 5d 5d 56 56 56 54 54 54 5d 5d 5d 69 69 69 70 70 70 62 62 62 5b 5b 5b 66 66 66 50 50 50 45 45 45 4c 4c 4c 52 52 52 12 12 12 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 06 06 06 43 43 43 7a 7a 7a 54 54 54 53 53 53 58 58 58 63 63 63 67 67 67 67 67 67 69 69 69 6d 6d 6d 72 72 72 74 74 74 74 74 74 6f 6f 6f 6f 6f 6f 6d 6d 6d 6d 6d 6d 6a 6a 6a 6c 6c 6c 6a 6a 6a 63 63 63 0d 0d 0d 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 44 44 44 7a 7a 7a 77 77 77 7b 7b 7b 7d 7d 7d 77 77 77 68 68 68 64 64 64 61 61 61 5e 5e 5e 5a 5a 5a 55 55 55 53 53 53 58 58 58 5d 5d 5d 63 63 63 63 63 63 57 57 57 5c 5c 5c 5d 5d 5d 4d 4d 4d 44 44 44 45 45 45 4b 4b 4b 09 09 09 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 2b 2b 2b 78 78 78 55 55 55 51 51 51 52 52 52 53 53 53 5c 5c 5c 63 63 63 61 61 61 60 60 60 60 60 60 5d 5d 5d 5c 5c 5c 59 59 59 5a 5a 5a 59 59 59 59 59 59 5b 5b 5b 5a 5a 5a 59 59 59 53 53 53 0e 0e 0e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 2e 2e 2e 63 63 63 60 60 60 62 62 62 62 62 62 62 62 62 61 61 61 5e 5e 5e 5c 5c 5c 5b 5b 5b 58 58 58 53 53 53 5b 5b 5b 5c 5c 5c 60 60 60 63 63 63 60 60 60 5c 5c 5c 5d 5d 5d 52 52 52 4a 4a 4a 46 46 46 40 40 40 2b 2b 2b 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 65 65 65 56 56 56 4d 4d 4d 4c 4c 4c 4f 4f 4f 4f 4f 4f 51 51 51 51 51 51 50 50 50 52 52 52 52 52 52 4f 4f 4f 4e 4e 4e 52 52 52 53 53 53 54 54 54 54 54 54 52 52 52 51 51 51 4d 4d 4d 10 10 10 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 25 25 25 5b 5b 5b 5d 5d 5d 5d 5d 5d 60 60 60 60 60 60 5d 5d 5d 5b 5b 5b 59 59 59 57 57 57 56 56 56 57 57 57 5f 5f 5f 57 57 57 57 57 57 62 62 62 71 71 71 67 67 67 61 61 61 5e 5e 5e 4f 4f 4f 49 49 49 39 39 39 12 12 12 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 3d 3d 3d 55 55 55 49 49 49 49 49 49 4a 4a 4a 4c 4c 4c 4a 4a 4a 48 48 48 45 45 45 45 45 45 47 47 47 46 46 46 44 44 44 46 46 46 4c 4c 4c 51 51 51 4b 4b 4b 49 49 49 49 49 49 46 46 46 12 12 12 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 1f 1f 1f 54 54 54 56 56 56 5a 5a 5a 62 62 62 6b 6b 6b 5d 5d 5d 56 56 56 56 56 56 58 58 58 5d 5d 5d 5c 5c 5c 56 56 56 50 50 50 4d 4d 4d 67 67 67 8f 8f 8f 85 85 85 6b 6b 6b 5f 5f 5f 4f 4f 4f 47 47 47 2d 2d 2d 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 29 29 29 4f 4f 4f 49 49 49 47 47 47 47 47 47 47 47 47 45 45 45 46 46 46 44 44 44 44 44 44 44 44 44 45 45 45 43 43 43 43 43 43 41 41 41 43 43 43 47 47 47 47 47 47 45 45 45 46 46 46 15 15 15 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 17 17 17 50 50 50 4f 4f 4f 53 53 53 59 59 59 5e 5e 5e 5a 5a 5a 56 56 56 53 53 53 53 53 53 53 53 53 53 53 53 4e 4e 4e 4c 4c 4c 4c 4c 4c 58 58 58 77 77 77 7d 7d 7d 64 64 64 5a 5a 5a 4d 4d 4d 46 46 46 1b 1b 1b 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 1f 1f 1f 4a 4a 4a 46 46 46 44 44 44 43 43 43 46 46 46 45 45 45 44 44 44 44 44 44 43 43 43 42 42 42 45 45 45 43 43 43 40 40 40 3d 3d 3d 3c 3c 3c 3b 3b 3b 3e 3e 3e 3f 3f 3f 3c 3c 3c 13 13 13 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 11 11 11 4d 4d 4d 4e 4e 4e 4f 4f 4f 52 52 52 51 51 51 57 57 57 58 58 58 53 53 53 4f 4f 4f 4e 4e 4e 4d 4d 4d 4b 4b 4b 4c 4c 4c 4b 4b 4b 4f 4f 4f 53 53 53 5c 5c 5c 59 59 59 53 53 53 4b 4b 4b 38 38 38 0d 0d 0d 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 17 17 17 43 43 43 46 46 46 41 41 41 41 41 41 43 43 43 43 43 43 42 42 42 43 43 43 42 42 42 42 42 42 42 42 42 41 41 41 41 41 41 3d 3d 3d 3b 3b 3b 39 39 39 3b 3b 3b 39 39 39 36 36 36 12 12 12 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 0c 0c 0c 4d 4d 4d 57 57 57 54 54 54 55 55 55 53 53 53 54 54 54 4c 4c 4c 4c 4c 4c 46 46 46 47 47 47 48 48 48 49 49 49 49 49 49 4a 4a 4a 4c 4c 4c 4d 4d 4d 52 52 52 58 58 58 4d 4d 4d 45 45 45 2a 2a 2a 06 06 06 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 11 11 11 37 37 37 46 46 46 44 44 44 41 41 41 45 45 45 43 43 43 43 43 43 42 42 42 42 42 42 41 41 41 44 44 44 42 42 42 40 40 40 3d 3d 3d 3a 3a 3a 39 39 39 3b 3b 3b 38 38 38 35 35 35 14 14 14 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 08 08 08 49 49 49 4a 4a 4a 46 46 46 45 45 45 48 48 48 48 48 48 46 46 46 45 45 45 44 44 44 46 46 46 48 48 48 47 47 47 49 49 49 49 49 49 4b 4b 4b 4c 4c 4c 51 51 51 51 51 51 4f 4f 4f 3f 3f 3f 1e 1e 1e 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 2f 2f 2f 44 44 44 46 46 46 3f 3f 3f 42 42 42 41 41 41 40 40 40 42 42 42 43 43 43 44 44 44 42 42 42 41 41 41 41 41 41 3d 3d 3d 3b 3b 3b 39 39 39 38 38 38 37 37 37 33 33 33 16 16 16 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 06 06 06 3a 3a 3a 42 42 42 42 42 42 41 41 41 42 42 42 3f 3f 3f 40 40 40 40 40 40 42 42 42 47 47 47 47 47 47 47 47 47 48 48 48 48 48 48 4a 4a 4a 4b 4b 4b 4f 4f 4f 4f 4f 4f 4a 4a 4a 39 39 39 0d 0d 0d 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 1e 1e 1e 42 42 42 49 49 49 40 40 40 41 41 41 41 41 41 41 41 41 40 40 40 43 43 43 43 43 43 44 44 44 41 41 41 40 40 40 3f 3f 3f 3d 3d 3d 3b 3b 3b 37 37 37 37 37 37 32 32 32 18 18 18 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 36 36 36 3e 3e 3e 3f 3f 3f 40 40 40 3e 3e 3e 40 40 40 41 41 41 40 40 40 45 45 45 47 47 47 48 48 48 47 47 47 49 49 49 47 47 47 48 48 48 49 49 49 4a 4a 4a 49 49 49 45 45 45 2a 2a 2a 05 05 05 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 11 11 11 35 35 35 46 46 46 41 41 41 46 46 46 45 45 45 4a 4a 4a 44 44 44 46 46 46 44 44 44 42 42 42 3e 3e 3e 3f 3f 3f 3d 3d 3d 3b 3b 3b 39 39 39 36 36 36 35 35 35 31 31 31 1a 1a 1a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 31 31 31 39 39 39 3d 3d 3d 3f 3f 3f 40 40 40 40 40 40 41 41 41 40 40 40 46 46 46 47 47 47 48 48 48 46 46 46 46 46 46 44 44 44 44 44 44 45 45 45 49 49 49 48 48 48 42 42 42 18 18 18 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 29 29 29 41 41 41 40 40 40 42 42 42 41 41 41 46 46 46 3e 3e 3e 41 41 41 42 42 42 40 40 40 3f 3f 3f 3f 3f 3f 3c 3c 3c 3b 3b 3b 38 38 38 36 36 36 34 34 34 2f 2f 2f 1a 1a 1a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 2c 2c 2c 38 38 38 3c 3c 3c 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 41 41 41 42 42 42 44 44 44 44 44 44 43 43 43 44 44 44 40 40 40 41 41 41 43 43 43 46 46 46 45 45 45 39 39 39 08 08 08 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 1d 1d 1d 37 37 37 40 40 40 46 46 46 41 41 41 3f 3f 3f 3e 3e 3e 3e 3e 3e 40 40 40 3f 3f 3f 3f 3f 3f 3f 3f 3f 3a 3a 3a 3a 3a 3a 37 37 37 38 38 38 34 34 34 30 30 30 1a 1a 1a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 26 26 26 36 36 36 38 38 38 39 39 39 39 39 39 39 39 39 38 38 38 3e 3e 3e 3e 3e 3e 3e 3e 3e 42 42 42 41 41 41 3f 3f 3f 3c 3c 3c 3e 3e 3e 41 41 41 45 45 45 44 44 44 23 23 23 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 11 11 11 2a 2a 2a 3b 3b 3b 43 43 43 40 40 40 40 40 40 3a 3a 3a 3d 3d 3d 40 40 40 3f 3f 3f 41 41 41 40 40 40 3e 3e 3e 3b 3b 3b 38 38 38 38 38 38 35 35 35 32 32 32 1e 1e 1e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 25 25 25 37 37 37 37 37 37 36 36 36 37 37 37 38 38 38 36 36 36 3b 3b 3b 3c 3c 3c 3d 3d 3d 3e 3e 3e 3f 3f 3f 3d 3d 3d 3b 3b 3b 3a 3a 3a 3f 3f 3f 43 43 43 3a 3a 3a 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 22 22 22 34 34 34 3e 3e 3e 40 40 40 43 43 43 3a 3a 3a 3d 3d 3d 3e 3e 3e 3f 3f 3f 40 40 40 42 42 42 3e 3e 3e 3b 3b 3b 39 39 39 35 35 35 34 34 34 33 33 33 22 22 22 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 21 21 21 35 35 35 35 35 35 35 35 35 34 34 34 35 35 35 35 35 35 37 37 37 38 38 38 3a 3a 3a 3b 3b 3b 3a 3a 3a 3c 3c 3c 3a 3a 3a 39 39 39 3e 3e 3e 42 42 42 24 24 24 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 13 13 13 2a 2a 2a 3a 3a 3a 3e 3e 3e 3e 3e 3e 3c 3c 3c 3b 3b 3b 3b 3b 3b 3d 3d 3d 3e 3e 3e 48 48 48 49 49 49 42 42 42 44 44 44 37 37 37 31 31 31 31 31 31 26 26 26 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 1b 1b 1b 33 33 33 34 34 34 32 32 32 32 32 32 32 32 32 35 35 35 38 38 38 38 38 38 3b 3b 3b 3a 3a 3a 3a 3a 3a 3d 3d 3d 41 41 41 42 42 42 41 41 41 34 34 34 0c 0c 0c 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 1f 1f 1f 31 31 31 3e 3e 3e 3d 3d 3d 3c 3c 3c 3b 3b 3b 38 38 38 3f 3f 3f 3f 3f 3f 4a 4a 4a 52 52 52 51 51 51 55 55 55 3b 3b 3b 32 32 32 2f 2f 2f 26 26 26 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 18 18 18 31 31 31 32 32 32 32 32 32 32 32 32 31 31 31 31 31 31 34 34 34 36 36 36 37 37 37 3a 3a 3a 45 45 45 60 60 60 70 70 70 6c 6c 6c 46 46 46 19 19 19 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0e 0e 0e 28 28 28 3a 3a 3a 48 48 48 3f 3f 3f 3c 3c 3c 38 38 38 39 39 39 3c 3c 3c 4f 4f 4f 5b 5b 5b 5a 5a 5a 5c 5c 5c 3b 3b 3b 31 31 31 2c 2c 2c 26 26 26 05 05 05 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 14 14 14 31 31 31 2f 2f 2f 2f 2f 2f 2e 2e 2e 2f 2f 2f 32 32 32 34 34 34 36 36 36 3e 3e 3e 5a 5a 5a 71 71 71 75 75 75 72 72 72 65 65 65 2c 2c 2c 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 17 17 17 2e 2e 2e 4b 4b 4b 4d 4d 4d 3e 3e 3e 3b 3b 3b 38 38 38 3b 3b 3b 4f 4f 4f 56 56 56 55 55 55 4f 4f 4f 30 30 30 2d 2d 2d 29 29 29 24 24 24 05 05 05 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 0e 0e 0e 2a 2a 2a 27 27 27 27 27 27 28 28 28 2a 2a 2a 2a 2a 2a 2f 2f 2f 42 42 42 5d 5d 5d 67 67 67 62 62 62 5f 5f 5f 5a 5a 5a 34 34 34 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 1b 1b 1b 30 30 30 41 41 41 3a 3a 3a 38 38 38 34 34 34 31 31 31 3b 3b 3b 3d 3d 3d 3b 3b 3b 24 24 24 1b 1b 1b 19 19 19 15 15 15 0f 0f 0f 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 05 05 05 09 09 09 0b 0b 0b 0a 0a 0a 0b 0b 0b 0c 0c 0c 0e 0e 0e 1a 1a 1a 22 22 22 25 25 25 21 21 21 22 22 22 22 22 22 16 16 16 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 13 13 13 20 20 20 22 22 22 1a 1a 1a 13 13 13 0b 0b 0b 0f 0f 0f 10 10 10 13 13 13 06 06 06 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
