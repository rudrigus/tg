-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- ***************************************************************************
-- This file contains a Vhdl test bench template that is freely editable to   
-- suit user's needs .Comments are provided in each section to help the user  
-- fill out necessary details.                                                
-- ***************************************************************************
-- Generated on "11/18/2015 21:55:21"
                                                            
-- Vhdl Test Bench template for design  :  ProcessadorImagemGMAW
-- 
-- Simulation tool : ModelSim-Altera (VHDL)
-- 

LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;

ENTITY ProcessadorImagemGMAW_TB IS
END ProcessadorImagemGMAW_TB;
ARCHITECTURE ProcessadorImagemGMAW_arch OF ProcessadorImagemGMAW_TB IS
-- constants                                                 

constant imagem_padrao0 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

constant imagem_padrao1 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

constant imagem_padrao2 : MatrizImagem := ((X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"49", X"49", X"49", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"9B", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"49", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"5B", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"A4", X"F7", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"52", X"5B", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"52", X"52", X"52", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"9B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"52", X"52", X"5B", X"5B", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"52", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"5B", X"A4", X"9B", X"9B", X"5B", X"5B", X"52", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"5B", X"A4", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"52", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"52", X"52", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"52", X"5B", X"52", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"52", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"5B", X"5B", X"9B", X"5B", X"5B", X"5B", X"5B", X"9B", X"5B", X"9B", X"5B", X"5B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"A4", X"9B", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"5B", X"5B", X"5B", X"5B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"5B", X"5B", X"9B", X"9B", X"5B", X"9B", X"5B", X"A4", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"A4", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"9B", X"9B", X"9B", X"5B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"9B", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"9B", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"9B", X"9B", X"9B", X"A4", X"9B", X"9B", X"9B", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"9B", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00", X"00", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"5B", X"00", X"00", X"00", X"00", X"00", X"00", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"08", X"08", X"08", X"08", X"07", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"07", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"A4", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"07", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"5B", X"49", X"00", X"00", X"00", X"49", X"49", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"9B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"9B", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"F6", X"F6", X"FF", X"F7", X"52", X"49", X"49", X"49", X"52", X"52", X"08", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"9B", X"5B", X"52", X"52", X"5B", X"F7", X"F6", X"07", X"08", X"07", X"07", X"07", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"F7", X"5B", X"9B", X"A4", X"F7", X"F7", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"07", X"07", X"FF", X"07", X"FF", X"FF", X"08", X"08", X"08", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"A4", X"F7", X"A4", X"A4", X"5B", X"F7", X"5B", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"49", X"A4", X"5B", X"9B", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"08", X"F6", X"F6", X"F6", X"08", X"08", X"08", X"07", X"07", X"07", X"F7", X"F7", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"52", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"9B", X"F7", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"F6", X"F6", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"F7", X"A4", X"A4", X"A4", X"9B", X"A4", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"07", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"F7", X"A4", X"A4", X"F7", X"F7", X"07", X"07", X"08", X"08", X"F6", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"9B", X"9B", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"08", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"F7", X"49", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"F7", X"A4", X"9B", X"A4", X"F7", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"FF", X"F6", X"F6", X"F6", X"08", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"FF", X"F6", X"08", X"08", X"07", X"07", X"F7", X"A4", X"A4", X"A4", X"A4", X"A4", X"9B", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"A4", X"5B", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"F6", X"07", X"07", X"07", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"9B", X"A4", X"52", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"5B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"F6", X"08", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"A4", X"5B", X"9B", X"9B", X"9B", X"49", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"9B", X"5B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"F6", X"08", X"07", X"08", X"07", X"F7", X"F7", X"F7", X"A4", X"9B", X"9B", X"9B", X"9B", X"5B", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"9B", X"9B", X"A4", X"A4", X"F7", X"07", X"07", X"08", X"F6", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"F6", X"07", X"07", X"F7", X"07", X"07", X"F7", X"F7", X"A4", X"A4", X"A4", X"9B", X"9B", X"5B", X"52", X"9B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"A4", X"A4", X"9B", X"9B", X"A4", X"F7", X"F7", X"07", X"07", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"FF", X"08", X"07", X"F7", X"F7", X"A4", X"A4", X"F7", X"A4", X"A4", X"A4", X"5B", X"5B", X"5B", X"5B", X"5B", X"52", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"52", X"5B", X"A4", X"A4", X"A4", X"A4", X"F7", X"07", X"F6", X"FF", X"FF", X"F6", X"07", X"F7", X"F7", X"A4", X"9B", X"A4", X"A4", X"9B", X"9B", X"5B", X"5B", X"5B", X"5B", X"52", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"52", X"9B", X"A4", X"F7", X"07", X"F7", X"07", X"07", X"07", X"F7", X"A4", X"A4", X"F7", X"F7", X"F7", X"A4", X"5B", X"52", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"),
(X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"49", X"49", X"52", X"52", X"52", X"5B", X"5B", X"52", X"52", X"49", X"52", X"00", X"49", X"49", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00"));

-- signals                                                   
SIGNAL ENDSIM : STD_LOGIC := '0';
SIGNAL clk_count : natural := 0;
SIGNAL brilho_maximo : UNSIGNED(24 DOWNTO 0);
SIGNAL in_clock : STD_LOGIC;
SIGNAL in_janela : STD_LOGIC;
SIGNAL pixel_entrada : STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL bloco_atual : unsigned(1 downto 0) := "00";
SIGNAL linha : integer range 0 to numcols - 1 := 0;
SIGNAL coluna : integer range 0 to numlin - 1 := 0;
SIGNAL reset : STD_LOGIC;
SIGNAL start_stop :  STD_LOGIC;
SIGNAL contador12b : STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL qtd_imagens : UNSIGNED(1 DOWNTO 0) := "11";
--SIGNAL fim_imagem : STD_LOGIC := '0';
SIGNAL frequencia_camera : real := 150.000E6;

COMPONENT ProcessadorImagemGMAW
	PORT (
	brilho_maximo : IN UNSIGNED(24 DOWNTO 0);
	in_clock : IN STD_LOGIC;
	in_janela : IN STD_LOGIC;
	pixel_entrada : IN STD_LOGIC_VECTOR(7 DOWNTO 0)
	);	
END COMPONENT;


-- Procedure for clock generation
  procedure clk_gen(signal clk : out std_logic; constant FREQ : real) is
    constant PERIOD    : time := 1 sec / FREQ;        -- Full period
    constant HIGH_TIME : time := PERIOD / 2;          -- High time
    constant LOW_TIME  : time := PERIOD - HIGH_TIME;  -- Low time; always >= HIGH_TIME
  begin
    -- Check the arguments
    assert (HIGH_TIME /= 0 fs) report "clk_plain: High time is zero; time resolution to large for frequency" severity FAILURE;
    -- Generate a clock cycle
    loop
      if (ENDSIM = '0') then
        clk <= '1';
        wait for HIGH_TIME;
        clk <= '0';
        wait for LOW_TIME;
      else
        wait;
      end if;
    end loop;
  end procedure;



BEGIN
  -- Clock generation with concurrent procedure call
  clk_gen(in_clock, frequencia_camera);  -- 166.667 MHz clock

  -- Time resolution show
  assert FALSE report "Time resolution: " & time'image(time'succ(0 fs)) severity NOTE;



	i1 : ProcessadorImagemGMAW
	PORT MAP (
-- list connections between master ports and signals
	brilho_maximo => brilho_maximo,
	in_clock => in_clock,
	in_janela => in_janela,
	pixel_entrada => pixel_entrada
	);

brilho_maximo <= to_unsigned(720000,25) after 0 ns;
in_janela <= '1' after 0 ns,
             '0' after 5 ns;

IN_process: process (in_clock) begin
  if(rising_edge(in_clock)) then
    clk_count <= clk_count + 1;

    -- avanca as imagens
    case bloco_atual is
      when "00" => pixel_entrada <= STD_LOGIC_VECTOR(imagem_padrao0(linha, coluna));
      when "01" => pixel_entrada <= STD_LOGIC_VECTOR(imagem_padrao1(linha, coluna));
      when "10" => pixel_entrada <= STD_LOGIC_VECTOR(imagem_padrao2(linha, coluna));
      when others => pixel_entrada <= STD_LOGIC_VECTOR(imagem_padrao0(linha, coluna));
    end case;

    -- marcacao de linhas, colunas e parada na simulacao
    if (coluna = numcols - 1) then
      coluna <= 0;
      if (linha = numlin -1) then
        linha <= 0;
        --fim_imagem <= '1';
        bloco_atual <= bloco_atual + 1;
      else
        linha <= linha + 1;
      end if;    
    else
      coluna <= coluna + 1;
    end if;

    if (clk_count = 3 * (numlin * numcols)) then
      ENDSIM <= '1';
    end if;
  end if;
  

--when -label end_of_simulation {end_of_sim == '1'} {echo "End of simulation" ; stop ;}
end process;


END ProcessadorImagemGMAW_arch;
 