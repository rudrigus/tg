 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 05 05 06 05 06 00 06 05 03 0b 11 12 17 18 0f 10 12 1d 1e 0d 25 2b 35 2f 24 20 2a 2b 37 39 2d 38 43 4a 44 4d 4d 51 55 4b 4a 45 44 49 59 6a 56 43 3c 45 52 4b 42 27 1e 1f 1a 1d 26 2a 38 37 2b 2b 24 2b 1a 24 29 20 18 1d 20 26 1d 0f 18 14 11 15 09 09 12 15 12 02 06 05 04 00 06 06 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 05 06 05 03 0f 06 05 0a 00 07 0c 0d 10 1b 1c 1c 0a 12 12 0b 1c 19 1f 21 2a 31 20 23 2c 33 26 33 33 44 39 3b 3b 35 36 49 43 5f 61 5d 70 63 6c 66 66 66 68 64 5a 5e 66 84 8f 7f 75 60 7c 7e 7f 61 42 35 2f 28 32 38 42 4f 6c 61 48 47 4d 42 31 34 3d 3b 30 1f 20 23 23 1c 24 13 1a 19 0e 15 1d 1b 1f 10 13 15 10 0a 05 0b 04 0c 05 03 0d 0e 05 03 00 06 10 08 00 06 05 03 02 06 05 03 00 06 05 09 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 15 0e 0d 00 06 05 03 00 06 0e 08 0c 0c 0d 16 16 0d 06 08 0c 0d 14 13 16 2e 3c 27 09 09 16 15 19 20 2d 4f 41 3b 2f 25 34 40 36 32 40 43 46 40 53 7d 89 87 85 71 67 74 7f 7c 80 7d 8a 8d 8b 96 9f 87 8a 9f a1 a4 9a 90 9f a4 8f 81 6f 5f 63 60 5d 62 5b 70 8f 76 7a 75 64 4d 45 40 52 51 4e 40 3f 2e 35 2e 29 2f 28 27 1c 19 21 1c 21 18 1b 19 18 0b 12 0f 14 0b 05 03 06 06 0a 11 06 06 0e 03 00 06 05 06 00 06 06 03 00 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 05 0f 24 1e 1b 0f 0d 05 03 04 06 05 0d 0b 06 06 09 12 0e 0c 0d 10 07 14 11 16 1b 1e 23 1a 16 1b 10 22 42 71 73 5b 45 2a 2a 33 3c 4a 5c 65 77 8e 79 8b a8 a5 b0 a9 a9 a0 a2 ab b0 b5 ab af b5 bc ce df d1 c8 c6 c6 cb c4 c4 b4 b0 a9 94 89 87 89 8c 8e 92 89 8b 89 76 79 6f 61 5f 58 50 5b 64 6d 65 5c 57 50 4e 52 47 3e 37 32 29 30 23 30 3a 35 35 26 15 1b 17 1c 1e 0a 10 0b 0c 0e 0d 12 06 0f 07 12 0a 0a 0b 03 06 05 03 06 06 07 03 04 06 05 03 02 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 08 1a 14 13 0f 0e 06 03 00 06 0d 07 04 06 06 03 10 14 20 2b 1d 17 14 1b 13 17 14 1a 20 28 23 20 30 4b 72 75 5e 3b 36 4a 60 72 88 b0 a5 ad ae a7 a1 a2 ac b1 a7 af c6 d2 db dd c8 bf bb b4 cd cb df db d8 da df d9 d8 dd c9 d1 cf bb b3 a1 9a 9d 91 9d 97 99 98 8f 82 85 80 80 75 73 78 71 6f 7b 7c 7b 76 6c 6b 60 64 4e 4c 48 48 43 3d 37 3a 34 2e 27 2a 1b 21 20 13 10 17 15 14 14 19 0d 0e 10 0e 0e 11 0a 05 08 05 03 07 06 07 03 00 06 05 03 00 06 05 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 16 0e 03 07 0c 05 03 04 0b 05 0b 0a 06 0e 0e 08 0e 1a 19 12 25 21 25 1e 18 20 34 29 35 2c 35 42 43 54 64 60 5c 62 78 92 a4 c2 c7 ce d8 d2 d2 d6 e5 df eb e0 e7 fd ff ff ff ff f3 f0 ef ef fe ff ff ff ff ff ff ff ff ff ff ff ff ff f2 d8 c8 c0 ba b4 aa bc a6 a3 a9 aa a4 9a 9d 9f 9c 9d a1 9b a7 aa a9 a0 98 8d 6f 75 6e 66 5e 68 58 52 3d 3b 1c 36 30 2a 28 20 22 22 25 19 1f 1a 1a 12 11 11 08 09 0c 02 0b 05 0a 05 0b 0b 09 08 06 0f 03 08 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0d 0f 27 24 07 05 07 05 0f 0d 07 05 09 0b 0e 13 18 1f 19 18 21 1f 22 2b 2a 30 2a 2d 38 38 44 45 4f 56 67 67 72 86 92 9c c5 dc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f3 e4 d5 d4 d1 d7 d1 d3 d4 cd d5 cc c4 bd bf c5 ba be bc b4 9c 91 89 90 95 90 86 6b 6b 67 71 62 4e 3d 3d 34 2a 28 2a 25 1f 20 25 20 1d 1f 1b 10 13 13 06 0b 0c 0b 0e 09 0d 0c 0d 14 03 06 06 05 04 00 06 05 03 00 06 05 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 12 03 0d 17 15 10 09 06 12 1d 1f 21 11 14 14 14 29 28 21 1f 2e 38 3a 4c 4c 3e 40 42 44 53 5b 5d 64 79 8e a1 a8 b2 c9 d9 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e8 e2 e2 e3 e4 df e4 e9 e3 e0 d0 c9 c7 bd b4 a5 a0 94 93 92 96 9d a3 97 86 8b 9e 9c 94 83 6c 68 5f 51 45 3e 35 32 2c 2f 24 27 21 1a 21 26 18 1b 14 12 10 08 06 12 09 19 31 07 0b 06 05 05 06 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 06 06 05 0a 04 09 0c 09 10 0e 11 25 24 18 12 18 1f 2c 34 29 34 3c 44 4f 5f 64 57 5c 60 65 73 71 71 7c 87 a0 b0 cf ea da e8 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ea dd e1 e1 d5 dc d7 d8 d5 ce c7 c0 b5 ac a0 9e 92 99 8a 82 8d 8a 8a 8d 8b 91 9f a2 9e 95 8e 85 7c 73 6e 74 5f 56 52 40 42 3e 2e 3a 2b 22 1f 22 1a 1e 14 13 17 0e 0e 11 12 06 06 07 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 09 05 03 05 06 05 04 0c 06 08 05 04 06 05 06 01 06 05 05 15 0e 08 12 1f 17 15 22 1a 21 1f 2b 35 3a 45 47 50 51 6c 73 77 6f 75 75 8f 9d 9d 99 99 97 99 a4 b2 b9 c7 d3 d4 db e5 e9 ea f3 fb ff ff fb fd fb f0 f7 f5 f5 f1 e2 eb ee f0 fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 df d5 d4 d6 c9 cc c3 c1 c1 bc af ac a5 9b 9c 91 95 92 8e 93 88 88 8d 8c 84 80 92 8b 93 94 9e a1 91 92 95 8e 93 93 8c 7d 80 68 67 58 4a 39 29 35 2c 23 26 20 25 24 1d 22 17 10 14 18 1e 12 13 11 06 03 01 0d 07 03 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 06 05 05 00 06 07 07 04 06 05 03 05 0f 05 03 07 0a 0e 0c 0f 19 1a 23 2a 27 20 1f 2c 2a 3e 43 57 66 6f 7b 74 73 75 87 90 8f 8c 95 a5 a0 b1 b0 a5 9c a5 a3 a0 a7 a6 b1 b4 b5 c2 c4 cd cb cf e2 dd e2 e1 e7 ec ef f3 f5 fb f6 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ed e3 d2 bf c6 ca c2 ba ba ad b1 b0 ae a6 a3 a3 9d 9d 99 9d 98 94 8e 85 8b 8d 88 85 8c 8b 94 8f 8c 8b 8b 87 90 93 93 99 88 9e 91 89 7f 74 5a 57 4f 47 47 42 33 34 39 31 30 2c 28 2a 1f 22 14 0f 1b 12 0c 12 0e 08 05 03 03 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 06 05 03 00 06 06 05 05 0a 07 03 0a 0f 13 15 18 1a 1d 2d 34 35 3e 47 50 52 5b 60 6f 8b 9d 9f 8a 8d 8f 93 9d 94 9d a2 9c a0 a4 a2 9f 9e 98 a9 a6 a8 a3 b7 bd b5 be c9 c9 cc d7 dd e5 f1 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fa f6 ef f5 e9 e2 e0 ce cf c0 bf be b9 ad a9 ac ae aa ae ab a5 a6 a4 a5 a6 a1 9d 9a 96 95 90 88 90 93 9a 99 95 95 88 86 87 8e 8f 88 89 8c 8d 8a 90 88 7f 7d 78 73 80 7c 71 59 43 35 37 3b 38 2f 42 32 2a 22 29 23 28 1a 19 11 11 08 05 0e 00 06 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 0f 05
 03 02 06 05 03 05 08 08 05 06 07 0b 12 18 1b 11 11 18 11 1b 1f 23 31 31 3c 43 54 61 66 6f 77 78 83 8d 9f 9c 8c 89 85 8c 92 90 97 9b 98 91 97 9a 9f a6 a8 b5 ac b4 b9 b7 c5 c9 c7 cc d2 dd e4 e7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f2 e8 df d6 df d2 d4 ca cb b9 c0 be ba ba b0 b7 b3 b5 a8 b1 ae ad af b1 b4 a3 a9 a5 9b 9e a0 98 a4 9f ac a8 a6 a3 a3 a0 96 95 94 92 92 96 8e 8d 8a 7e 80 8a a1 b7 b4 9d 8b 76 73 5e 56 5e 5e 52 4c 47 32 34 2e 32 2f 2b 26 1c 22 15 09 09 0a 0c 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 0d 08 08 03 03 06 06 07 08 0b 0e 03 06 12 08 18 1c 1b 14 16 23 19 29 39 49 56 5a 63 69 78 7b 7b 82 84 82 83 80 86 81 80 89 84 83 88 8d 97 94 92 9f a2 b0 af b9 b9 b7 c1 bd c6 c6 d5 d3 dc de e9 f1 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa eb e1 dc d4 d6 d2 c6 cb c5 c8 cd c0 c3 c1 c0 c0 bc b6 b9 b5 b9 c2 bb b8 b1 aa b2 ab b1 af a5 b6 ae b3 b6 b6 aa ab ab 9d a6 a1 9e 99 9a 89 81 84 8a 95 b2 c5 cf c7 bd a0 8d 9c 8d 88 89 75 6e 5e 58 50 3b 42 39 32 34 33 26 20 18 15 0a 09 0d 0c 05 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 06 06 03 06 07 0f 0b 0f 11 17 16 1d 1b 22 26 2e 31 40 54 66 7a 79 87 86 75 79 77 7e 85 82 7e 7e 7b 7f 80 81 81 7f 8f 92 99 9d 99 9f aa ac b7 bc c6 c8 c5 ce cd d4 e0 e4 e6 eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e6 dd e2 e0 da da d7 da d0 d0 d0 cf c6 c8 c0 c5 cb c0 c1 c4 c0 c1 bf b4 bb c5 ba c1 bf bb be ba be c1 b6 b8 b1 ae ae ae a2 9e 91 80 7a 89 80 95 a2 ae be c1 c9 c4 ba b4 b3 a6 a0 96 7e 78 71 64 56 56 52 47 42 3f 31 30 1b 0f 0c 14 09 08 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05
 06 19 0b 0b 07 09 06 09 17 16 18 20 1f 24 23 2d 3b 42 4e 55 6c 93 b5 94 84 79 75 79 7d 83 83 82 88 80 84 88 8b 83 89 93 97 95 a3 a4 b3 b1 ae bf c9 d1 d9 d4 da e2 e9 e7 f1 ea f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f8 f2 e6 e4 e4 e5 e0 d8 e6 df dd d9 d3 cb cf d1 cb ce c6 c9 ca d0 c8 cb cf d0 d1 c4 d1 cd be c4 bd bd bf b6 b8 ab 9b 9d 96 81 83 80 89 84 8c 8e a1 af be c2 c9 cf ce c4 d0 c0 b3 aa 99 7e 76 71 6a 69 62 57 39 2b 23 22 18 15 11 0e 06 0b 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 06 0c 06 06 0e 12 18 0e 0f 11 0f 1a 21 1d 28 22 2c 25 2e 36 38 48 5c 61 74 81 a0 c3 a2 84 70 79 7e 81 8f 7e 87 80 86 81 98 89 97 92 a1 a1 a1 b2 b3 be bc ca d3 d3 da e3 e2 f4 e9 fa f1 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 ff f4 f4 f1 f1 ec e9 e9 e1 e5 dd dc d2 de d4 d5 da de d6 e0 db da df d4 d4 d4 ce ca c9 bd bc b3 bb b5 ad ab 9f 9f 96 92 84 87 90 8b 88 86 93 9a 9e ae ae af d1 d5 d0 cf ca b4 ab 8d 7c 7c 85 7e 6e 5f 4f 36 33 24 1b 18 19 12 0e 0e 0d 09 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 07 05 06 00 06 08 09 00 06 0d 11 1a 13 1d 20 1c 2a 25 2b 36 2d 34 34 3e 4e 55 66 7a 91 94 8e 99 b5 9b 7d 85 82 81 83 81 84 8d 8e 8f 90 94 90 99 9e a7 ac b2 b8 bd ca cc d1 da da ea ee f7 f6 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe f8 f8 f3 ed ea f0 e7 eb e2 e2 db e4 e2 e3 ed eb e6 e1 de db d8 cb cf cb cb bd bf bc ad b3 a5 a6 a9 a0 97 98 91 8b 8f 96 95 8d 8a 8c 8f 96 96 a9 ae b3 b7 b3 b7 ac 9b 94 9a b5 b1 9f 84 72 56 4a 37 34 20 19 10 0c 11 0a 06 0a 07 05 03 00 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 06 12 09 0d 09 10
 11 16 17 20 26 2f 34 3a 3d 3d 41 53 59 6c 76 84 89 8e a0 9d 9f 9c 96 7f 79 80 84 8a 85 87 8d 8b 92 98 9f 99 99 a0 aa ad b4 bb c4 c9 d1 d4 db e5 ec f0 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff fe f0 f4 ef f2 f5 f2 ee ef f5 f7 f3 f0 ec dc de d8 d6 cd d1 c7 be ca b5 c1 b8 ba b5 bb a5 a6 a2 a4 9f 9f 98 9d 97 95 91 8d 8c 8c 92 90 8d 8e 94 93 98 a8 b0 cf e5 dd bf 9f 8f 7e 6e 5e 4f 39 29 0d 12 13 0b 03 0f 06 06 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 04 06 0c 08 05 08 0c 08 13 11 1b 25 29 2b 3c 41 57 5e 6c 6a 6b 74 82 90 97 9e a0 9c a0 a3 9c 94 8c 89 87 8b 8d 8e 88 8a 8e 94 92 96 97 9e a2 a5 af af b0 bd bb d0 db d9 e0 ea eb f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff fd fa fd fe fb fd ff f4 f0 e5 df e0 df d7 cc d4 c4 cb c4 c2 c3 c0 c1 b7 b9 b4 b5 aa a2 ab a8 a3 a6 a2 9e 98 9d 8d 94 9f 94 95 8e 8d 8c 93 aa e2 f2 ff e9 ca ba a5 8d 82 69 4b 3f 25 1e 12 0c 06 07 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 09 0e 07 0f 15 10 1e 20 2f 33 4c 5f 79 83 93 a0 a9 a7 aa a8 ae b3 c2 b5 ad 99 8b 87 7f 85 88 90 91 94 90 99 99 94 9a 9a 97 9c a3 a8 b4 b0 b6 be c0 ce d0 d5 e0 e9 f4 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f6 f0 eb ed e8 db dd da d7 d3 d4 c9 cd ca cf c7 c6 bc b7 bf b5 b3 b6 b1 ac ad a7 a6 a2 9f 9e 97 9c 96 91 90 90 87 81 92 c7 fa ff ff fb e1 c7 ba 9a 8a 68 56 41 2c 1f 1a 0c 0f 06 06 03 00 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 07 0c 0e 14 0e 20 21 2a 2d 30
 35 4e 74 8b 9a b5 c2 ca c6 cb ca cd cf d4 ce c5 ae 91 8b 8c 8e 91 95 9b 9d a2 99 a4 9f 9b 9f ac ac ae af ba b2 b8 bb cb d5 d6 d6 e1 e1 f1 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f6 ec eb e8 df dc d5 d7 d3 d3 da d4 d2 d2 d1 cf c4 c5 be b9 ba bc b2 aa ac ac 9d a7 a5 9f a3 a2 9c 99 8e 8f 82 8c 9b d5 ff ff ff ff f1 df d1 bb 98 7b 61 50 35 27 18 0d 08 05 03 06 06 05 03 01 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 08 09 0d 15 19 1d 24 27 2d 2c 36 3b 51 77 9a b0 c0 d4 e8 f5 ee ea e4 df e0 d9 cf c0 9c 8c 8a 89 91 9e a3 a7 b2 b6 b5 b1 b4 b2 af b6 b7 b8 bf c0 b9 c1 c6 d7 de de f0 e8 f2 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f7 f9 e9 eb e2 e5 e3 de d9 d5 dd d9 db db d7 c8 c6 c8 ce c6 c4 bf be b6 b1 ac b0 a7 a8 a8 a0 a0 8f 98 90 8c 91 99 a2 d0 ff ff ff ff ff fa e6 b7 8a 79 6d 60 3d 35 22 16 06 0e 09 06 07 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 05 07 0e 09 0a 12 15 21 21 2b 2a 35 37 41 56 55 8a aa b6 d3 dd ec ff fd f3 ee e0 d5 d1 bc b0 a2 93 96 93 9c 95 a7 ac b2 ba ba b6 be ba bc c4 bc c5 c6 cb c9 c8 cd d5 dd da e6 f1 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f7 f6 fb f9 f0 f2 df e9 e4 e1 db e6 d8 e2 d8 d8 d5 d0 d3 c6 c8 c0 c2 be ba c0 af b1 b1 ad ac a6 a5 98 9a 94 8f 99 98 a6 c7 f1 ff ff ff ff f6 c5 ac 91 87 79 62 57 38 23 0d 05 03 0b 05 07 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 08 05 03 06 06 05 05 11 1d 0c 1c 29 29 35 34 31 2c 3a 52 64 6c 92
 b1 c6 da e2 e7 f2 f7 e7 d8 d2 be b8 ac 9e 9b 94 93 97 99 a7 aa ae ae b9 be c1 c6 c6 cb cf c6 cf d2 cf c9 d5 da d6 e3 e2 ef f4 f6 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff fe fc f2 ea ec ed e9 e9 ed ec e4 ec e4 d2 da d4 d1 d6 ca c9 c7 b9 bb b9 ba c0 b6 ae af a8 ac a5 9d 92 8e 94 97 96 96 b2 d0 e2 f7 e6 dd d4 c5 b3 a6 9d 84 63 4e 35 1a 0f 02 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0b 05 05 13 14 17 1f 23 30 3b 42 40 41 32 32 35 3e 58 71 69 86 a2 b9 ca d2 cf dc db cf cf bc b6 a8 9b 9c a0 95 9a a3 a0 a5 ae a8 b5 c3 c5 ca cf cd d7 da d6 db db dc d8 da e5 e2 e0 dd ec f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f2 f3 ed ea ed ed eb ec c7 e3 db dd dc d7 d5 d1 d1 ce c1 bc c7 cb bf bf c0 b0 b5 ad ab ab a6 97 9a 96 92 93 89 97 a7 b6 b6 b6 c8 d7 d2 cc c4 a0 7f 67 4c 31 25 13 0c 0c 09 0a 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 08 06 08 19 17 1c 1f 24 37 49 52 50 4c 44 42 43 47 51 5c 71 6b 70 8c a4 b9 b5 ad b0 af af af aa a6 9f a1 99 9f 9a 9b 9f a2 a4 a9 b9 b1 bc c2 c4 db d1 dc d9 db e4 e2 e5 e5 ec e8 f3 f2 ee f8 fc fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 f7 f4 ea e9 f5 eb e9 f1 e0 e6 de d9 d2 d6 cf d5 d4 cb cb cb c2 c1 c8 bc b6 b7 ad b0 a4 a3 9b 98 95 8f 8b 8f 93 96 9b 9e 9a a6 b9 d9 df d1 bb 99 71 54 44 32 21 14 06 11 00 06 0c 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0c 1e 1c 1f 20 1a 37 48 4f 53 4f 47 3d 40 40 57 69 70 7e 84 85 91 9a
 a6 96 8c 97 95 98 9c a0 a4 a6 9a a6 98 9f a2 a5 a4 a0 af b6 bb ba cc d1 d4 d0 dd e0 e5 e3 e9 e9 f0 ee f2 f5 f0 f7 f2 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 f1 ee f0 e8 ec f2 e4 ec e6 e1 e3 dc d7 d0 d3 cc cd c8 c6 c2 c2 c2 ca c0 ba b3 a9 a5 ac a0 9c 98 96 93 8f 84 8f 91 9c 9a 97 96 9a b9 d7 db d0 b1 90 7a 58 49 29 1b 18 07 03 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 0b 0d 14 16 22 27 2c 2a 3c 53 59 4f 41 41 44 48 52 67 77 83 91 93 94 9c 94 89 8d 8a 87 8f 97 97 9d 9f a7 a0 a4 a0 a1 a8 a9 b1 ae ae c2 bd c6 c7 d2 d8 d6 dc e4 e8 f4 f1 eb f6 f5 f9 ff f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f9 f5 f6 ed eb e6 eb ec e3 de e0 e0 df d8 d5 ce d2 cf c8 c5 ca c8 c7 bb c5 bd b4 bc ac a9 ab 9f a1 9c 96 96 99 90 9a 99 95 8d 94 90 93 b6 cf db c9 b4 95 74 52 3a 21 18 0f 0a 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0a 06 08 0c 0d 21 28 33 33 3b 48 53 57 56 38 42 51 4c 63 73 7b 82 88 8e 8a 92 93 8d 8e 8b 93 95 9b 95 a9 9e a7 a9 ab ad ad b3 ae b3 b1 bb ba c7 cf d5 cd e2 dc e1 ef eb e9 f4 fc f8 f6 ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f6 f1 f4 e6 eb ed e7 e6 e5 e5 e2 e9 d7 d8 d1 d2 cc cf ce c8 c6 c1 c3 ce c3 b8 b6 b1 b1 a5 aa a6 a1 9d a0 98 9b 9c 94 9a 9b 99 90 8e 90 96 a3 c5 d4 cc a7 92 6c 49 2a 1f 14 0b 0f 07 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 08 10 20 30 2e 3d 3a 4f 6c 6e 5a 4d 54 5e 5b 6e 74 74 77 88 8f 8f 8f 89
 91 8e 90 8f 92 97 a1 9f 9d a7 a9 aa b3 b6 b4 b9 b4 c0 b9 c0 cd c6 d5 d4 dc de e1 e4 eb ea ee f7 f8 fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 fe fd f6 f7 e7 e5 e8 e9 ee ea dd e6 df db d7 de d2 d3 ce c7 cb c5 ce c6 cb c1 be b5 b3 b1 ab a4 aa a7 a1 a2 9e 9b 9e 97 a3 9d 99 9e 93 8a 8d 8b 9b bc d0 cc a5 7a 5a 35 24 18 21 1c 0b 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 06 05 03 0b 07 06 11 1a 1f 2b 40 46 4d 62 6f 79 69 57 5e 6f 75 7b 7b 78 84 88 7c 8c 89 8e 8d 8b 95 9d 9b 9a a0 a5 a4 aa b1 a9 ba af b8 b9 c8 c5 c7 c1 cc d1 da dc e4 e8 e3 ef e9 eb f1 f6 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd f9 f8 f1 e9 e8 f1 e2 ed e4 e3 e1 d7 da db d9 d5 cc d1 ce d1 da cf c6 cb bb be c2 b7 b3 a9 a9 ae a3 9b 9d 99 a1 9d a2 9f 96 98 93 88 8d 81 8f a4 c2 d0 b7 89 56 34 20 25 1f 1d 15 08 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 0b 15 07 0c 1d 23 3a 40 56 60 71 78 7b 7c 7a 6c 73 76 7d 7c 85 80 87 86 8c 8d 92 94 9e 9f 97 98 9c a1 ad a8 ab b2 b2 b1 b7 c1 c0 c9 c5 c5 c1 c7 d8 d4 de e4 e2 ea ed ef ea f0 ef fd ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fb fd fb ee ea e5 e9 f2 f2 e6 e6 e4 df dd da e1 d5 d3 d0 d7 d3 ce d3 d0 c5 c5 c5 bf b3 b3 b0 a4 aa aa a5 a4 a1 a1 a3 a5 98 9e 92 90 8b 88 87 87 98 9f b3 b7 9a 65 37 31 2b 1a 1a 10 03 00 06 05 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 08 0c 03 06 08 03 0b 0d 1c 2a 39 42 53 68 7b 80 87 7a 76 75 6f 70 73 80 7e 7d 82 82 87 8b 90 a0 a8
 aa a0 9e 9f 9f 9f a6 a9 ab b2 ad b7 bb b5 c8 c2 c3 c9 d2 cd d4 d8 e2 e9 ed e5 f3 ea f4 f3 f4 ee fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fb f9 f4 f4 f0 e7 f1 ee e6 e4 e8 e3 dc e2 db da e0 d4 d7 d1 d3 cc d4 cd c7 c4 bf b5 b3 b6 ad b2 ae ab a5 a9 a6 9b 9f 9b 95 94 8f 8c 8f 83 85 8e 90 aa c5 a7 7a 54 40 34 25 15 08 0c 05 06 06 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 06 0a 12 05 0d 19 1c 2d 48 54 60 70 71 80 80 8b 7e 82 70 72 79 6e 75 7b 7c 7e 7f 8b 93 93 a4 a8 ab a4 a0 98 9d a4 a7 aa ae b2 ae b9 b9 bb c0 c2 ce d1 d0 da d9 df e5 e3 ea eb ec f3 f3 f7 fc f7 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f6 f6 f7 f8 ed eb f0 f1 e5 e7 e7 e5 dc e1 dc e0 dd d7 d4 d5 d1 d3 d4 ce c9 c8 c1 b8 b5 b0 b2 b0 b1 af a9 aa a3 97 ac 9f 9d 8a 87 85 8e 86 88 87 90 9a bb c0 a3 81 6a 4c 29 13 0a 0a 09 06 06 06 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 10 0c 12 17 1a 19 30 42 5e 6b 78 86 80 7d 7f 88 83 87 7b 7c 7b 79 7c 85 83 8d 8f 92 95 9f 9f a6 b0 a8 9f 9c a0 9d a8 b1 ad b6 b6 b5 be b9 c6 ce cf d1 de e0 e0 e0 ea e7 ec ed f6 f9 fd f9 fc fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f8 f1 f5 f2 f4 f1 ea e5 dc e0 de db db e0 e1 dd da d4 d5 d0 d0 c9 c6 be b6 b8 b0 b7 b4 b3 b8 b5 ae b0 a2 a5 93 94 92 87 82 84 83 80 83 83 97 c6 d3 c4 ae 88 6e 45 27 13 0a 0a 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 0a 0a 0c 10 0f 13 1b 2c 3b 5c 6f 74 85 92 8d 84 7f 7f 78 73 7e 79 84 81 80 83 8a 8b 92 8d 98 9d a5 a1
 ab 9f a2 9f 9d 9b a7 ae b3 b8 b9 b9 b7 c9 ca d5 d5 d4 e0 e2 e6 ee f0 ed f8 f2 f6 f5 f9 f5 ff ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 f7 f8 f5 f2 ed ed ea df e2 e0 db e2 db dd da e0 d2 d4 ce d0 c6 c6 bc b9 bd b9 b8 b9 b4 b8 b5 a4 aa 9c 9e 93 91 91 90 81 88 81 81 84 87 8a a2 ba c5 cb bd 8d 5b 41 1e 19 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 06 05 03 09 0b 0a 09 10 14 1a 28 44 51 6f 80 86 95 94 a1 93 85 83 7e 75 72 7e 81 86 86 8e 89 8d 94 98 9b a5 a9 a8 a7 a7 a8 9f a2 9f a5 a9 b5 bc b7 bf be bc cb cb d8 dd e2 eb ef ef f4 f1 f9 f6 fd fc fd ff ff ff ff fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f9 fb f6 f7 ff e8 ea ec df e5 e8 e3 e1 e0 db de da d8 d1 d3 c9 c8 ca c0 b7 bd b0 b8 bc b9 b6 ae aa a1 9b 94 9c 97 8a 90 89 8e 84 85 87 7f 7e 88 94 98 a3 b2 a9 84 5d 35 1a 14 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 06 0a 1d 1e 1f 27 43 54 62 7c 99 a5 a9 ad a7 a3 97 8c 7f 7a 76 77 7e 8e 91 96 93 92 8d 98 99 9b ab b1 a8 a6 a5 9e a5 ab ad b4 b4 bc b8 bf c7 cc cb d6 d5 dc e5 e7 f0 f4 f6 f6 f5 fa fe ff fa f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa f8 f4 f6 ed e4 eb ee eb db df e0 e3 d9 cd d1 cb d4 c1 c0 bf c1 bb bc bd be bb b7 af ad a8 ab a9 a2 9e 9d 95 94 8d 8b 8a 85 86 80 89 83 90 8f 86 89 a8 99 7a 50 2b 1a 06 0e 03 00 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 07 12 12 18 1b 29 38 4f 60 7e 93 a4 b3 b1 b0 a9 b0 a3 9d 76 79 86 86 7e 8c 88 83 96 8a 91 a5 9c a0 a6 a3
 ad a7 a4 9c a7 aa b0 b8 ba bc c0 c9 cf d1 d4 da db da ed f7 ea f6 f7 f7 ff fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff ff ef f7 f2 ec ed ee e9 e3 dd d5 db d7 d2 ca d2 c9 c2 c3 c0 b8 bd c3 bf bb b9 b5 b2 bc af ad a6 9d 9a 97 9b 94 98 8a 84 8b 8b 8a 8c 8a 89 8e 8d 9c ac 96 74 3e 1d 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 07 05 07 04 0b 1f 1f 25 43 54 6a 82 97 b0 b6 bb b5 b2 ac a7 ab a2 93 87 80 7e 89 89 8d 90 8e 9d 9a 98 a0 a7 a3 a6 a5 ad a7 a8 ad a1 af b7 bb bb c9 c8 d4 d6 d1 db e6 e2 e3 f5 f7 f0 fd ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fe fa f6 f1 ea ed eb e3 e4 db db db d5 d2 d0 c4 c9 c5 be c0 bd ba b8 be c0 c1 b8 b5 bc bb b6 a6 a2 a3 a0 95 98 9e 8c 8d 8f 8f 85 8a 86 87 8b 86 92 a6 aa 8c 5d 27 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 05 09 1b 11 20 2f 46 5d 76 98 a2 b1 b5 c6 c5 c7 b4 a9 9f b0 9e 9a 89 8c 89 90 8f 96 9e a2 9f 9e aa a2 a3 a8 a2 ad b4 ae a5 a5 b1 b2 bf cb be cd cc d5 dd de db e1 e7 ed ef f3 f8 fd ff fd fc ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff fb f3 ee ee f0 ee e9 dd d7 d4 d9 d2 d4 d1 c7 c7 c9 c5 c2 c4 c1 c4 bf c4 be bf b8 b6 aa b3 aa af a2 a9 97 9b 96 98 98 93 90 93 8f 90 87 8e 90 94 ab 9c 62 3c 19 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 04 08 06 08 14 15 1f 25 4a 69 80 94 aa b5 c7 c7 d2 d0 c7 ba a1 a0 98 9c 8c 91 90 92 8e 92 96 94 9e a1 a4 b1 ac a3 af b2
 af b1 ae ad b0 af b8 b7 c6 cc cc d5 d5 e5 d3 e1 eb eb f1 f1 f8 fb f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f4 f8 f1 ed f3 e9 e1 e2 e1 dc d9 d4 d3 d2 d0 c7 c6 c5 c4 c7 c8 c4 c4 c4 bc bf b7 b6 b2 ae a4 a8 a4 a6 9b 9e 91 9e 95 95 8f 8e 8d 90 85 8d 87 97 8b 6e 3e 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0a 09 08 08 12 17 24 3b 65 8d a6 b1 b1 cb cf d9 de d1 c8 b1 a5 97 95 8d 92 99 94 90 92 90 98 95 9b 9b a5 b4 aa b1 b2 b4 b7 b8 b4 b3 bc b0 c2 bf c7 d0 d7 cd d9 dd e4 e2 ea ec e5 ea f1 fd fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f7 f6 eb f7 e5 eb e5 dc df d3 ce d1 ce d1 cb d6 c5 c9 c7 c5 cb cc c6 c9 bd ba b3 b8 b0 b1 a5 a5 aa a4 9f 96 9c 96 8f 90 92 8d 87 8c 8b 85 8c 85 84 6b 41 15 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 04 0c 06 11 25 29 4b 76 a5 cc d6 da d9 e1 e1 d6 c9 b6 a4 a4 a0 90 96 94 92 92 98 96 96 9c a2 a4 a3 a5 b6 b7 b4 c0 b6 bf bf bb be b6 bc c5 cb ce de d7 d8 dd dc e2 e5 e9 e9 f1 ef f0 f8 fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f8 f2 ef f1 e7 e7 e4 e3 e4 dc d5 d1 d4 cb c7 c7 ca ca d0 c9 c5 cc c6 be c4 b7 b7 b0 b1 b0 a6 a9 af a1 9e 9a 97 94 97 8d 9c 97 8d 88 8b 8d 80 8d 8b 75 43 1a 05 07 06 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 06 0d 0d 0b 10 0e 1e 25 43 66 8a b9 e1 ea f2 eb e6 d6 c4 b0 9f 9b 9e a4 9e a1 9d a0 96 9b 91 99 a1 a3 a6 ac ac b7 bd c2 c1 c6
 c3 bd bc c5 c7 cc d5 d2 d3 d9 d4 e3 e2 df e9 e1 e7 ec ef ef f6 f8 f6 fd ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f9 f9 f4 f3 de e3 e7 db de da d1 d2 d0 cb cc d2 d1 cb d3 c9 c9 be b3 b1 bb ac ae ae aa aa a6 97 a3 9c 9b 9b 97 96 90 93 8e 8e 8f 90 8e 8f 87 77 41 15 0c 07 02 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 09 16 1b 28 56 7d a3 ca f2 fa ee e9 dd c5 b1 a0 99 91 97 a2 a5 9d 9e 9c a1 98 99 9d a9 a3 a6 ae b3 bc bb c6 c1 c2 c9 ca c4 cc ca cf d5 d6 d7 db de e3 dd df dd e4 ec e4 ed f0 f3 f8 f2 f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fd f4 f3 df e1 d5 d6 dd d9 d4 d2 cd d1 c9 c7 d5 cc ce c5 bf be bc b0 ad b4 ac a3 a4 99 9b a1 97 97 98 9a 95 9b 92 8e 92 96 8f 8f 8c 84 80 69 3c 1f 0d 09 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 0b 10 19 20 36 5c 9b c4 df f1 e4 cf ce c0 ac a8 9d 9e 99 95 98 a2 a1 a2 a9 a7 a1 a6 ab ac ad a3 b3 b7 c0 c1 c1 c6 cb cd c9 c9 ce d0 cb dd d9 da e1 e4 df e5 e5 e5 e6 e9 e2 ed eb f3 f7 f9 f6 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 fa f6 f3 f0 eb de de df df d3 d8 d2 cb d1 cf c9 d1 d3 cd c2 bd b9 ba ad af a6 a2 a9 9f a2 9a a1 9e 96 9b 97 99 99 95 91 94 91 9b 9d 91 84 83 60 3c 19 0e 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 01 07 05 0d 12 15 22 24 43 61 aa d7 e5 d6 b0 aa a1 9a a3 9c 9d 9c 99 94 a0 9a aa a3 a7 ad a7 aa b0 b0 b8 b5 bf b5 ce d2 cb d2 d3
 c4 cd d5 d2 d3 d2 db d1 dd ec ea e5 ed e7 e8 e7 ed f0 e8 f1 ec f1 ff ff f9 f7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fd f9 f3 f1 e8 e8 e3 dd e1 de da da d0 d3 db d5 d2 d1 d0 c1 c7 b9 b6 ad ae ac a9 a6 a4 a1 9a 9d 9b 94 98 97 92 96 95 98 92 96 98 99 95 88 7d 78 64 32 1c 07 05 09 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 0f 0b 1a 19 33 4d 70 9f cc d1 ad 9d 97 99 95 93 97 96 95 98 9a 9f a5 a2 a9 aa af b8 ae b2 ae bc b8 c1 c2 c4 c2 ca ce c9 d4 d0 ce d0 d0 d5 d6 da e4 e0 e5 ed eb ee ed e9 ec e7 f0 eb f3 ff f9 fc ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f5 f7 ec ec e3 e3 dd d9 db e1 db db d9 da da cc cb c6 c4 bf b7 bb b1 ab a5 a6 a7 a4 9e a0 94 9e 94 9b 99 98 92 94 8f 96 97 92 8d 8c 84 81 7b 57 24 13 13 0b 09 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0f 10 13 25 3c 5b 7e 91 ae b1 99 99 8d 9b 95 92 96 97 9f 96 97 a1 9e 9e a2 ab af b1 b3 ad b9 bf c4 c4 c1 cd c9 ca d3 ce d5 d0 d7 d0 d0 d8 d9 d9 db f4 e8 ec f0 e6 e6 f0 f0 eb f5 ee f4 f7 ff f9 fd fa f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f4 f6 f6 ea e3 e3 dc e4 d7 da e2 df e2 d9 e0 d9 c2 c8 bc c7 c4 b2 b3 b5 ab a4 a7 a4 a3 a1 9a 97 9a 93 8a 95 92 93 99 96 8f 90 8f 85 91 80 80 76 49 2b 16 11 09 03 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 07 06 0c 0d 14 15 33 52 73 95 94 a6 a8 a2 97 95 9a 94 9d 9c 9f 9f a3 95 a4 a5 a5 a0 b0 b4 b4 b7 b3 be c2 bf c8 cb c9 c9 cc c6 ca
 d8 d0 d4 d9 d3 d9 d8 d5 e5 e5 ec ee ed f4 f3 ee fb ec ec f9 f7 f9 fe ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 fb f1 f0 ed f2 eb df e7 e2 e7 e9 ec e2 da d1 d3 cc cc c7 bf be b4 bd b8 b5 bc a6 a8 a2 a3 98 9b 98 90 94 96 98 90 96 8c 92 94 86 8a 8b 89 7f 74 48 21 0f 0c 0f 07 06 05 03 05 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 08 0f 0f 1a 2c 58 86 a9 ac b2 ab 9b a1 9b a3 9b a1 a3 a0 a3 a4 a5 ab aa a7 ad ae b2 af b4 b6 b7 c2 c4 c0 c1 c9 cc cf ce d4 d4 d0 d0 d3 dc d2 d4 dd e4 eb ec ef ef f0 f0 f5 f6 f3 f5 fd f8 ff fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 f8 ef f2 ed ee ed ed e2 e8 e7 e5 e2 d8 d7 d5 cc cb c6 c5 c2 c0 ba b9 b8 af b1 a0 ac 9d a1 9b a2 9b 92 8d 96 8d 8c 96 91 90 8a 8e 8f 8b 8d 80 70 39 1f 0e 10 0f 06 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 01 06 09 07 13 22 42 62 97 b4 bd af a3 9e 97 9f a7 a3 a2 9d a0 a4 a5 a5 b0 a9 ae b3 b0 b6 b5 b3 b6 bc bc c1 bf bf c3 c1 ca cd cd d4 cd cc d0 d1 d2 da dd df e0 df e9 ec f3 f6 f7 f7 fd ff fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe f8 f2 f0 f1 ef e6 ed ee e6 e3 e6 e1 e2 dd d2 d2 cd d0 cb c8 c5 bc c6 bc b4 b1 aa aa ab a2 a7 9a 96 a0 92 9a 94 9a 8e 8c 8b 8d 91 92 8a 8a 7f 77 64 28 14 13 07 0b 06 0c 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 08 03 0b 06 0e 0f 13 25 3e 6d 9c c4 c9 c2 b4 a5 9d a5 a0 a6 a5 a9 a5 a6 a0 ae ab b1 b0 b7 b7 b6 b2 ba b8 bd bb b6 be c1 bf c6 ca ce c5
 ca d1 d3 d1 d7 db d6 df e2 e7 e3 ed f1 f5 fa f7 f8 f2 fd ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 f3 ef f3 f2 ec ed e7 e0 e0 dd da da d1 d5 d6 cb ce c9 c9 bc c3 c1 b5 b4 ae b0 a9 a4 a5 94 9a 9a 9b 96 9b 96 8e 95 8f 95 8f 8f 8a 8b 84 81 5f 37 23 12 0b 06 01 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 03 0e 0b 12 1c 21 33 46 70 9c cd c8 be ac a9 99 a2 a7 a0 a1 a7 a6 a4 a4 a9 ae ae b7 ae b1 b4 be b4 ba b9 c1 c0 bc bf c1 c6 c7 cc cc cc d3 d0 d4 d7 d9 da dc df e6 e4 e2 f0 f4 f7 f4 f2 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fa fb f4 f6 f0 f5 f3 eb eb e4 e0 df e1 de de db d3 cc d0 c8 c9 ca c3 c2 b5 b6 b8 bb b4 ac a3 9e a8 a1 9b 9d 99 9b 98 9b 94 98 94 95 8f 8a 82 73 4a 32 24 15 14 10 09 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 04 04 07 08 15 1c 31 57 71 aa cd ca b9 af 9b 93 9c 9e 9e 9b a3 a0 a5 ac a3 a9 b0 b2 b3 bd bb b1 c1 bd bb c0 b9 c3 be c4 ca be cb c8 d4 cb d9 d4 db d8 d6 d6 e4 e4 e5 ea ed f0 f5 fc fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 f3 eb f7 f1 ed eb e4 e8 e2 dd e1 db e3 dc dd db dc d6 ce d4 d3 c7 cc c6 ba b4 b2 ba af a2 ab a5 a4 9d 9e 97 9b 9d a0 9b 98 90 91 96 8d 87 7c 65 4f 30 35 22 16 0f 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 00 10 13 16 25 3c 5b 88 af ca b2 a6 a2 9c 93 9a 9a 94 9d a2 a6 a5 a5 ac aa af b1 b4 b0 bb b1 b3 b7 be c1 bf c0 be c1 bb c4 c6 c6
 d1 d3 cd d5 dc dd d7 dc e0 e9 e8 ea f4 f0 fd f7 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff f5 f5 f2 ea ef f3 eb e9 dd e1 da e1 df e1 e7 e5 e1 dc df d0 cc d3 d5 d4 d2 c8 bc b5 be b6 aa b5 ae ab ae a6 a2 a0 97 a2 a6 97 99 9b 8b 8d 8b 7f 75 72 59 4f 3e 2d 18 0e 05 06 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 07 0e 09 11 1d 1e 3e 61 91 b2 c0 a6 9f 98 9a 9b 9d 94 95 9e 9f a4 9d a2 a5 ad ad b0 b0 b1 b2 b5 b6 b8 c3 bf c3 c2 c2 c3 c5 ca c8 cc ce d2 ca cd d4 dc dc dd e0 e5 ec eb ef f9 f0 ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff f5 f7 e7 ec ec e8 e5 e0 dd df db d4 db e2 db e4 e4 df e2 d9 dd d4 db d6 d0 d2 cf ce cd be bd c0 b2 b1 b6 aa b4 a5 a6 ad a2 a5 9b 9e a2 96 97 8d 84 79 6c 6f 6e 5b 4c 2c 22 16 06 06 05 07 01 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 08 0a 1b 28 39 66 98 b9 b0 9a 95 92 97 95 93 94 92 9b 9a 99 99 9f a4 a9 ab a6 ab ae ad b6 bb c1 be c0 c1 be be c9 cd c5 bd ca cd ce cd ca d0 db d3 e3 e2 dd ea e5 e7 f1 f2 f4 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f4 f4 ed ee f5 e8 ea e3 e2 df d7 dc d2 d4 d2 d5 d5 db d3 e0 d8 df d6 d2 d8 d6 d7 d2 d1 d3 cf ca c8 c0 b8 b8 b4 bc ae b2 a8 a9 a0 a8 a1 a6 9b a1 9a 8f 83 7b 71 66 69 75 61 47 35 28 18 11 07 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 04 09 0e 13 1a 27 43 65 9b bb b0 91 90 92 95 94 8b 97 8e 96 a2 99 a4 a6 9c a3 9a a8 b1 a8 ba b4 aa b8 be c4 c1 c1 c6 c5 c6 c9 c6 ca
 cd ce cb ca dd d3 d9 de dc e5 e6 e6 f1 f5 f3 fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fc f0 f2 ed ec f4 f5 e4 ee e2 d8 d6 dd d9 d1 d5 d6 d6 d4 d5 de e1 d3 dd df db d9 dd dc d0 d4 d3 d2 cc c8 cb bc c1 b4 b5 a9 b0 ae a6 a5 a0 a0 9e 9f a0 91 86 89 73 70 68 74 7a 68 5f 44 2b 21 11 09 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0c 09 0a 06 16 20 20 3b 64 9a b5 a3 94 92 8b 90 95 94 90 94 94 98 9d 99 a3 a1 ab a1 ad a9 b0 b4 ad b3 b5 bc b9 ba bc c0 c6 c2 c7 bc d2 cd ca c9 cb d5 d3 d9 d1 df e0 e6 e2 f0 f0 f4 f8 fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f5 f0 ed ed ee e6 e6 f4 e5 e5 e5 d7 d1 d3 d0 d2 d6 c6 cb d2 ce d5 d3 dd d7 d5 d9 d9 d5 d6 de d8 cb d3 cc ca ca c0 b6 b9 ba b8 b5 ac ae a6 a3 a3 a3 9a 99 91 85 77 74 6c 73 73 82 75 54 42 34 1c 10 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0f 0c 16 25 3d 6d 95 b5 a7 89 8b 90 89 8f 93 98 90 8e 9a a1 9c a3 a0 a9 a3 a3 ad a4 ad a8 af ba b2 bc ba b7 be bc ca c3 c1 c7 c7 c4 ce d2 d5 cf d8 db dc d9 e2 e7 e8 ef ef fb f7 f4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f5 f0 ea ec e5 de eb ea e2 e2 de e4 cf d8 cd c5 c6 c8 cd cd cc d3 d0 d2 d3 d1 dc d4 ce cf d4 d3 e0 d1 cf cf c4 c8 c3 c2 be bb b4 ab b1 ae aa a5 aa 9b 96 96 8a 81 70 79 70 6f 72 86 74 61 43 29 1c 13 07 06 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 0a 0b 07 0a 23 2b 3a 61 95 b2 a2 8c 92 8e 8f 93 8d 96 96 95 a5 97 a0 a0 9b a4 a7 a2 a3 a6 b1 b2 ae af aa b8 b7 b5 b1 aa c0 bc c8 cb
 cf cd cc ce d9 d9 dd d6 e1 e2 df f3 ed e4 f2 f5 f2 f3 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 f3 ec e4 df e8 de ed e1 e3 dd df dd d1 d3 ce c3 bc c3 bd cc c7 ca cb d2 d9 d6 d4 d9 d4 d7 d2 d0 d7 c9 d4 c4 be c7 c3 c5 b6 c0 b5 bc b2 ae aa ad a2 99 99 8c 77 74 76 6b 73 66 77 7f 81 6e 4b 40 23 10 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 04 09 0a 16 25 2a 3e 66 8d b1 a7 92 8d 8b 93 9e 96 9f 9a 95 9d 95 96 9f 9a 9c a1 a2 a2 a8 aa ae b2 b0 ad b6 b6 b1 bb bf bf be ca bd c6 d0 c8 c6 db d6 da e4 e9 da ea e8 ea e4 ea e8 ed f3 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f1 f0 ee ea e6 e2 e5 e4 e0 dd d3 db d3 cc d4 c4 c7 c7 ba c5 be c5 c5 d0 d3 c8 d5 ce d1 d0 cb d4 d9 d4 d4 cf cd c0 c6 c1 c5 ca b4 b8 b6 b0 ae a7 a6 a1 9c 92 91 73 70 71 6a 67 78 71 89 7a 66 57 37 26 20 0d 08 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 06 05 09 02 0a 10 1b 24 31 5a 85 9f a7 a0 96 91 98 92 99 96 97 94 9a 95 96 97 9b 8f 97 98 a5 ab a6 a1 aa b1 ad ae b0 af b2 bb b8 c6 c8 c5 cb ca ce ce d9 db de e4 e3 dc df e5 e7 ea e9 ec e5 f4 f0 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb ea ee f0 e7 e7 e4 eb e0 e9 e4 da e1 d4 c8 cd c5 c4 bd ba bf be c4 c7 cc c6 ce d5 d1 cd ca cb cd c9 ce cf cb ce c6 c4 bc c0 b6 bb b7 ae a8 a5 a0 a5 97 98 85 7c 70 6d 73 74 70 6e 70 83 7c 6b 5d 35 28 15 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 09 09 10 18 20 36 4c 7d 9d 9b 91 8c 92 96 8d 90 97 95 92 8b 93 95 93 95 9b 91 97 a3 a5 a7 a5 9c a6 a9 b4 b2 b7 b7 bc bc be c9 c3
 d0 cb d1 d9 d5 d9 d8 df d9 e3 e4 e6 eb ea f1 e6 f4 f2 ec fe fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f6 ff f0 ef f5 f6 f6 f9 f9 eb f1 e1 df dd d4 cc c5 c7 c3 bc ba c3 c2 c2 c7 c6 c4 c9 d1 ca d0 cf ce cc d2 d1 cf cd ca be c1 be ba bd b4 ac b4 ae a5 a3 a0 91 8e 84 7e 77 74 6f 70 71 65 69 7c 87 74 56 44 25 20 0c 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0b 05 07 0b 0b 1a 2a 33 50 77 96 95 8e 88 84 85 88 84 86 86 90 99 93 91 95 92 96 95 9b 99 a5 a4 9e 9e aa ab ae ae b1 af b4 b9 c2 cc cd ca cd d0 dc e0 db de e3 e4 e2 de e3 e5 eb f3 e9 f3 f1 f9 f7 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f4 f9 f8 fa fa f5 f6 f0 e5 f0 e6 e9 df d1 d0 c8 c8 c2 ca b8 c1 c4 bc ba c2 bf c8 c2 c4 c6 c9 d2 cd d4 cb ca c9 c6 c0 c3 bd ba bd bc bb ae b5 aa aa a0 9d 8d 85 7f 74 6d 76 76 77 6f 6f 6a 84 84 7d 54 45 34 15 11 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 06 0c 14 1e 30 4d 76 91 95 87 8a 81 80 83 81 85 85 8d 91 93 90 8b 91 91 98 93 97 a0 9f a5 a4 9f a4 ae a8 b0 b8 ba bf bd be c3 d4 cc d6 d5 e0 d5 e1 e0 e3 ed e9 e8 e9 e6 e7 f3 f1 f5 f6 f7 fd fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f8 f5 f3 ed e8 e2 e1 e0 e0 da d7 da d4 cf cb c0 c5 c0 c0 bc ba bc bf bc c4 bb c8 c2 c4 ce d0 cc cd cf cd ca cb c8 c9 c6 c0 bc b7 b8 b8 b6 b2 a7 a7 9a 94 8d 7b 7b 76 74 72 67 6d 71 6d 71 82 7f 74 53 49 26 1a 0f 05 09 06 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 09 03 0d 06 11 1e 20 2d 49 65 84 8f 87 7f 83 82 80 88 8c 8e 90 8b 8f 94 94 97 91 96 96 93 98 98 9c a7 a2 b0 ae b3 b0 bf bc bb c6 c7 c2
 c9 cd d4 d7 d3 e4 d8 e2 e3 e6 e3 e8 e3 eb ee ec ed ef f4 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f7 ec e3 e0 e7 df e9 e8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fb f4 f0 f0 f2 e9 e6 de db e0 d8 d4 cb d3 cf c6 c7 c4 bd bb be bd b9 bb b9 bb b7 bd bc c0 c6 ce cd ca c7 d2 c8 cc c1 bd c0 ba c0 b6 b7 b3 b8 b4 ae 9f 9d 95 90 8a 82 7f 7a 77 79 7a 73 72 6e 75 7c 89 74 5e 45 2a 10 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 08 03 0a 06 0c 1a 1e 31 3e 67 77 83 8a 85 86 84 7d 80 88 8f 91 90 8e 8e 90 9b 94 92 94 96 9d 9e a3 9c a6 a7 b5 b5 b3 bb be c2 c6 ca c9 ca cc d8 d0 df d8 dd e1 e8 e1 e7 e5 eb e5 e4 ee f0 f5 f3 f8 f7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe e1 ca ca c7 bf c5 b9 b0 b9 b5 b1 bb d1 e3 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fe f9 fb f1 ec eb e6 db e1 d3 d7 d6 c7 d4 c6 be c5 c1 be bd c2 bb bd bd b1 bd b4 b6 be bf bf c8 bd ca c9 d0 c5 c9 c5 c7 c3 c1 be c0 b2 b1 b4 a5 ac a3 a1 91 81 89 82 85 7e 7c 7d 77 71 76 6c 70 88 89 70 62 4a 2a 19 0a 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 06 05 09 00 08 13 1b 1a 27 3f 54 6e 7d 84 7e 89 8a 86 8a 86 8c 89 8f 98 8d 8f 95 9a 96 94 95 90 94 a1 a1 a3 b1 ac b1 ae b8 be b9 be ca ce d1 cd d5 da de dc e3 e0 e2 ed df e4 e9 ec ee ef f4 fa f9 fa f6 fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 c5 ab af a7 a6 ab a2 95 96 97 98 99 a4 a0 b3 c8 d6 de f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f5 f5 f4 eb e9 e4 e9 e7 e0 db d0 ca cf d5 be c3 c0 ba bb bf bd bb be b3 bb b5 b4 b7 b8 c1 bb c6 c0 bd c1 bf bf c5 bd be bd b4 c0 b2 b2 b4 af ad aa 96 a0 9b 8c 89 80 80 7d 7f 81 78 78 6a 7d 7d 8b 8e 7b 59 3f 2e 1a 0f 05 04 04 06 0a 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0b 15 21 25 3b 4e 72 7f 7d 81 7d 86 81 84 8d 8c 8f 92 8f 94 97 94 8e 9a 9c 92 9a 9e 96 a6 9e ae ab aa b1 af bc c1 c1 bf cb
 cb cd d4 d4 da df db de e3 df e3 e8 ea ee ee ee f1 ee fb f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 cf b8 ad 92 99 8b 96 92 91 8e 8d 84 84 79 85 8b 98 a7 b2 be d2 e0 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff ff fd fd ff f8 f1 ed f1 e7 eb e2 e4 e1 e0 de d7 d4 c4 ce c1 be bf b3 be ba b7 bc b7 b0 b6 b3 b4 b4 b4 bb b1 b4 bb be bb c2 c3 c3 b9 b8 b8 b4 b7 bb ae b5 b1 a6 a0 a2 99 90 87 87 7e 7b 7e 7f 73 74 77 74 75 82 92 8d 74 55 3b 25 1c 08 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0a 06 0a 1a 19 26 3b 4c 69 7a 7b 7d 80 85 8b 81 85 8b 91 90 98 92 90 98 98 96 9a a0 9f 9f a5 a5 a6 af a5 ae af b9 bb bf bd c6 c6 cd d1 cf d5 db d9 df df e0 e2 e7 e6 eb e7 ea f5 f6 f4 fe fc f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 d2 b1 a2 96 8e 8c 80 81 77 71 79 78 74 7b 73 79 80 86 8a 8f 99 ae bf ce e8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff fc fb fe ff f7 f3 ff f5 f5 f2 f0 f4 eb e3 e2 e6 e1 d3 d3 cf c9 c4 ca c4 c0 bb bc b2 b5 bf b9 b2 b9 b2 b0 ae ae b6 b0 b6 b8 ba b8 c3 b5 be ba bb bf b5 bb af ae a5 ab a7 a3 a2 9c 90 8b 86 88 80 83 81 73 71 76 79 7b 85 95 8a 73 5e 48 24 1d 0f 05 03 09 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 06 05 03 05 06 0e 13 1c 29 33 49 6a 71 81 72 78 86 85 84 8a 8d 89 97 96 8f 94 95 99 95 98 9b 9c a3 9f a5 a8 a3 a7 b0 b3 b6 c1 b9 bb bd c2 cd d0 d0 d4 d5 dd dc d6 dd e2 e1 e6 e9 f0 ee f5 f0 ed f9 fa f4 f8 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 c9 a8 98 85 83 78 75 73 6b 61 63 65 69 69 64 63 65 6a 6d 7b 7f 83 94 99 ad c9 e4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 fc fa f3 f3 f2 f8 f1 f5 f2 ec f0 ea ef ee e9 e9 e4 e0 da d5 cf cc d0 c6 c1 bf bb bd be b4 bb b0 af b4 ad ab ae b0 b4 ae b3 bf b1 af b8 b9 bb b1 b4 b8 b3 b5 b5 ae aa a3 a2 9c 9a 95 96 94 84 8b 8a 87 83 7f 6f 76 7c 82 8a 9c 8b 74 55 38 29 17 0b 05 08 04 06 06 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 0c 1c 25 37 51 60 74 6c 75 74 73 7b 84 8d 86 8c 8f 90 93 90 9c 99 a0 9c 98 a0 a5 a4 ad a5 a5 b0 b2 ad b3 b7 bd be c0 c4
 d0 c9 d4 cf cf db d6 de e3 e2 e9 eb ef eb f0 f4 f2 f1 f9 f5 f3 fc fd ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 c9 ab 92 84 7f 72 66 60 60 5e 5a 56 53 56 57 5b 48 54 5b 5a 65 6b 6a 74 85 90 a0 c7 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f8 f7 fc f2 f0 f7 f3 ef ef f2 f4 ef f4 ed ed ec ea e4 e4 df e2 e1 d9 d2 d7 d3 cc c2 c0 bc b2 b8 b6 ac bc b5 a8 af ac ac a8 ad b3 ab ad b0 aa af ac b1 b9 b7 b4 b1 a6 aa b0 a5 a9 a0 9d 9f 93 99 8a 8d 8f 8e 87 75 80 7a 77 6f 7d 81 8d 96 84 70 5a 44 30 19 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 08 10 17 30 3a 4d 61 70 6d 70 73 74 7f 85 89 86 8b 91 91 9a 94 9c 9e 9b a0 9b 9e a3 9c a6 a9 a7 ab b4 ae b5 c2 b9 c3 cb c7 cd cd d3 d5 d5 d9 df e1 e3 df e8 ed e6 ec ea f2 fa ee f7 f5 f5 f9 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 bf a9 9d 8e 77 6f 5b 59 50 46 46 49 46 3b 4d 45 47 4c 48 49 51 58 66 6d 6d 70 7c 86 a9 ce ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f8 fb f5 f3 ef ec f5 ee ef ed ed e7 f0 f3 ea ea e9 e1 e0 e3 da e0 d2 c7 d4 d1 c2 ca bf bb b2 b8 bc b0 b1 ad a6 ab ac ab a9 ac 9f a9 b0 a6 ae af a6 b0 a8 af ae a9 ab a8 a5 a3 9f 97 9a 93 91 95 8c 90 85 7e 85 76 76 76 7b 84 7f 97 9e 89 75 5e 40 34 1a 0d 05 03 03 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0a 07 00 07 06 12 19 2c 36 4c 5f 6c 6f 66 6c 74 74 7f 82 86 89 94 96 98 93 9c 9e 9e 9f a1 a3 a6 ab aa ae a3 a7 a6 ad b3 bc be c1 c2 c5 d2 ce d3 d3 d8 d8 db e0 e2 e2 e3 e9 e9 f1 ed ea ee e9 f3 f3 f2 f1 f9 fa f6 fa ff f5 fe ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 cd af 96 87 75 5d 5c 4a 4c 46 3d 42 40 46 40 3f 3e 44 3a 49 48 4d 48 52 57 61 65 76 85 9f af cc f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f5 ef f0 f3 ee f0 f3 f6 e4 f0 e4 da e2 e5 e2 e9 e3 e7 e3 e0 dc d9 d7 ce d2 c6 c2 c1 be ba bb b4 b0 b0 ac ae ab a4 ad a5 ac af ad b7 ab a5 a7 af a6 b0 ab a9 a6 ab a4 a7 9b 9e 99 9d 92 93 93 84 87 8a 7c 7d 81 78 79 7b 7d 7f 94 9f 8b 78 5a 3e 22 19 13 05 03 05 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 10 06 07 14 17 25 34 4b 60 66 69 65 62 70 6b 75 79 80 8a 93 93 95 97 95 9b a1 a0 a6 ad a4 a7 aa ae ae ab ab b0 b6 b7 b6 b6 c2 b9
 ce cd c7 cf d5 d8 dd db dc e3 e0 dc e3 e8 e6 e7 f1 ed eb eb f3 f0 f6 f5 ff ff f5 fc fb fa fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff db b5 98 8b 71 62 52 51 4b 3f 40 38 3d 35 3a 38 3e 3a 3c 38 3d 3f 45 4b 3b 45 49 59 68 78 80 9a ab d9 fe ff ff ff ff ff ff ff ff ff ff ff fa fe f2 fa eb ea f1 ed e6 e7 e8 e6 e7 e9 e7 e6 e0 dc e1 df e5 e4 e2 de dd d6 d5 df ce d1 c4 c0 c0 bd b9 ba b0 b1 ad ad af ac a6 a8 a8 a3 a9 a1 a1 a2 a1 a7 96 a1 9f a7 a4 9f a2 a0 96 99 9c 9b 97 95 8b 90 8b 89 89 82 7a 73 73 78 75 7a 7d 95 9c 85 6d 58 33 24 13 09 05 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0a 06 0d 0f 22 23 35 47 61 6c 72 67 5d 64 70 72 7d 82 83 8c 93 95 9a 9a a2 a2 a3 9c aa a4 ac a3 aa ab ac b3 b1 b3 b6 b6 bd cd c7 ca c8 cb c9 d4 d4 d2 d8 de d9 db e6 e2 e3 e6 ec ed f1 e5 f0 e6 ef f7 f2 fb f5 f3 f5 fd fb ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c4 a6 8c 71 5d 4c 50 42 38 36 3f 3e 37 31 34 33 2f 30 2d 36 36 3f 37 38 41 45 48 52 51 64 73 83 9b bf e7 ff ff ff ff ff ff ff ff ff ff ff ff f5 f5 ed f1 ef ea ed e4 e3 e6 e1 de dc ed e5 e3 da da da db e4 e5 de e4 da d4 d2 ca d1 c4 c0 bd bc b4 b2 ae b5 ae a9 b1 ab b3 a8 ad a7 a0 a4 9d 9f a0 a0 a3 a7 96 9c 9c 9b 9e 97 9b 9e 99 93 96 9b 90 89 8c 81 80 80 7c 73 7b 77 7f 76 7d 8d 9d 82 73 54 38 25 1e 08 05 06 00 06 06 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0b 05 03 08 07 0d 13 13 2b 34 49 61 73 6c 5f 63 66 65 6f 7a 78 85 8a 91 94 8f 95 9b 9a a5 ab a9 ae ae ae ae b8 b4 b0 b3 b9 b9 b3 c3 c1 c0 c1 c5 ce cd d1 d5 da e1 de db e3 e1 e0 e3 e6 e4 e8 ef f0 f1 ee f0 f6 f2 f4 ee f6 f7 fc f8 f8 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 b6 95 7c 65 5c 3b 3f 3c 3a 3d 38 30 32 31 34 31 31 2d 2c 33 2f 30 34 33 31 3d 4d 52 4d 56 65 77 82 ae e0 ff ff ff ff ff ff ff ff ff ff ff f9 f8 f4 ee ed e8 eb e6 e8 e1 dd dd de e6 e2 e2 d9 df da e0 e5 de e4 dd da e1 d6 cc d5 d3 c6 c1 c4 bb b8 ad aa a9 af af aa ab a9 a8 a6 a0 a4 a6 a5 97 a5 9a 9a 9d a0 a0 9d a3 96 97 99 9a 93 98 90 8a 8e 90 88 83 7f 85 7f 7d 7b 7e 76 74 7d 92 9f 8c 6f 56 3a 2f 11 08 05 04 06 06 05 06 02 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 1a 1e 22 35 49 66 68 6a 67 64 62 62 6e 6d 76 76 82 8b 90 8d 99 96 9b a5 a7 a4 af af a6 a7 b6 b0 b4 b6 b5 ba be b9 c1 c3
 ca c5 c8 ce d1 d0 ce d9 d7 e0 e2 e8 e0 e6 e1 e8 ea e4 e6 ec f0 ea ee f5 f2 ea f4 f7 f5 f6 fe f2 fa f8 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d5 a3 83 66 59 47 3d 37 2c 34 27 29 27 2a 22 2b 28 1f 21 2a 24 29 2f 24 33 36 38 3c 3c 41 48 5c 65 72 9b cd ff ff ff ff ff ff ff ff fd fc f6 fc f8 f4 ef e7 e9 df e0 e8 df de db d4 e2 e1 e4 d7 e2 f0 e4 e6 d4 db db da d6 d9 d2 d2 cf c6 c2 bc c0 bb b1 b2 b2 af ae a8 a8 a6 a4 a4 9d 9b 9d 97 95 97 9d 9e 94 98 98 98 9c 91 98 93 94 8e 93 95 88 8e 84 87 88 89 7f 81 7b 7b 77 72 74 76 82 9c 87 6f 55 37 22 0f 19 05 03 09 06 05 06 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 07 14 11 2a 39 43 60 65 65 66 5c 61 68 69 74 76 7a 83 84 89 91 93 95 9b 9e a5 a9 a9 af b4 af b3 b2 b4 b1 b6 c5 b5 bb c1 ba c4 c1 c5 cb d1 cf da df de db e2 dc e5 e0 e5 e9 e6 e4 e5 ea f0 ec ea e3 f1 f1 ea f1 ed ef ee f5 f7 f4 f7 fa fb f8 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff c8 a3 7b 5e 4d 45 36 2e 2a 31 25 25 23 1b 1e 21 1f 1f 1c 1f 19 1e 1c 24 23 27 2c 25 3c 3e 41 47 54 61 82 c5 fc ff ff ff ff ff ff ff fe f9 f5 ef f6 f2 eb ed e2 e9 dc e3 d9 d8 d8 dd de d8 d9 de e8 f5 f3 ef e0 d8 dd d9 d1 d2 d5 d5 d0 c4 c8 b5 ba b8 ae b0 aa b0 aa aa a9 aa a4 9b 9d 91 9a 99 9d 9f 9e 9a 91 a3 8f 9b 90 97 9b 95 9d 91 90 91 8f 8c 88 83 87 7a 80 83 7b 7a 7b 79 6b 6e 7b 8b 81 6f 4f 35 22 19 0d 05 0b 07 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 01 0b 0a 0f 1f 25 30 4b 5c 69 6d 67 5f 66 64 68 6b 73 6d 7d 85 88 8d 8e 93 99 9d 9d a2 a6 ae b0 a8 ad af b3 b3 b0 be b6 b3 bb bf c1 c0 ce d0 c9 d0 d2 de e7 dd df de de d9 e5 e8 ee e6 e7 e7 e9 e1 e9 eb e9 ec ed eb ef f2 f1 f0 f5 f1 f2 f7 fc f4 fd fb ff ff ff fb ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff bf 85 6d 54 3e 43 39 30 29 1e 1d 1e 21 20 16 17 1d 1e 19 22 1c 1a 1a 23 21 29 2d 39 32 37 35 46 47 58 7d b5 ec ff ff ff ff fe ff fb f5 f5 f0 fb ed ec ec e1 e2 e2 e3 e0 df db d9 d6 d7 d6 d6 e0 e8 eb f6 f0 e4 d3 ce d4 c5 cb cd c6 d2 c1 b8 be bd b3 ae b4 ad a9 ab a7 a2 a7 a5 a0 a0 96 9f 98 95 9a 8f 95 98 94 99 a2 91 a0 94 94 97 9b 98 90 86 8d 89 8b 8a 7f 84 84 80 78 78 77 76 6f 77 89 7a 72 4f 35 27 14 18 0d 05 0c 06 05 03 02 06 05 03 02 06 05 05 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 12 1b 20 3e 4d 5c 6c 67 62 60 66 66 67 6e 70 75 7b 7e 81 86 8e 96 99 9a a2 a0 a1 a7 a8 b0 b1 ae b0 b7 b2 b9 b3 b6 b8 c0
 be bc c2 c7 c7 d3 d7 d2 db db e0 dd e2 df dd e1 df de e9 e8 e4 e2 e3 e3 ea ea f2 e5 ec ec e0 ea f0 ef e6 f0 ea ef ef f5 ff f8 fd f9 ff f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff bd 85 66 50 3a 34 25 23 22 1d 1a 1a 13 20 1b 08 1a 0e 11 10 16 1b 10 13 18 21 1d 30 2c 28 2d 39 4c 4d 6c 9a de ff ff ff f8 ff f3 f4 ef f8 f2 eb f2 ea e4 e4 e1 d8 d9 da d8 d5 d0 d6 d7 d2 cf d5 da ea f2 f7 e9 d9 cf ce ce ce ce cc c7 c7 c7 ba b1 b6 b1 b3 b3 ad a5 b0 9c a6 9c a2 a8 99 93 91 92 98 92 8e 95 95 96 97 97 91 95 93 91 90 96 89 90 89 89 86 8c 84 84 88 7f 78 74 6c 6d 6e 75 84 7a 6c 51 35 1a 19 11 05 03 01 06 0b 03 02 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 10 12 19 21 36 45 55 72 6d 63 65 61 64 67 68 67 69 77 79 79 84 8b 8b 92 99 9e 9d a6 a4 a0 ab ae b1 ae aa a8 af b7 ab b2 ba ba b7 c1 c3 c5 cb d6 cd d4 d2 de e0 da e1 e1 e0 e0 e0 e5 e4 e3 df e3 e5 ea dc e3 e5 e8 df e5 ea e1 e4 e3 f0 ee ee e9 f1 f1 ea ef ed fe f4 f9 f7 ff fd fe fe f7 fa fe fc fd fe ff ff fc ff ff ff fe ff ff ff b1 79 60 46 31 27 2a 1b 1a 13 17 12 14 15 14 11 0f 10 11 0f 0e 12 15 15 1b 13 1b 1f 27 22 28 31 45 5f 67 9a df ff ff ff f1 f0 f1 f5 f1 f4 ee e5 e6 dc e6 db db dd d6 d8 de cb d0 c9 c9 cf d1 d4 d5 dc eb f0 ec e1 ce ce ca ca c6 cd cd c1 c1 bf b4 b3 b3 af a4 a4 ab a5 a7 9e 9a a0 9e 94 9a 98 91 8e 90 8f 90 8f 8f 8c 91 94 8f 8d 8c 90 8b 90 8f 88 7f 84 86 82 86 7d 6e 70 6e 75 6d 5e 6d 75 78 68 43 2f 24 0e 15 0b 05 08 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 06 0c 0a 1a 2b 2e 48 59 6c 74 63 62 5d 66 68 6c 67 6c 66 79 7a 82 8a 8f 91 96 9c 9c a0 a8 ab a6 a9 ac b3 ae a8 aa af b0 b8 bf bc ba ba c2 c8 c9 c3 d0 d0 d5 da e0 da de de e0 e6 e3 d7 dc df e2 e2 df e7 e2 de e2 df d9 e1 e4 e2 e4 e6 eb e6 e0 ea ea f5 ee ed e9 f7 fd f4 f9 fc f2 f8 f7 f4 f0 f1 fa ef f8 f4 f1 f4 fc fb fa ff ff ff ff ad 74 5e 49 34 1e 18 11 13 13 17 1a 13 10 16 0f 12 13 12 09 0f 12 14 16 0d 0a 15 21 26 26 2f 28 3d 51 65 95 da f8 fd fd ed f0 eb ed e6 e4 ed e3 d7 db d6 d9 d7 d2 cf da c5 c8 ce cf cb c7 d1 c5 cb d5 e2 f1 f0 e6 d0 c9 c8 bb c2 c3 c1 c5 c4 bb be af ab af b3 aa a9 aa a1 a2 9c 9b a2 98 96 8d 94 90 9c 98 8e 93 8b 92 8e 93 92 94 92 91 7a 8d 85 85 8a 83 83 88 82 7c 77 6e 6b 6e 67 62 69 75 75 66 47 32 26 1d 10 06 03 00 06 05 03 01 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 07 08 0c 12 14 21 35 4a 65 6c 74 6b 66 65 62 62 6b 68 72 73 70 75 7d 80 8a 8a 96 9c 9a a3 9e a6 a5 9f ac ae a4 ad b5 b0 b1 b2 b9
 b8 ba c1 bf c4 c3 c4 ca d5 d6 d9 da d9 da d9 da d9 db da e1 df df e1 db db e0 da d5 dc d9 db dd df e3 e2 e4 db e1 e6 df ed e5 eb f0 ee ef f3 e7 f2 e5 ef f5 ec ee f0 ea f0 f3 ed f0 f1 f0 f3 f1 f2 fd ff ff b8 76 5b 47 25 20 1d 14 19 10 0e 17 0b 0b 0c 0b 0d 1a 14 13 0b 0d 09 0f 19 19 16 20 1d 20 22 29 35 50 69 8d d8 f0 f1 ee ea e4 e9 e4 e3 e5 da de de d4 df d3 d3 cd d0 cd c6 c9 c6 ce be ca c6 c9 ce d2 d8 e6 ef ed d7 c4 c2 b2 c1 c8 c5 bd c2 bb bb ae b8 a9 ac a8 a8 a0 a5 a4 9a a3 9a 95 99 92 8c 92 8d 8e 8f 98 8e 8e 8d 93 91 93 91 95 8f 91 86 8b 85 87 8a 80 81 7e 78 78 6e 6a 6b 61 64 6f 6b 61 4b 42 27 17 10 06 09 04 06 05 03 00 06 05 03 07 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 0b 14 18 2f 34 46 52 6b 71 66 6b 66 64 67 60 66 67 73 6e 73 80 78 7e 87 89 97 94 94 9f 9e 9f a9 a6 a7 a2 9d a8 a8 ad af b3 ae af b2 b8 bc bd c1 c2 bc c6 c8 d5 c9 d2 dd d4 d8 d8 d5 d9 da d7 d7 da dc d4 dd d9 d7 db dc d8 e5 d6 d6 d5 d8 d9 e1 e6 e3 ec e7 e4 e9 f1 e9 eb ee ea df e7 e1 ea e0 ec e8 e4 e6 ec e9 fb ef f4 fa f4 ff ff b8 6f 5b 47 20 1a 15 09 09 10 0a 0d 0a 04 0d 0f 0a 0a 06 0e 0a 11 08 06 10 09 0f 0a 17 1c 1f 2a 31 46 68 94 d3 e3 ec ed e5 dd e0 df db de db dc d2 d3 cb cc cc cb c9 c9 c1 c2 c5 c5 c8 c8 c1 c8 c9 cf d6 d4 e5 e2 e0 ce bb b4 ba ba bf bf bc c0 b1 ad a8 b3 af a5 a2 97 9e a0 9d 9f 99 94 9b 8c 8e 87 90 91 91 95 8d 94 90 85 8e 87 8b 90 91 8f 8f 8b 87 89 83 78 80 72 77 6b 71 67 6d 60 61 62 69 6a 4b 3d 23 17 12 08 03 00 07 05 06 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 07 0e 0b 15 1d 21 2f 42 5c 6d 7f 6d 6f 6c 68 60 64 6a 71 71 7c 6f 74 73 80 82 8f 8c 95 99 9d 9d 9d 9e 9e ab a7 a1 ab a5 ad ad ab b7 b3 ae b6 b8 b9 c0 c3 c4 cd c7 cb cd d0 d4 d1 dc d7 cc d7 d4 d0 d5 d5 da d6 cf db d7 da d9 d6 dc d0 d7 da de d8 e0 de e0 ea dc e1 e3 dd eb e5 e2 e8 e1 e2 de df de e0 df e1 e9 de e3 e9 e9 ee f9 f5 f3 ff cb 76 5c 4e 21 17 13 06 12 12 12 09 08 03 0c 0d 09 0a 0b 05 0a 0d 12 0e 08 0f 13 0e 16 1e 17 26 28 4b 74 9a d8 e4 e3 e5 d9 dd de dd db d0 d4 cd cd c9 d0 d0 c8 cc c4 bd cc bb c3 c5 c7 cb bf c8 cd c5 c9 d1 dd df d5 cc bd b8 b8 bc ca c1 ba bf b0 b0 b3 b3 aa ae aa a5 a2 9f 9f 9a 94 90 90 95 90 8f 91 93 8d 8f 8f 8e 94 90 92 88 8a 88 8b 8e 8d 88 84 86 84 7d 77 7b 78 6f 75 6a 63 5f 64 64 69 61 4c 3f 2a 20 16 07 07 00 06 05 03 04 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 07 0a 0e 1b 24 37 42 60 66 74 7a 67 65 64 60 6e 67 6e 71 74 7d 71 6f 7a 85 85 92 90 94 9f 98 9a 9d a1 a7 9f a7 a9 9f a8 b0 a9
 b3 b1 b2 b1 b7 b4 bb ba bb cb bf c5 cc d2 d1 d3 cc d6 cd d3 cf d3 d4 d3 d5 ce d0 d3 d0 cd d6 d9 cd d7 d3 d7 da d8 d7 da e4 d8 e2 df de e0 d9 da de e0 d5 d4 da d7 d5 de db d8 e0 da e3 ea ea f7 f4 f0 ee f5 d0 7d 61 42 23 19 0b 05 04 12 14 09 06 00 06 0b 0e 04 0a 07 04 05 06 0e 08 0e 13 13 1a 12 18 24 2c 4f 84 b7 d1 d8 d8 d6 d6 da d8 d5 ce d8 ce d0 d2 cd c7 d0 c6 ce c8 c3 bf be bd c1 c0 be bf c4 cb ca c8 c4 cc ce cb c4 b6 b9 b6 bc bf b4 bd bd ac b0 b2 ae af ab a4 a8 a6 a0 a0 9b 9c 98 93 93 8e 89 95 8a 89 8a 8f 9b 90 89 8c 8d 8f 8d 87 8a 89 82 81 89 82 76 78 70 6d 6f 6a 68 6c 69 64 62 6d 66 56 39 32 13 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 12 1b 27 34 48 51 6d 74 79 63 6a 6b 60 69 68 69 77 76 7e 75 73 72 77 84 8b 8f 93 92 95 99 95 98 96 9d a0 9c a1 99 a8 a1 ab af b4 ae ac af b6 b6 c0 c4 bd c4 cd c8 cd cd c5 cd cb c9 c3 ce cd d3 cd cb cc cb c5 ca d1 cd d2 d0 cd d5 d4 d3 d6 d5 d4 db d6 d9 d6 d8 d6 da d8 d2 ce d0 cc cf d6 d7 de d0 db da dc e2 e1 e7 ea e3 d5 e3 d7 89 63 3b 22 0e 06 05 0b 09 06 0c 08 02 08 05 03 00 06 05 06 0c 06 05 0a 10 09 12 16 12 1a 18 1f 45 8b bc cf d9 ca d1 c5 d0 d5 d3 cb cd c6 c7 c9 c9 be be c8 c1 c1 c3 b6 b6 bb b2 b8 bc ba c8 d0 c9 c3 c3 c0 bd be b7 b7 b2 b5 b7 b1 b7 b0 b2 b5 b1 a5 ad a7 a9 a7 a5 9b 97 91 a3 94 96 99 8c 8c 8d 8a 8f 91 91 90 91 85 85 89 84 8e 88 87 94 83 87 86 7b 76 76 71 70 73 68 76 69 6d 69 65 70 63 65 5b 40 27 1a 17 05 08 02 06 05 08 00 06 07 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 0e 1b 25 2e 43 5c 6d 7a 73 68 63 65 6a 65 6a 68 76 74 7b 7b 7a 72 78 79 83 85 8a 94 8c 95 96 9c a1 a0 a4 a2 9b 9f a1 a5 a5 a2 a5 ad ac b5 b3 b6 b2 b4 bc ba c0 c4 c3 c2 c5 c5 d0 d2 c7 ca cd c3 d5 c8 cb cc cb c9 c4 cc c6 c9 d3 cc d3 d0 ce d6 d6 d5 db d7 d3 cf cf d1 cd c3 c8 ca c9 cb ce cb d2 d7 d2 d6 d0 dc e7 e7 d8 d3 c9 c6 cd a0 6b 43 19 0b 06 09 0c 0b 0b 0d 0b 09 0c 08 0d 05 06 06 0a 09 06 0d 08 0e 11 10 0b 0e 14 1e 25 48 91 be ca ce c4 ca c9 c6 c4 c0 ca c9 c0 c1 c0 c4 c0 c6 be bb b1 bd c2 b1 b6 b7 b4 b1 af bf bf ca c5 c1 be b8 b6 b7 b4 a6 aa b4 ad aa b5 ad a7 ad b6 a8 b1 b0 a7 a2 9a 9f a6 95 94 8e 8e 8e 8f 90 93 90 87 8e 93 93 92 8a 96 85 90 8a 8d 8a 87 88 84 84 79 78 68 68 69 70 71 6d 6c 64 6b 65 67 6a 51 48 33 1f 17 05 07 06 06 05 03 00 06 05 03 00 06 05 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 04 06 05 03 06 06 10 10 16 25 38 42 5b 6f 7c 70 70 69 6a 6b 69 72 69 6b 7c 7b 7c 7c 7a 7f 83 86 83 8a 8c 8c 90 94 9a 98 9c a4 a0 a7 99 a0 a4
 a4 a4 a8 ac b3 a5 b3 ab b2 b1 b7 b8 b8 c2 b6 c1 c0 c6 d0 c5 c6 ce cd c1 c6 c6 c3 c3 c7 d0 c2 cd ca c7 c8 d1 cd d0 d6 d5 d7 d2 d9 ce ce cd ce cc cf bd c4 c5 c4 d0 d0 db d6 cd ce cd c5 d1 de dd cb ca c6 b4 bb a9 75 41 16 09 07 09 09 08 06 0c 0d 06 07 0a 05 07 09 08 07 03 06 0d 12 04 13 13 0f 12 10 1c 20 3c 8e bf c3 c8 be c4 c2 bd c3 c3 c3 c3 b9 b9 c4 c5 c0 c0 b9 bb b9 bd bb b6 b2 b2 b9 ae b9 bc c5 c7 c9 c0 bb ba b6 b3 ac ac a9 b0 b1 b5 b1 b5 af ac b4 ab b1 ab a0 a3 9e a8 a3 a1 9e 94 95 93 91 8b 90 95 85 9a 8e 93 94 94 89 93 8e 92 89 8a 87 87 78 71 6d 70 6c 6b 6a 67 75 68 6a 64 61 64 6e 68 60 4e 3b 22 0b 0e 07 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 04 06 05 0e 13 1f 2f 3f 54 6e 70 71 6d 5e 64 67 64 69 6d 6b 6d 72 72 6d 71 7e 83 8a 83 85 84 87 8d 8d 91 95 92 9f 9b 94 9f 9a 9e a3 a3 a9 a5 a5 a9 a7 ab b8 ae b6 b4 b3 b1 b3 c1 b9 c0 be c3 be c5 c5 be c0 bb c1 c2 ca c0 bd c3 c6 c6 c6 c5 ce c2 c4 d0 ce ce d2 d0 cd c4 d0 cd c1 bf be c3 bd ce cb c5 c4 bd c1 bf cf d6 d6 cb c9 c7 ba b4 ab a0 70 3f 1f 10 0a 07 03 0c 0b 05 09 06 06 08 09 01 06 05 05 00 07 05 05 0f 06 12 11 10 13 18 1b 41 97 b8 be c2 bb bc b7 b6 b7 b9 b3 bb b7 b6 ba b2 bc bc bd b6 b3 ba b6 b2 b3 b2 b4 b1 b6 b0 bb c9 c8 be b2 b3 b0 a5 a1 a8 9f a8 a8 a5 a6 ae a5 aa ae a8 ad ab a9 a6 a4 9e a7 99 9b 9a 92 90 8f 94 90 87 92 90 9a 9a 8e 99 8a 95 93 8b 94 86 7e 7d 78 76 6e 69 6f 6f 6c 69 69 6f 6b 67 5f 65 69 68 5d 47 3a 21 1d 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 07 14 19 29 31 46 55 6e 7b 74 6f 61 66 69 6c 70 6a 6d 70 6d 80 73 78 7d 7c 80 7d 88 88 87 8d 94 95 97 94 9a 9a 99 9f a0 9c a1 a1 a3 9d ac aa a4 a7 aa ac af ae aa b0 ae b6 b6 b9 be bf bd c0 c4 c2 bb b9 bb c1 b7 b7 be c6 c8 c3 c6 ca c5 c8 c5 d0 cb ca c2 c7 c1 c5 cd cd ca b9 bb c2 c4 c6 c6 c9 bd bf c1 c9 cc cb c5 ba ba b7 ad b1 a4 9d 7c 4c 1f 10 06 05 05 09 0a 0f 08 04 06 05 07 01 0b 06 03 08 06 05 04 10 09 0c 18 12 15 16 20 3e 88 b3 b7 bc b2 b7 ad b9 b5 b2 af ae b0 b9 b2 b6 b2 b8 b4 b3 b1 b3 b4 b1 b5 b3 a8 ad a9 aa b8 bd be be b3 ad b0 a6 a5 a2 a6 aa b0 a0 a3 ad a4 a1 ac aa af ac a5 a6 9a a1 99 a1 9b 95 9a 93 90 90 92 93 93 92 91 95 97 99 99 94 96 8f 8a 81 7c 78 72 6c 6b 6f 66 6c 67 64 6e 6f 6a 5f 67 5d 61 6d 5a 53 39 26 19 15 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0f 11 1f 1d 2b 4b 57 64 7b 79 60 69 61 66 6d 72 6d 6f 72 6f 74 7c 7d 83 84 83 7e 89 86 88 83 91 94 95 96 95 9d 98 95 9d 9e
 9e a1 a0 a1 a8 a0 a5 af a5 ad ad a7 ac b2 b6 b7 b8 b3 be bc be b6 b4 b8 b8 b5 bd b7 b1 bd b6 c0 bf b7 c1 c4 c3 c8 c4 c4 c7 c6 c1 c4 c7 c4 c1 c5 c1 bf be bd be c2 c6 bc ba b9 bd c8 c5 c9 ba b8 b7 b0 ad ab a7 9a 76 4a 23 0f 06 07 05 0b 0f 05 03 06 06 06 09 05 06 05 0a 0a 06 05 03 08 06 08 10 14 1a 17 22 3b 77 ab ad b2 aa b7 a8 b2 b3 a7 b2 ac b2 ac b4 b0 b1 b7 b0 ab b0 b2 aa ab a8 a7 a3 a7 a8 a6 a9 b6 ba c2 b2 af a5 a4 a1 a0 a6 a2 ad 9d 9e a1 9c aa a0 a5 a6 a8 aa a5 a1 a7 a0 a3 9c 9c 97 9d 8e 97 96 9b 94 9a 92 99 90 98 9a 95 88 84 85 87 7b 75 71 6d 71 6b 68 6a 73 6d 77 64 61 5e 5e 6d 6a 6e 5c 58 44 2f 21 12 0d 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 05 12 1a 25 2f 46 56 60 74 71 6e 67 64 61 69 6c 6d 72 6f 6a 75 78 7a 81 88 86 7e 85 86 88 8d 92 94 8b 8a 97 91 96 9c 99 96 9f 98 a8 9b a3 9f a8 a2 9e a2 9f a1 a9 a9 ab b3 ae ae bd b7 ba b0 b6 b0 b1 b5 ba b0 b8 b4 ba c5 bf c2 b9 c9 c7 c5 bd c0 c3 c4 ba c1 b7 c2 c2 cc c3 ba be be bd be c4 bc b5 b6 ba c1 ba bc b0 a8 b3 aa a4 a8 9a 99 70 4d 1d 10 06 05 11 06 09 09 06 04 06 05 03 07 06 05 05 00 06 05 05 06 0e 0c 10 0f 0a 19 1e 2c 7c 9c a8 b1 a8 b3 ac a1 a9 ae ac b2 a8 ae a6 ad b6 b0 ad ac a7 ac a6 ac a5 a7 a3 9f 9e a4 ab ae ab ad b1 a6 a6 a3 9b 9d a2 9a 9d 9e a0 a5 9d a1 a9 a6 a4 a6 a6 a1 a8 a0 9d a2 9d 9f 98 94 94 90 92 89 90 91 91 98 8e 8f 88 8e 7e 7f 81 73 70 71 6f 6b 66 66 66 6d 6a 65 6e 6b 61 5c 5f 62 6e 6e 65 55 40 2e 20 0a 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0b 25 30 39 47 4d 5d 6c 6c 5f 5a 64 5c 64 70 71 75 78 6d 72 6b 75 7b 7e 84 84 82 81 81 85 8e 8a 91 94 89 95 94 96 97 9b 96 9a 9b 99 a0 a9 a3 a4 a1 a1 a0 9d a7 a6 a9 b0 a7 b3 ab b5 a8 b3 b5 b2 b8 b2 ab b1 b1 b4 b2 ae be c0 bc bd bb b9 be b5 c4 c4 bb b7 bb b8 bc c4 c6 bc b7 b1 b6 bf ba b5 af ad b2 b4 af a9 af aa a3 a4 a3 a4 9d 98 79 57 23 10 06 05 09 06 06 09 04 03 06 05 07 01 06 05 03 05 06 05 03 09 0a 0e 06 06 0d 09 19 2f 77 a2 a5 a6 a2 a5 a3 a1 a1 a7 a4 a6 af ae 98 a5 aa a7 ab a2 a4 9e a4 99 9b a0 a0 9b 9b a0 a6 a7 ad ac ac af a4 9e 9c 9c a0 9e a0 9f 9b 99 98 a1 9c 9e 9f 99 a1 a5 9e a0 9d 9e 96 92 8d 97 8b 8f 96 94 8a 84 84 8c 8d 8f 85 82 79 79 75 71 6e 65 6d 69 6a 63 6b 69 67 6a 65 68 57 5f 5d 5e 6a 6d 6c 54 47 27 21 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 03 06 0a 0e 1a 2b 3a 49 57 6a 74 6a 5b 63 60 62 6b 68 79 72 78 78 75 7a 7a 7e 7d 81 8a 87 87 80 85 83 8c 92 94 97 9d 9b 9a 97 96
 9f 9b 98 a2 95 9d a5 9d a1 9d 9e a1 a1 a3 a2 ab b0 aa af ad ab ae b4 ae b2 aa aa ac b7 af b1 b5 bb b9 bf c8 c4 b3 b5 b4 c0 b7 b6 b2 b3 b6 b4 ba c4 b0 b6 b3 ba b1 b9 b5 a2 a1 a4 a7 a9 ad a1 a3 9e a4 a0 97 9b 90 7d 5b 21 0f 07 05 07 09 07 0b 03 00 06 05 04 07 06 06 05 02 06 05 03 05 06 0d 0f 10 12 11 1b 2f 71 9b a3 aa a0 a4 9f a8 a6 a5 a9 99 a0 a2 ac 9f a9 a2 a7 a2 9b a1 a2 9e 98 a5 97 9f a2 9d 9b 9f a8 a3 a9 a1 a1 97 9d 9c 9d 9b 99 9f a2 a4 a1 98 9b 97 9e 9b 93 a3 9b 9d 8f 97 97 97 95 91 8a 93 8d 86 89 8b 8d 90 83 85 83 7a 85 72 75 6f 69 70 6d 65 6e 66 66 6a 6e 6c 6b 5b 59 5f 60 5d 66 70 67 53 4a 33 20 17 06 05 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 05 16 20 24 44 40 59 68 68 62 60 62 5d 65 62 63 70 75 72 79 7b 70 7a 7d 82 83 86 85 8b 88 91 87 8e 8b 87 91 94 94 97 92 98 9e 9e 9d 99 95 99 98 a0 9a 9e a4 9d 9a a3 9d a6 ad a9 ac a2 a9 a3 aa a3 ae aa a9 b3 a5 af b2 b9 ba b9 b8 b5 b7 ad b6 b8 bc b6 b0 af b3 b0 b0 b5 ba b0 ad af b0 b4 aa a9 a0 a0 a6 a6 9e 9c 9a 9e 9f a2 a2 98 9b 90 86 5f 25 0e 06 05 04 09 06 05 03 04 06 06 03 00 06 05 06 00 06 05 03 04 0d 0c 03 07 11 1c 10 31 6c 99 9e ad a1 a5 a0 a2 9c 98 a1 a1 a1 a4 a2 a1 a3 a0 a0 95 98 9a 95 96 8b 9f 94 99 98 95 9f a2 a4 a9 a5 a7 a2 9a 93 95 96 98 9c 95 9d 9d 9c 99 9b 99 91 94 95 9d 90 92 8f 90 8b 8b 8d 89 89 87 86 88 8a 89 85 85 85 78 7b 73 77 69 66 72 62 68 6d 69 67 66 66 67 5d 5f 63 61 5f 56 5c 57 62 71 6a 57 4d 30 25 0b 05 01 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 19 24 2a 34 42 5a 5d 62 66 5e 61 5c 59 66 67 6c 73 73 82 73 7a 7e 7d 80 80 82 84 82 80 87 89 8c 8b 90 95 94 8e 99 98 9c 9b 95 9a 95 94 93 8d 9b 9e 98 93 9b 98 9b 9e a1 a5 a0 a2 a6 a1 a5 a4 ad af b0 a3 b3 ae ad b5 b5 b1 b5 b1 bb b2 b1 aa ad b6 a8 b0 a9 a5 af ad b5 af af a8 ae af a9 9e a6 9e 9f 99 a5 a3 a2 a4 98 a3 9d 94 a1 8d 8f 80 64 20 10 06 05 03 07 08 05 03 03 06 05 03 00 06 05 03 02 06 05 03 06 08 09 09 0f 13 14 1c 2b 6c 9d a1 a7 9e a2 9a a0 95 98 99 a3 9e a0 98 9e 9f a0 9d 94 95 96 99 96 93 94 91 8f 96 93 97 92 95 9c a1 a0 97 a0 98 91 95 89 9a 90 97 95 99 9c 9a 8f 8b 9b 93 92 8a 8f 8f 8d 90 82 8e 8a 85 86 81 84 83 85 83 7b 75 7a 71 6b 70 6c 73 6a 6e 6b 70 67 6d 62 66 62 5b 63 5e 56 56 51 56 5f 68 6f 66 5b 48 39 21 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 10 11 1d 33 3f 4a 5a 5b 5e 57 54 66 60 5e 64 5d 68 68 79 7d 7e 80 7e 75 7b 79 7f 84 80 8d 84 86 87 8f 89 8e 93 8e 97 8e 95
 95 92 92 97 95 96 9b 94 92 9b 9a 9b 9b 98 9a a0 98 91 98 a4 9c a0 a8 9a a9 a5 ad aa ad a6 ab b3 b1 b0 b1 a8 a7 ab a9 b4 b3 a7 aa ab a4 b2 a6 a9 b0 a2 a3 aa 9e a0 98 9a 92 a0 9e 9b 9f 9d 97 96 92 98 9e 95 94 94 81 60 2e 0d 06 05 03 0a 06 05 03 06 06 05 03 05 06 05 03 00 06 07 03 08 0a 07 08 07 11 0c 12 20 67 98 ab a8 9f a5 9f 9c 9a 97 99 9f 9a a1 94 98 94 9a 95 93 99 89 93 96 90 94 8d 8f 89 8d 95 99 97 95 96 9a 9d 95 92 93 95 97 9f 8e 97 9c 95 98 93 98 93 94 92 91 89 8b 88 8a 8c 85 89 82 7d 80 8a 89 84 81 77 7c 74 70 6d 6b 70 68 68 74 6a 6a 6a 64 6a 61 5d 57 5a 55 67 58 5b 54 5c 55 60 72 6e 57 4a 30 1c 12 04 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 12 1b 19 2f 48 42 5a 65 61 57 56 5a 64 60 64 65 61 67 6d 6f 70 7a 81 7f 87 7a 76 83 7d 7a 82 83 87 91 91 93 95 92 8f 92 9c 99 9b 97 91 97 9a 98 8c a3 98 8f 96 9b 97 9b 9f 92 96 99 9c 9c 9e a2 a3 ab a3 a2 a8 a8 aa aa ac ad ac a3 a9 a8 ab a2 a7 ad af a5 a9 a9 a5 9d a5 a4 9b 9e 9c 9d 9e 91 97 9a 94 9b 99 9d 9c 9b 9d a1 9b 92 9c 8d 8c 85 60 25 10 06 07 03 0b 06 07 04 00 06 05 03 00 06 05 03 00 06 05 07 01 09 0d 09 06 06 12 13 24 5d 8d 9f a0 9e a4 94 9a 98 9e 9a a1 96 8e 91 93 8a 93 90 94 91 95 8b 87 96 8e 92 90 8c 91 90 8a 8d 86 92 8f 8c 94 8d 93 92 8c 94 8e 97 92 87 8a 98 94 92 8e 84 8c 8e 7f 82 8a 88 88 82 84 80 84 84 86 84 74 7a 74 6c 6f 70 6c 6b 6b 6f 6c 6d 71 73 63 62 65 59 63 61 59 66 60 55 58 4e 5e 61 73 6c 5c 4b 32 1e 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 0c 11 2b 38 43 57 5d 61 5f 52 51 54 60 5f 68 5f 68 68 5e 70 73 76 7e 76 88 7e 81 7d 82 81 7f 85 86 80 8b 8b 92 8f 8f 93 8d 95 97 8c 95 9a 8f 8c 91 91 93 8e 93 93 96 92 91 8f 9c 91 9b 9b 9f a7 a5 ac a2 a3 a5 a1 a1 a8 a4 aa a2 a4 a8 98 a4 a5 a5 a7 a1 9b a3 a0 a4 9e a3 a1 9e 98 9a 8e 8f 95 96 a3 97 99 94 9b 99 96 92 99 99 95 97 92 96 89 5c 24 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 09 03 00 06 05 0a 0b 0c 0a 12 20 56 93 a4 a5 a1 9d 95 9b 9e 94 96 9d 93 96 92 91 97 8f 89 8f 93 90 8c 8f 8e 91 8f 91 90 90 8a 8e 8a 89 92 8c 8b 91 8d 89 8a 8b 99 89 95 93 8c 8b 8e 8e 8c 8d 84 86 85 84 86 88 7c 7b 81 87 81 81 82 79 74 72 6d 6a 62 68 66 64 6a 5c 68 72 6f 6c 68 61 68 57 5d 63 5b 5f 5d 5d 4e 59 51 52 68 6d 68 53 3e 34 1c 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 06 0e 21 21 31 41 4d 5f 63 5a 59 60 5a 5d 57 6a 66 72 65 69 6e 64 72 73 77 80 83 84 85 83 7b 7b 85 7f 86 8e 8a 8a 93 8b 96 90
 93 95 8d 8e 95 98 90 98 8f 8a 92 93 93 90 91 91 8b 92 99 8d 99 a5 a4 a4 9f a1 a2 a4 a5 a5 a2 a4 9f a3 a0 9c 9b 9c 9c 9e 9f a0 98 9e a1 9b 90 9a 9d 95 92 94 89 91 92 8d 92 8a 96 96 96 95 97 95 9a 95 96 a8 93 8e 88 5c 29 0d 07 06 03 04 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 0a 0d 05 05 05 17 12 10 1c 4a 88 9d a3 a5 9c 9c a0 9c 9b 95 99 8a 8f 8b 96 8c 90 8f 8d 8d 91 8b 8b 88 8b 8d 90 8d 8b 8d 88 92 88 8f 87 85 8a 8a 88 8d 8a 95 8d 87 96 94 8a 87 88 8c 82 91 8e 7f 82 82 8b 80 85 83 7a 7b 83 80 74 74 74 70 67 64 5f 66 6a 63 6f 68 72 6e 66 6a 5c 63 5f 61 58 5b 5f 67 58 5c 56 5e 5b 62 74 69 4d 3c 2b 19 15 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 06 09 12 19 21 31 49 58 5f 5f 59 50 54 64 5d 62 61 5f 67 6c 67 6b 5e 64 73 6f 7a 7b 7b 85 83 85 85 7e 7d 8b 81 8b 88 84 87 91 92 8f 93 90 92 94 87 89 8d 96 90 8d 90 8f 89 8e 8f 8b 93 90 9e 9a 9e a3 9c a1 9a a0 9d 95 a0 9b 9d 9f 96 98 9e 9a 9f 99 9c 9e 95 90 9a 90 99 96 8f 8c 87 88 93 87 8d 90 8c 8b 8f 91 91 92 95 91 9c 95 93 97 9b 8c 8b 83 68 31 09 07 05 03 03 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 09 06 11 08 0e 10 1a 55 8b 9f a3 a2 9e 98 a1 96 97 95 9c 8f 92 8c 8e 94 8d 8f 8b 8a 90 85 8d 8d 89 83 8c 87 83 8b 84 8b 85 83 85 89 89 8f 8a 8b 86 90 8b 8d 8e 88 88 8a 8b 84 86 86 86 85 85 85 84 80 7d 84 81 7d 76 6d 74 6b 6f 66 67 61 6d 60 6a 66 64 6b 6e 6b 65 63 5b 5c 5d 53 5a 5b 5e 67 56 56 54 53 61 6c 6e 64 50 39 29 17 12 0a 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 09 0b 1d 2a 41 49 53 60 61 5d 59 55 55 61 59 62 66 5d 70 6a 61 67 63 6f 74 76 7a 77 83 82 80 81 8c 90 7f 89 85 85 7b 83 94 91 8f 94 94 8b 8d 8e 8d 84 8f 8c 88 88 8a 8d 8c 88 8d 8c 97 97 9c a1 93 9c 9c 9c 99 99 8e 88 91 92 98 95 90 9b 93 90 9c 95 93 94 8d 8d 95 86 8f 92 8f 8b 8a 88 87 89 86 89 85 8c 8e 91 96 91 90 8c 92 93 95 8e 89 8b 81 5e 29 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 09 13 0e 13 38 84 9e a2 a5 9c 95 95 97 9a 97 90 91 8f 84 89 86 86 8a 85 87 86 85 89 84 8b 7f 84 81 7f 7e 88 7b 7f 83 7e 7c 7b 81 7f 80 8b 83 89 87 8e 84 89 8b 7f 7f 82 7d 84 7c 7f 82 7f 7d 7a 80 70 6e 73 6c 70 71 65 67 69 63 68 5e 65 63 6d 69 69 62 5f 5d 59 59 5f 5b 53 58 5f 5f 63 5f 5a 56 63 69 6c 5f 47 32 25 20 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 09 0f 20 27 37 48 55 62 62 60 5c 55 58 58 4e 5b 5e 64 6a 65 68 69 69 6c 6a 71 76 76 7e 79 7a 82 88 8c 87 89 7e 88 87 88 95 86
 8a 8f 8a 87 96 85 90 8d 8d 9b 85 88 95 90 90 88 8e 93 96 9c 99 94 99 8f 94 93 94 9b 90 94 8f 8b 95 94 96 96 94 94 94 8c 9c 96 93 93 94 8e 85 85 8a 8f 88 87 85 7e 7f 88 8a 87 97 8a 8e 8e 8b 91 9e 95 92 8c 95 8e 8c 62 32 05 06 05 03 08 06 05 03 00 06 05 03 00 06 05 04 00 06 06 03 04 06 0c 10 03 0c 0e 0f 14 37 7d a7 a0 a5 9e 99 9b a1 8c 95 94 95 89 8a 80 83 8a 87 8f 86 86 8b 7e 7e 84 84 7b 83 7f 7e 7e 7b 80 85 80 81 7e 85 84 7e 87 83 84 8c 88 89 81 84 8b 85 7e 81 80 7e 7f 83 77 84 79 74 70 68 6c 68 6d 68 66 61 61 5d 5e 65 5f 68 66 6b 76 66 63 5a 4e 5b 54 5d 59 5a 60 61 63 5c 52 5e 65 6c 63 52 3d 2f 22 19 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 02 0c 1d 23 28 3d 48 59 60 66 5a 59 56 58 55 5c 60 61 5a 65 61 70 71 66 6e 6e 6e 75 6f 6a 74 7a 76 85 87 91 8a 88 8b 86 82 8b 86 8a 8f 8b 8c 88 8e 85 89 8f 8c 90 8d 8e 8f 90 8b 95 9b 9f 95 94 92 87 8d 8b 8a 8e 8e 8e 89 8c 8d 92 94 94 94 8d 91 94 94 97 8d 98 91 89 8e 89 85 89 79 87 7e 90 86 86 84 8c 89 89 89 8f 92 92 95 97 9c 94 93 8d 8f 85 58 27 0a 06 05 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 0b 0b 14 12 3a 84 9e a9 ac 9f 94 9c 9b 90 90 92 83 90 81 85 88 80 88 8b 7f 86 7d 86 7f 81 7e 7e 85 82 7e 81 80 82 7c 7a 82 7c 87 81 7d 83 87 81 85 8a 7d 7a 85 80 7d 80 7b 7f 82 7e 7b 86 7f 79 79 6f 6d 63 68 68 63 69 62 5c 65 6d 5e 68 66 6f 62 64 5a 5e 5f 56 55 57 61 60 55 58 5b 5b 5d 54 5c 60 66 5e 43 35 2f 33 19 15 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 10 23 36 3c 4c 62 5e 5e 52 52 57 52 4d 5c 5d 61 65 64 63 64 70 67 60 6f 6b 6b 75 70 6f 71 70 72 76 7b 81 86 8d 89 7e 82 89 87 83 85 89 87 8d 85 8f 88 8b 8e 8c 8b 8e 92 91 98 93 8d 8f 8a 90 86 7e 86 82 83 84 82 8a 8b 8f 8d 86 8b 8c 91 8c 8a 8b 96 86 8c 8c 84 89 85 86 8a 81 7c 82 7e 7d 83 82 83 82 89 85 8a 87 87 89 8b 92 94 90 8e 90 85 63 32 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 0a 12 0d 38 74 a5 a0 9f 98 8e 99 92 8f 90 8b 88 7b 7f 7b 7e 84 7d 7a 79 75 7b 7f 7a 7f 78 76 7a 7c 79 75 7c 7d 77 70 7c 7f 7a 7c 82 79 80 7c 79 86 7d 85 81 80 7d 79 7c 80 74 87 79 75 77 6f 6f 67 5d 62 5f 65 5f 61 64 66 60 65 62 60 67 66 65 5c 57 5a 52 4d 50 54 57 5c 52 56 55 56 50 55 5c 60 5c 4e 3a 2b 25 29 14 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 09 18 1e 2a 3d 4f 5d 5e 59 55 56 51 60 57 5b 5f 5b 5c 6a 60 65 64 64 63 6c 67 7a 73 6e 6f 70 71 6f 75 6f 76 74 7d 7b 86 86 80
 81 86 85 86 8d 80 8b 82 87 90 87 89 91 8a 89 94 92 8e 92 85 91 89 83 7f 85 84 81 88 81 8a 8e 90 8c 8b 8a 8e 90 8b 8b 8e 8e 8d 87 89 88 81 7f 7e 7f 87 82 7b 79 83 7a 7e 7e 80 8c 85 83 8b 84 82 85 8d 8a 89 99 89 8a 64 28 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 03 0e 0b 0b 0e 13 2c 7c 9d 9c 9d 9f 91 9f 8f 8e 8a 83 81 83 7a 73 79 73 7c 7e 7a 7d 7a 77 75 79 7d 75 80 7f 75 7c 7f 72 7c 7a 7e 74 7a 74 79 77 7d 79 7e 82 7e 79 7a 7d 79 7c 74 7c 7f 7d 76 79 72 75 68 5f 5b 60 5d 57 5f 60 5e 60 5b 68 64 66 66 63 5b 5b 56 55 51 54 55 50 5b 59 56 55 53 4c 52 4e 56 59 51 45 32 2c 29 20 1a 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 06 0e 24 24 31 44 59 56 65 5d 59 58 5b 55 56 53 5b 5b 5e 68 60 64 69 6b 63 65 70 70 6e 6b 70 6a 6f 7e 72 6c 78 78 7e 7a 7d 82 82 79 7c 82 7d 85 84 81 84 84 89 8c 86 8e 89 92 91 94 89 88 88 7c 86 84 7f 83 82 7f 85 85 7f 82 87 85 7f 8c 8e 8a 86 8c 8a 8e 8f 86 89 86 8d 7d 80 84 80 86 7e 7e 80 7d 81 8a 7c 85 85 87 86 85 86 94 8d 85 90 8c 89 81 69 24 0a 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 03 00 06 05 03 0e 06 14 0f 10 27 71 a4 a4 a3 95 91 94 8d 84 89 8d 89 84 7b 75 77 7e 76 76 73 73 77 7b 81 75 79 7b 79 7e 6f 7b 78 7b 7d 7a 7f 7a 77 75 7a 80 7e 79 82 83 7a 7e 7d 81 78 78 85 79 7b 71 75 6e 71 6f 63 62 62 60 67 5e 5a 61 63 60 62 66 64 66 66 5e 5c 59 56 58 54 55 5b 58 5b 5d 56 55 51 4c 4d 4f 54 58 41 3b 35 25 23 1d 13 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 07 01 18 12 22 38 40 54 61 66 67 55 58 56 52 5b 53 61 5b 63 66 61 64 67 65 60 6a 68 6b 70 70 6b 6c 6e 71 75 71 74 73 75 6f 73 7c 75 71 82 77 73 7b 81 77 81 87 87 7e 7c 86 89 85 87 8c 81 7e 86 86 83 84 85 83 7e 7e 83 83 83 85 81 84 89 85 8b 8b 87 87 8b 88 81 7d 83 86 7b 85 81 86 7e 7b 6f 79 80 78 7c 7f 79 7f 80 78 83 8c 8e 7f 87 88 84 95 88 82 64 2a 0c 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 0c 09 16 0b 0a 25 71 9b a1 a1 9e 95 94 8c 87 85 84 7b 79 77 7c 7a 76 7f 7a 72 73 6f 74 7a 76 7a 7b 77 75 7b 78 7b 78 73 7a 73 77 77 72 7a 74 74 6f 74 80 7b 7e 7e 70 75 78 78 7b 6a 6c 6a 6a 5e 6d 59 5d 56 59 62 5e 5b 5d 62 63 62 65 5b 64 59 5f 56 56 57 55 5a 57 56 52 56 58 52 50 49 4c 4b 4f 4c 4e 37 2f 2d 25 24 19 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0f 1c 2f 39 45 57 54 61 61 5b 51 56 59 58 59 5a 59 60 63 61 61 5b 60 65 6a 65 68 67 6b 6d 75 70 75 74 70 70 73 6e 6f 6f 6a 74
 6e 6c 74 71 6f 72 71 76 78 78 7b 75 80 85 84 89 88 79 80 88 7f 87 85 79 89 77 84 7a 80 80 7e 7d 87 85 84 87 7c 81 8b 82 7f 89 84 8d 7e 85 7e 72 80 7c 7c 80 80 80 7f 78 75 79 78 7b 83 7a 85 85 86 87 87 87 8c 89 87 63 26 05 06 05 03 00 06 05 04 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 07 00 06 05 0c 0c 23 66 9e 9d 96 94 8d 92 81 7c 7a 79 81 77 78 6f 7b 7b 73 6d 76 7d 73 78 69 75 6f 74 73 71 7a 6b 70 72 73 78 75 7a 74 72 6f 7a 71 74 77 77 78 70 78 78 77 7d 6b 75 6c 6e 66 68 62 5b 60 5d 58 5d 60 5b 61 5d 59 64 5c 69 62 5d 5c 56 5a 4f 5d 47 50 5b 52 4c 56 4e 42 50 53 45 4a 49 47 43 33 3c 30 25 1e 1a 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0f 16 31 33 52 5e 60 5f 5b 5a 4e 5a 50 56 59 53 5f 5c 5a 5f 61 64 5b 5f 66 60 63 6a 6b 70 6f 76 77 72 6f 6f 71 6c 68 6f 6e 6b 6d 70 6f 6b 73 74 7a 71 72 71 76 77 76 7c 74 78 7c 89 85 84 7c 7f 7e 8d 7e 81 87 7e 7e 86 81 84 80 85 8a 85 86 88 85 83 85 81 8a 84 85 85 79 79 7f 76 78 79 7d 80 75 77 79 7c 7c 7b 7e 7a 7d 83 7e 82 85 83 84 85 88 5e 2a 09 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0a 0d 14 17 5c 92 98 99 8e 87 8c 84 80 7b 76 75 79 6f 75 74 74 76 6f 71 6e 6d 6f 6d 77 6e 6e 71 6a 70 72 72 6a 6c 70 69 72 71 73 72 75 77 72 76 75 72 78 7a 70 77 6b 76 6b 66 69 61 60 58 5f 61 5f 5f 57 5f 5c 61 66 64 65 57 63 5d 5b 51 55 52 52 51 51 54 58 56 56 4f 53 51 52 57 4d 4d 45 4b 40 38 30 22 25 27 1b 16 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 19 22 2e 39 48 58 5f 69 5d 55 49 57 54 5e 4f 59 58 5d 62 62 61 60 5d 5f 65 64 67 65 6b 71 73 6e 73 6f 6e 75 6b 6e 6c 62 67 68 66 65 6c 66 66 70 65 6d 71 76 72 6e 6f 71 77 76 79 75 7b 7c 76 7c 7d 81 7b 71 7e 7c 7c 76 80 84 87 87 7f 85 85 8e 7a 88 84 80 7e 82 7f 81 80 80 80 7a 7e 75 76 75 76 7a 75 71 7b 76 77 83 7c 7b 7d 82 86 84 83 87 7a 60 21 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 00 06 05 03 06 09 05 03 03 1f 5c 8d 8c 93 8a 80 80 7d 7a 77 75 77 74 74 6e 72 75 72 6f 70 73 70 70 67 72 65 72 70 61 6f 68 6e 70 6f 6a 69 6e 6b 6c 6d 64 72 70 78 74 74 73 72 71 74 68 67 59 5d 62 5e 5e 59 5d 5c 57 54 54 58 5f 5b 5a 60 5d 5e 56 5f 55 58 54 54 5d 50 59 5b 52 52 53 53 4d 52 4f 50 49 49 46 44 42 3b 31 29 25 22 18 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0b 0e 1f 1d 2a 3b 49 56 59 68 5a 54 51 4f 58 51 55 5e 4d 54 5a 5a 59 63 64 62 59 64 60 5b 72 67 6f 69 6e 72 70 71 6c 6c 70 66 64 65
 61 6e 69 68 5e 68 66 62 6a 64 67 6c 6e 60 73 75 6f 76 77 7e 74 76 7b 76 77 80 76 75 7e 7d 7b 7f 82 7f 85 88 82 86 85 7f 83 7e 84 87 79 84 7c 81 76 71 7c 7e 72 79 7b 70 76 79 7d 7c 76 7b 7a 79 7f 7b 7f 82 7a 83 83 63 23 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 0f 05 09 1a 52 8a 8f 93 89 86 75 76 7a 75 7b 78 74 74 7d 71 75 6c 73 66 6e 61 70 66 6a 62 6d 70 68 72 6b 69 72 61 6a 6e 67 70 61 6f 6e 6e 70 78 72 71 6f 6f 6e 6b 68 5c 5f 5a 5f 5b 66 57 50 53 56 57 5b 52 54 5c 5e 62 5a 55 5a 56 50 5a 5c 51 54 4f 52 54 54 4f 56 4d 48 4f 4b 47 4b 47 46 38 41 2f 34 24 1f 1d 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 13 1b 22 2f 38 4c 60 60 6c 61 59 55 5b 4e 4f 55 4f 56 5b 5b 58 61 5a 68 5f 5c 5c 5f 68 68 69 6c 6f 65 77 6e 65 70 6a 65 63 68 6b 61 6d 65 61 66 68 6d 68 62 63 65 65 66 72 6a 6c 68 70 73 70 70 6d 72 6b 79 78 70 7c 78 78 7c 82 80 89 7f 7f 7c 83 82 86 8b 84 86 8b 78 7e 7e 72 7b 7b 7b 75 75 70 72 76 7d 71 7c 73 80 74 7d 7c 7f 82 82 84 84 7f 7a 5a 1c 05 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 07 0f 4f 81 8d 8c 86 83 7d 7c 72 78 74 75 79 6f 6f 69 6a 6e 69 66 72 65 71 6a 67 6b 6b 6a 6b 63 6b 66 67 5f 65 6a 64 63 6d 63 72 7a 6f 71 74 70 6f 6f 65 63 67 60 60 62 5f 58 57 59 5f 56 5b 52 53 57 5d 62 5f 63 5a 55 53 58 55 55 5f 4d 5e 54 54 5a 50 56 51 4b 54 4f 53 4e 52 4f 46 41 3a 34 2d 23 23 1b 13 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0c 1d 39 3e 51 60 60 6c 64 61 59 56 52 5b 56 58 5b 5b 5e 63 64 5a 61 60 5e 69 67 64 64 60 67 6d 6d 73 72 62 63 63 6a 65 6b 62 61 63 64 67 62 5f 64 69 64 6b 62 61 69 64 68 67 64 6f 6d 6d 6b 6a 75 65 6f 71 6f 75 73 70 7c 7f 7c 80 84 83 78 7f 83 82 81 7d 85 87 8c 82 81 81 7b 78 78 82 7b 7d 7a 80 77 71 80 73 72 7a 84 81 7c 79 80 78 78 7f 7b 5d 20 0a 06 05 03 02 07 09 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 04 00 06 05 03 0a 14 49 7a 8d 87 86 7b 7c 83 79 79 6f 75 6e 74 73 71 6e 61 66 65 66 69 62 65 66 69 6a 67 62 66 60 5f 5f 6e 64 6b 64 64 60 66 5f 6e 69 67 75 5d 6d 64 61 64 60 5e 5c 59 55 5d 5a 59 5c 5d 55 52 57 60 5b 5a 5b 5d 52 50 5c 53 4f 52 5c 56 52 50 54 59 4b 53 52 4c 51 4b 4e 4a 4b 4e 44 44 3b 2a 30 24 29 16 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 05 0f 0f 24 26 35 4b 5a 59 65 6a 64 53 4f 56 4d 4d 5a 53 54 51 5e 5b 57 60 5d 60 64 60 66 5b 5f 64 62 6d 6b 6c 6b 65 64 68 64 65 63
 66 60 5d 60 5e 61 63 65 5f 65 5c 69 62 60 63 67 60 60 67 66 67 65 6d 6f 75 6f 68 6f 71 75 77 77 79 74 6f 83 7f 77 78 7f 89 72 8a 7f 7a 82 7b 83 7b 76 7d 7a 75 7b 77 75 7e 76 79 76 75 76 70 77 7c 7d 77 7a 74 7b 71 5c 25 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0e 40 77 7d 81 80 7b 82 7e 7c 78 73 70 6c 67 71 69 6a 69 6f 61 67 69 67 5e 5c 64 65 63 62 62 68 6a 65 5f 5b 62 60 5d 62 60 65 63 5f 62 65 60 61 65 62 5c 5d 5e 59 53 5b 5a 55 59 51 53 5e 4d 4f 5a 5c 60 58 4d 54 4c 54 4e 55 50 59 4f 5c 45 51 4f 4d 50 55 4a 51 47 4d 4b 49 44 3d 42 41 29 24 1d 20 17 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 18 23 26 38 47 58 5d 6f 69 67 5d 59 4d 53 4c 5a 51 59 53 57 5c 5d 53 5e 62 64 65 5f 5a 59 61 63 67 6d 68 65 62 65 64 65 65 66 60 65 56 63 65 5b 68 64 66 5f 60 64 62 62 6a 65 5c 63 62 62 60 60 63 68 67 6b 73 6e 70 6d 69 72 76 77 7d 7c 77 76 77 75 7d 80 7f 80 7c 89 88 84 83 81 79 84 81 75 7d 7f 74 76 76 77 6e 78 78 7f 76 76 7d 7d 79 7c 76 5e 1f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 04 04 13 3d 79 84 86 84 82 80 7c 6f 69 6e 68 6f 6b 66 69 67 65 61 61 64 67 69 65 66 5c 63 5d 68 62 5f 5e 63 62 5f 5f 53 5b 65 5f 5f 64 62 65 64 59 5b 5c 60 62 5f 56 5b 5c 5a 5a 5b 58 54 56 58 5f 58 62 5e 5a 56 59 5c 56 4f 56 54 51 50 5e 54 49 4e 4e 54 53 4c 4f 4d 44 46 49 42 43 3f 43 36 34 2b 24 16 12 08 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 08 0c 17 23 1d 31 47 50 58 6a 66 6d 5d 59 56 52 54 53 52 4e 55 4d 55 54 51 5a 5a 5e 62 5f 60 5e 59 63 65 67 6c 68 63 62 63 5c 5f 5d 62 63 67 5c 59 5f 61 5b 5b 64 5e 60 65 69 62 5f 62 63 64 64 61 60 66 62 62 66 69 65 61 68 74 72 79 72 77 75 75 75 78 79 7b 79 7c 7a 7a 7f 78 7a 81 7e 7f 79 7a 7d 7d 7f 77 79 79 75 72 7e 7a 77 75 78 7e 78 76 76 71 58 1a 06 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0b 05 02 14 34 70 88 81 80 74 73 74 77 6f 6e 69 6c 62 63 6b 6a 62 69 64 65 62 62 62 63 5b 61 59 62 65 5f 58 61 64 5f 61 5b 59 56 5e 5c 62 5d 63 5b 66 5f 5b 5f 5b 5b 5b 52 5b 5e 5b 57 55 54 55 59 59 61 62 54 52 57 57 62 52 58 4f 50 4c 59 59 5c 55 49 4b 46 4c 4d 49 52 4b 4d 4c 48 4f 40 3c 3a 2e 24 1c 19 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 06 03 0b 0a 22 1e 33 47 4c 5c 60 72 66 6a 61 50 48 44 4c 52 54 58 53 5b 4f 57 50 5b 56 5b 61 5b 5f 5b 5f 68 68 60 60 67 6a 65 61 69 60
 5e 5d 5c 5b 5e 58 5f 63 61 5f 61 5c 5b 62 5d 64 66 60 5a 63 5c 5f 61 63 68 61 63 5b 61 67 6b 68 6b 6a 69 71 70 74 67 72 73 6f 72 76 71 76 6d 76 7b 7a 7c 7b 73 7d 77 78 71 6f 7b 76 7f 73 7b 7c 73 78 86 80 73 79 75 67 1e 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0e 3a 6f 79 83 7b 73 74 77 6f 6f 6d 6d 6a 6c 62 68 65 6a 6e 6a 67 68 5c 61 63 55 65 5e 63 60 5f 60 62 5d 5d 5d 5c 54 58 55 58 5c 5a 60 5a 5d 5c 5e 5d 59 5a 54 56 5b 56 51 59 58 56 61 5c 5b 5b 56 53 57 56 4e 52 4e 4d 47 4f 55 4f 4f 4b 48 4d 54 43 49 48 51 40 51 51 49 4d 49 44 40 32 24 1b 1a 15 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0f 13 1c 25 2d 3e 47 53 60 6c 75 6e 63 59 4a 4e 4c 4d 51 50 5a 50 54 53 5a 65 59 5e 5f 57 60 5c 5e 6a 64 63 61 5f 61 65 64 5f 63 65 62 65 62 65 5e 65 69 5c 65 5d 60 64 64 5b 61 64 5b 69 61 58 5c 5c 5e 64 6b 5c 67 62 64 6a 6b 70 75 72 71 65 6a 6c 6d 6c 6f 6f 72 6c 6e 72 75 7a 75 76 7a 76 77 72 6d 76 72 6a 79 77 72 76 75 77 72 84 8b 7b 76 7c 5c 20 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 2a 67 70 75 71 67 74 72 6b 70 72 6c 73 66 6d 72 68 72 62 61 5e 5e 62 5b 62 5c 5b 5a 5d 59 59 51 54 52 53 5f 5e 5e 61 5b 60 5b 60 65 55 57 59 56 54 5d 55 5a 55 5a 56 55 54 57 56 5d 54 53 57 57 53 5c 54 54 54 4b 4f 4f 53 5a 51 4d 4f 4d 48 4e 4a 50 4f 4c 45 4a 49 4d 56 4c 49 3f 3a 24 20 17 0c 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 09 15 12 22 26 3c 45 52 5d 5d 66 70 65 56 4e 4d 51 54 54 5b 58 57 4e 5e 54 62 54 59 5f 62 56 5a 60 5e 63 62 5e 5b 58 59 5e 5a 64 60 66 63 61 64 5f 64 5b 6a 61 57 5f 5f 62 5b 67 62 64 5e 64 5e 63 5f 5f 56 5b 66 64 67 60 65 6c 65 66 6e 6b 6f 71 67 69 74 6b 72 6c 6d 6c 72 75 6e 70 69 71 74 79 75 72 7a 78 81 76 73 7a 73 76 7a 75 7b 80 78 6e 77 5d 1f 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 00 0a 28 5c 70 6b 75 64 70 72 70 65 6b 6d 64 65 66 6d 6d 63 6a 67 64 5b 63 5b 5f 59 5d 59 5e 56 5a 61 55 56 5a 59 50 59 59 5a 5c 5d 5d 58 66 62 58 5d 5c 56 57 61 51 55 5a 5a 5e 5c 5f 59 53 51 56 5b 53 55 53 52 47 4c 4e 51 4b 4a 56 51 57 50 54 4d 4f 50 4d 49 4c 4b 4f 53 52 4e 44 33 35 30 20 19 0b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 14 17 1d 2b 2c 45 43 46 5c 65 6a 67 61 50 4d 50 51 53 52 4e 56 46 47 50 55 5b 5e 50 5b 59 5b 5b 5b 60 5f 5a 5a 64 52 54 59 61
 5b 66 5f 62 63 66 63 68 65 64 58 66 5e 54 64 60 61 60 61 62 63 56 62 5d 62 59 5a 5d 5c 60 69 65 65 64 63 6a 63 68 66 66 72 62 67 6b 70 70 6f 71 73 68 6d 70 6e 74 72 6e 73 66 70 70 6d 73 77 72 75 75 7b 7b 7b 71 7a 5f 23 03 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 1f 54 61 6c 6a 5d 62 66 65 6a 68 5b 67 68 62 65 5e 6c 6a 67 65 63 57 58 5a 51 5e 55 5b 5a 55 59 57 54 5c 52 53 53 59 52 58 51 5d 5b 56 57 55 5d 62 59 5a 54 57 4a 5a 55 53 53 51 52 5f 50 51 5a 4d 56 50 51 4c 50 4c 55 4e 4c 54 4d 4a 4f 47 47 49 50 48 4d 45 50 52 4f 50 4a 38 3e 2d 2b 1d 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0b 1a 18 24 2d 33 40 39 4c 5c 63 5f 55 50 55 4c 58 4f 51 4a 50 54 54 57 55 5e 63 5d 55 58 67 5e 5c 62 55 5c 59 5c 5e 5f 67 67 69 61 63 65 5a 60 5d 63 66 62 60 63 5e 62 54 61 63 58 60 5d 5d 63 56 61 5c 62 5e 62 5c 63 63 62 5f 64 61 67 60 61 66 68 64 6b 73 67 66 68 65 6b 70 6b 6e 6f 6d 69 6c 69 6f 74 73 70 6b 6f 6b 77 77 7a 7b 6d 74 75 74 65 21 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 1c 53 5e 5e 6b 5d 68 67 60 64 61 62 64 5d 61 64 64 6a 68 62 63 59 5f 4f 57 5b 5d 54 5f 53 59 55 51 4d 5a 53 56 58 5c 58 59 5b 52 57 52 50 50 57 54 5b 5b 59 55 5a 5c 58 5c 55 50 58 52 52 54 52 51 58 53 4e 45 4e 45 48 54 49 4e 4e 47 53 4c 46 46 47 4a 47 48 48 4d 53 4c 4a 34 34 32 23 18 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 0f 16 1b 1f 2a 34 39 35 3f 48 4f 61 55 50 52 56 51 56 51 57 53 5d 5e 5f 5d 58 57 62 61 54 5b 50 58 5d 5b 5a 5c 60 57 5e 63 69 6b 71 6e 66 62 5e 69 66 62 6d 68 62 5d 60 5d 59 5c 63 5f 65 5c 60 65 5f 68 59 5b 5f 67 5f 62 64 5f 69 5d 6b 67 65 62 6a 64 6e 67 6c 6d 65 6c 6f 65 71 72 65 68 6c 6b 6c 68 6b 72 73 6c 70 71 70 70 6f 72 76 74 77 72 5b 24 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 07 06 06 17 4f 59 5b 63 56 61 66 67 5a 64 66 64 61 63 6b 64 66 6e 67 64 64 5d 57 5b 57 50 60 5e 55 59 5b 5b 52 56 56 56 56 56 55 55 57 5a 5a 61 5b 52 61 58 5d 5b 58 54 4f 58 58 56 5b 54 53 56 4f 52 55 54 56 52 53 50 53 53 5a 59 4b 4e 41 52 50 4e 4f 53 43 4e 51 51 57 49 50 48 3d 37 2e 2a 22 10 12 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 1a 16 1c 2b 2a 2e 38 36 35 3f 42 50 4b 4a 54 4c 4b 55 55 4f 63 5f 65 62 60 61 5b 57 56 53 52 57 4f 51 50 56 63 57 5b 5c 69
 73 77 6a 65 67 5e 63 64 62 63 5b 65 64 5e 60 62 56 63 5a 63 57 5f 5e 5b 5c 55 5c 62 57 5b 60 64 5b 5e 58 5a 63 65 58 66 61 68 69 66 68 69 64 5b 6f 65 6a 71 6a 69 6a 6c 6c 6d 5d 60 63 63 6a 6e 71 69 68 64 68 6e 66 5c 27 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 1d 42 62 61 5d 5c 61 5d 55 60 5b 5d 60 5f 59 60 54 63 65 66 67 61 59 53 59 4f 5a 55 59 5c 57 55 54 54 4f 59 56 5f 5d 54 53 56 50 5a 59 54 55 59 5b 56 55 54 52 57 4f 59 58 57 53 55 56 52 4a 45 4d 59 55 57 4c 4e 48 4b 4f 4e 4e 4d 4c 47 47 50 40 47 4d 55 56 54 4a 4b 4a 45 32 31 25 1b 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 10 0a 18 1e 25 2b 2b 2e 33 3c 41 45 4b 43 4e 4d 4b 4f 4b 59 56 5b 64 63 68 61 5d 56 61 52 57 58 54 4c 58 4f 58 5c 64 70 67 64 6c 62 69 67 66 64 64 67 68 5f 5c 5d 5c 61 61 60 5c 60 5e 5e 55 59 55 5c 54 5b 5c 5c 5b 59 58 5f 64 5f 68 64 5f 5d 66 62 69 69 5a 62 64 60 69 63 5f 63 6c 69 6a 66 67 62 6c 6a 64 62 65 6d 63 63 66 6a 60 5d 58 60 51 20 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 46 5b 55 5a 54 51 58 5c 57 56 58 57 60 59 5e 5f 64 63 66 62 65 59 59 55 50 52 60 56 57 5a 57 5b 57 58 64 5f 5b 59 59 58 56 53 5b 52 52 54 5b 57 59 54 55 5d 5b 5d 59 56 53 51 58 4e 4f 51 56 46 4a 4d 53 4b 4a 51 4a 48 4b 4a 49 50 49 4f 47 45 50 46 55 54 52 4e 48 45 37 38 25 1f 0f 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0c 13 22 2b 2e 2f 32 31 36 3a 38 46 40 48 40 4e 47 54 4d 55 52 54 62 5f 5d 60 57 53 52 56 59 58 61 5a 55 58 51 62 6b 61 69 6b 66 63 5f 60 5d 65 5b 6a 61 62 67 5f 65 58 5b 60 65 60 5b 5c 58 60 5b 5b 64 5e 64 61 54 5f 60 5b 61 62 5c 61 65 62 65 5c 5e 62 64 5d 64 66 67 69 69 5e 66 6d 70 64 6c 6d 66 6b 6b 6b 65 69 59 5f 62 57 53 60 52 48 25 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 43 50 5b 54 4d 56 59 5c 5c 61 54 53 5a 62 62 63 68 68 60 65 5a 5d 54 5c 5a 58 50 59 57 55 61 54 57 5d 57 57 59 5d 5b 50 53 50 56 50 52 5c 54 60 5b 5d 56 56 51 59 58 5a 5e 52 51 50 4e 4e 54 4e 51 5a 56 58 49 4f 4b 49 50 59 4e 51 46 4b 42 4c 4c 56 5a 56 52 49 51 44 3b 2b 30 24 07 0b 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 1a 18 1e 23 26 33 30 33 39 3b 3e 42 46 3c 49 45 4d 4d 45 48 53 50 61 5f 62 5f 56 57 59 5a 5a 5a 51 52 51 56 5d 5e 62
 5f 65 60 5c 62 63 64 64 6a 5d 64 5d 64 67 5d 59 65 5d 5e 58 5f 5e 58 61 61 5a 55 55 5f 5c 59 63 64 62 5b 60 50 5e 64 5e 66 58 60 60 67 5a 5d 61 67 69 63 6c 64 64 68 5d 68 66 5f 5d 60 6d 63 61 60 64 5a 5b 4e 53 51 47 21 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 37 54 5b 59 4c 5d 5e 4c 60 58 64 5d 5a 5e 5b 61 5e 5a 5e 56 57 54 52 55 4d 55 50 5c 5a 5c 59 54 59 5e 5b 60 5a 5a 55 54 56 54 51 50 4e 4e 56 5c 56 58 51 50 58 58 58 54 56 51 51 59 50 55 55 59 51 56 53 48 45 49 4c 44 49 4f 49 49 42 48 44 46 4b 50 55 53 4c 53 47 43 34 2f 26 1b 07 02 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0e 14 21 1e 23 29 30 2a 36 34 3e 36 39 42 46 44 4e 4b 45 4c 4d 51 54 59 5f 5c 5b 52 5f 56 52 59 4f 55 59 5b 61 5f 51 59 60 5a 52 5c 5c 5b 59 5d 5f 64 58 5c 5c 56 61 5d 5d 5a 57 5c 5a 65 54 5c 58 5c 58 5c 5c 5c 64 60 5d 63 55 61 60 62 5d 62 5a 64 63 57 5b 5f 64 62 64 5b 54 60 5e 61 62 61 65 5f 61 56 62 63 64 5c 56 52 4d 4d 4f 48 44 1f 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 0f 38 4f 56 55 53 5b 52 58 51 5d 53 5b 58 5e 5f 5c 65 6a 62 64 5b 5f 54 54 4f 4e 54 55 52 5a 63 63 61 61 5e 59 51 5d 51 5a 50 4f 54 54 50 4f 56 58 53 4d 4b 4c 50 55 52 58 50 53 4d 54 51 58 4b 4a 53 53 4d 4f 48 4f 54 51 53 4b 4c 46 49 4c 4e 49 4d 50 4d 54 53 4b 4a 38 2e 22 1f 16 0d 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 16 17 24 20 23 30 32 33 31 39 40 39 35 3d 44 46 42 43 3f 45 4f 51 57 60 5a 54 4e 4c 58 55 58 55 4f 52 5b 5f 5b 5a 60 5f 5a 5d 5a 5f 58 64 5b 5f 5a 5c 5e 5e 59 57 62 5c 61 5b 5a 5f 59 61 5a 5d 5c 54 52 62 56 5f 5e 54 55 63 60 60 62 53 5d 62 63 64 5d 63 58 60 5e 57 60 66 5c 5d 65 5c 5e 59 66 63 5a 5f 58 57 55 5a 55 58 51 4b 4e 45 22 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 3b 4f 5f 5e 5b 57 56 59 53 5f 5b 5b 5c 56 5c 61 5f 63 5a 54 5c 54 50 55 4f 54 51 62 53 65 68 64 65 63 60 5d 50 55 52 58 52 54 52 4b 4b 53 56 54 4f 53 50 57 55 51 4e 4d 4e 4c 4f 56 4f 58 50 55 56 5a 50 4f 51 4c 4c 46 50 50 42 4d 47 4b 4a 4b 4f 49 4c 50 47 55 3b 39 32 22 1b 11 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 02 10 14 1c 2b 2a 26 27 30 35 3f 3c 39 42 3c 44 4d 40 43 47 43 47 52 5e 63 5c 4e 53 4f 57 5e 5c 55 5a 59 59 58 57 5c
 5d 60 60 5a 5a 5a 5c 5e 56 5c 5b 61 61 5c 5d 55 63 5d 56 5f 58 5b 53 58 57 5c 57 5f 56 56 57 58 5b 5a 55 5a 59 58 56 59 63 59 5e 67 62 56 60 63 60 61 61 66 5c 62 69 60 59 60 62 62 5d 5f 5a 5a 57 5f 59 49 51 4d 53 48 26 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 32 52 59 59 50 55 58 5c 5a 5d 56 58 59 56 61 60 62 63 62 5d 55 50 52 55 46 55 63 58 60 5b 5c 63 57 59 5f 54 5d 5b 59 57 57 53 56 54 4d 45 55 54 4e 51 4a 54 53 50 45 54 51 4f 5a 53 51 50 4d 53 59 5e 55 55 50 54 4b 4c 4c 4f 4a 45 52 46 42 44 4b 4f 4b 4f 46 45 3e 36 35 26 15 0e 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 09 12 12 1e 25 28 2f 38 37 34 32 3c 35 3e 3b 41 3b 47 40 47 52 50 58 63 5e 51 50 4b 55 56 52 44 4a 58 5b 58 56 63 61 61 59 55 55 5c 53 52 57 57 5a 52 5d 56 68 5e 58 56 65 59 5e 5c 59 60 62 60 56 5c 50 56 57 56 54 57 57 5a 5c 5f 5f 59 61 5d 64 5d 5b 63 65 5d 5c 65 67 5a 60 61 66 64 5b 5b 5c 5f 55 5b 56 56 55 4f 54 52 53 49 4d 44 26 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 27 59 51 54 55 58 61 5d 60 5f 5a 5c 61 57 62 61 56 61 60 59 57 53 51 54 5b 55 5d 59 5e 5b 5f 5e 5a 5d 5b 4e 52 52 50 52 4c 50 4a 4c 4f 4e 4b 4d 49 4b 50 51 51 48 45 50 4f 55 57 50 51 52 50 58 5e 5f 54 52 4f 53 4b 4b 45 4b 4b 4b 4b 45 40 45 49 42 43 47 41 45 3f 30 25 1b 0b 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 0b 19 22 24 1e 36 34 35 37 33 34 38 40 3e 3d 41 42 41 40 45 47 4c 55 60 5b 4c 4d 4f 50 54 50 57 5c 4d 5a 57 5c 6b 5f 58 54 53 59 57 54 5a 5b 53 5a 4a 61 5a 57 5d 5a 56 60 58 52 61 56 5a 5b 5f 5b 56 59 55 56 57 58 5a 5a 55 52 5a 61 62 60 5d 5d 5e 60 62 58 62 5a 62 5e 5f 57 5d 56 53 5f 5b 57 59 5b 59 53 52 55 53 48 49 4d 49 42 27 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 35 51 61 5d 5a 61 5a 5c 63 61 60 5d 61 5c 5e 59 62 5a 55 57 5a 55 56 56 59 60 5e 65 69 5e 5c 52 52 4e 4d 4b 52 4f 4d 51 56 54 55 4b 52 56 4d 4a 49 49 48 51 4f 46 52 4e 4e 4e 50 56 4c 50 53 59 5f 5f 66 57 52 4d 47 43 49 5b 46 49 47 50 49 44 47 45 47 41 3d 36 38 2a 2d 13 06 09 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 10 1c 1d 25 25 29 38 34 3c 33 38 36 3b 45 42 42 43 36 3f 42 50 46 55 57 56 4e 47 51 4c 4b 4d 54 55 59 55 4f 5a
 5f 55 58 52 51 53 49 4c 55 52 59 5d 54 50 56 50 56 58 54 62 59 56 5e 51 5e 59 54 59 53 5c 61 59 5c 58 5e 5c 57 5c 5b 5e 5e 5c 59 5c 5f 57 61 5e 60 60 61 5b 5e 5f 56 5c 56 60 5d 5d 51 56 51 4e 57 58 51 45 4b 4b 49 46 1e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 2b 5f 57 61 4e 55 5b 5b 5c 5e 63 5e 5a 5e 5d 59 59 5d 5e 54 56 54 55 5c 59 57 55 5a 5f 58 59 52 49 4d 54 50 53 4a 4e 4c 52 4a 4f 4b 40 4e 47 50 45 47 4c 4a 53 4b 53 54 50 4f 51 4d 51 54 53 57 5d 62 5b 61 52 4f 43 44 4e 50 55 4e 4b 4d 42 44 3f 3c 3e 4a 3d 35 36 2a 1e 10 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0e 11 1b 21 27 2a 2a 31 35 33 35 3c 3d 42 45 46 47 43 40 41 42 3f 4b 4a 4c 4b 43 41 4f 44 48 50 51 50 50 56 57 54 5d 59 53 4c 4b 48 50 4a 4e 45 55 54 4c 4d 54 4f 57 52 58 4e 54 5d 64 60 59 5c 54 50 4d 59 56 57 5c 53 52 58 52 50 54 57 56 59 5a 59 64 65 60 60 5b 5c 5e 5c 56 5c 54 54 55 5a 5d 58 5b 4f 53 50 53 55 4a 4d 44 51 47 24 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 27 4e 5e 65 5f 5a 64 56 60 60 5e 5a 56 5b 56 54 5d 57 58 52 52 5b 53 59 5a 55 56 60 52 5c 4f 46 4c 47 4b 48 48 4e 4f 4e 4d 41 40 4d 43 45 40 48 45 41 4f 52 47 54 4f 4f 50 50 4e 4a 50 51 55 54 55 4d 50 5c 4e 4f 4c 4a 49 4b 40 4c 47 4e 4a 45 49 43 45 48 3c 3b 33 20 17 0c 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 12 21 1d 1e 31 2b 2c 35 32 34 3c 45 47 44 38 41 3e 3e 43 42 45 41 4f 44 4a 4d 49 44 44 50 50 52 58 4a 58 58 57 58 5c 58 52 50 4a 4a 50 4b 53 4a 4b 4e 56 4e 4b 51 55 56 51 54 59 59 55 54 56 51 56 56 5a 5a 5c 5c 51 54 51 57 5c 59 60 53 58 58 58 5d 5e 5e 55 5a 5e 5f 52 62 57 55 5b 52 53 4e 5c 52 59 53 4e 4d 4f 54 49 52 4a 48 2f 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 28 4c 5b 62 53 5f 61 5e 52 55 58 5c 59 56 58 4e 54 5c 56 55 4d 5f 56 57 59 5b 55 58 57 53 50 45 47 4b 50 4c 3d 54 4d 4b 4e 47 40 50 45 42 45 46 40 43 4d 47 4a 52 4b 52 55 51 4f 4c 53 4b 4d 4b 49 51 4e 4a 58 59 4e 4a 4a 50 4d 4b 49 46 45 44 4a 41 4b 3b 3f 33 32 22 16 0c 0b 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 07 10 18 26 24 37 32 2e 39 3a 3b 3e 46 44 41 40 3a 3e 3a 39 4a 46 46 45 3f 41 49 45 50 4c 4f 4f 4b 54 58 59
 5d 5a 5c 60 60 53 4b 4f 4d 51 4a 49 4f 53 50 5c 53 53 50 54 58 52 50 53 58 56 4f 51 53 56 58 51 55 51 4d 5d 4f 59 4f 54 5a 57 59 5a 5a 5c 5d 5a 63 5e 5b 59 5b 5a 50 53 56 50 5a 59 4a 5a 55 54 59 53 55 4d 49 4a 50 4d 27 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 24 56 5d 63 54 5b 5c 59 5e 5a 53 59 5e 54 52 54 52 54 51 52 57 5f 4b 63 53 60 58 5d 55 54 51 4e 4a 40 48 4c 47 49 45 46 46 49 45 45 47 48 4e 44 4d 48 43 4e 4a 50 43 4a 5b 4e 4d 44 4f 4e 48 43 4c 4c 53 57 4c 50 52 44 4d 56 41 4a 4d 46 4a 3c 45 46 4b 3e 3a 30 30 25 12 07 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 10 17 20 28 2a 28 2c 35 35 37 41 4a 45 3d 36 3e 42 3b 36 3a 41 44 44 43 42 49 4c 46 47 4d 42 48 47 49 52 52 5c 56 5a 52 4b 48 50 52 41 50 49 48 51 4d 52 53 4f 58 55 48 59 54 54 4c 4f 55 50 4d 4c 50 4d 57 53 56 55 4f 56 54 4f 5a 54 56 5e 62 5a 5b 5c 5c 55 60 54 51 56 58 54 56 4f 53 4f 59 4f 56 59 58 4c 44 4f 51 51 4f 45 22 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 22 4a 5b 64 53 58 57 5c 52 5b 5a 5c 52 50 52 4d 53 59 57 5f 50 58 51 5b 5c 59 59 51 4f 4c 4b 49 3f 49 42 44 49 46 45 48 54 44 46 4b 41 45 44 40 3f 44 4e 4f 4b 48 46 46 4a 49 42 48 44 46 45 45 4c 4b 53 52 4a 4b 51 4f 4c 41 4a 44 3c 4a 49 41 47 44 45 3b 35 31 28 13 1a 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 1c 24 2a 26 34 31 30 2f 3d 44 4f 4d 3c 3f 37 43 3b 39 3e 49 41 44 43 45 49 47 45 46 49 4d 48 4c 4c 53 4d 56 52 4b 50 52 56 4e 44 4f 3c 49 49 4a 57 52 52 4f 52 4f 48 4f 54 4f 4f 51 53 50 4d 50 56 5b 5f 5b 52 52 4f 4f 59 55 53 58 58 5b 5d 5a 50 5e 5e 51 59 57 56 4e 4d 51 53 56 54 5d 55 5e 4e 55 4a 51 4c 4c 4c 51 59 4d 2c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1d 45 56 50 4c 57 59 54 52 4c 56 54 4f 55 49 4d 4d 53 57 5a 57 54 53 63 53 58 52 5a 4d 4b 47 54 4b 48 4d 3e 48 48 48 4e 4b 4a 44 49 49 46 47 48 3f 46 41 49 4a 4d 4d 47 48 41 44 49 43 47 44 46 4e 44 4e 47 4c 4a 55 47 48 46 4a 40 4c 4c 47 45 3b 43 3a 39 35 2c 22 17 0d 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 15 19 27 2b 35 2f 34 35 39 42 4d 49 3b 3f 45 3e 3e 45 3c 3b 43 41 42 41 46 42 46 4b 4b 46 4c 4b 4f 50
 53 4b 4e 4b 59 50 45 4e 45 4a 4e 4c 49 51 49 44 4f 4e 4e 4e 52 4f 54 48 53 54 5a 50 50 54 51 5c 51 53 51 52 4e 54 54 4e 51 51 58 59 5a 58 5b 58 57 58 5b 52 5a 50 54 54 51 55 57 50 50 55 56 56 4c 50 45 51 4a 5e 52 4d 32 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 1c 4c 4c 4b 49 4c 4d 4b 53 51 59 55 54 53 56 54 57 53 51 59 59 53 55 55 56 5a 56 51 56 51 4c 4e 4e 44 3f 49 46 4d 4a 43 45 44 44 45 4a 4c 4b 46 40 45 4b 4c 4d 52 45 46 51 4f 4b 3e 40 47 47 46 4c 48 4f 4a 4c 5e 49 44 44 4a 48 4d 3e 4c 43 3d 4a 3e 43 34 33 21 21 13 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0f 16 22 28 31 2f 2b 3b 3a 3a 4b 48 42 3e 39 44 3a 3d 40 4a 43 40 3f 3e 43 44 42 47 44 49 42 49 49 53 49 49 4d 4a 51 52 4a 54 49 4d 50 4b 47 3d 4e 49 48 47 49 50 4f 44 4d 4d 4b 51 4b 4f 47 53 5f 5a 5b 59 4f 4e 5f 56 57 4e 52 59 5d 5c 56 50 57 57 5a 56 55 57 53 4d 54 53 52 51 54 4c 50 52 56 55 52 46 4b 48 4a 49 56 4f 24 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 42 46 47 46 4c 4f 48 54 4f 50 57 52 50 55 4d 4a 56 52 54 49 5e 4d 58 4d 50 4b 4b 47 4e 4f 48 48 49 49 44 3f 4b 3d 3f 4f 41 40 49 46 47 47 48 4f 42 47 44 49 4c 4d 45 45 4a 47 47 42 42 44 4b 4b 50 4c 4a 4a 40 4b 43 44 4c 47 44 46 45 4b 41 40 43 3e 3a 2d 25 22 0c 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0e 1e 21 34 31 2f 3c 31 44 42 45 3e 39 3e 3a 42 4a 3a 42 3c 3d 43 39 42 40 3d 45 47 47 4f 53 54 4a 4f 4a 46 53 4d 4c 4c 45 4f 45 45 49 43 49 49 4b 50 4f 4f 41 50 43 47 4e 4b 4b 4c 49 52 4f 57 55 4d 5a 59 52 50 56 4b 4c 4f 51 54 5a 4a 50 4f 51 4e 4f 4f 4c 4f 4d 57 52 4a 53 51 50 54 4e 4e 4e 4b 54 45 46 50 52 47 2d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 36 3e 45 4a 4a 46 4a 47 56 4f 53 4d 51 51 4f 51 53 55 4f 52 52 4e 4e 50 4e 44 4a 44 54 48 47 45 42 43 42 45 3b 3c 44 45 49 3f 43 45 4c 45 3f 4e 3f 49 4d 3f 49 42 48 45 47 42 42 44 4d 47 46 48 50 49 4e 45 43 42 46 47 4a 47 49 3a 41 3b 3e 43 3a 3f 2f 29 22 15 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 15 1f 23 31 32 30 37 3b 3f 3d 47 45 3e 40 45 43 38 43 42 3a 41 43 43 4b 40 44 47 47 41 4c 4e 4d
 45 4b 4c 54 56 57 51 4d 4a 4b 45 49 4c 43 46 47 4f 50 4a 4d 49 4a 53 44 54 4a 4e 49 44 4d 4d 57 56 4d 52 55 52 59 50 52 56 51 4e 57 55 4c 4c 4e 52 4f 52 4d 50 4d 5b 53 52 53 57 56 54 4e 50 46 54 51 50 54 4d 50 4d 4b 2e 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 2f 42 46 48 48 47 3e 4e 49 57 55 4d 54 55 52 57 56 4b 55 4f 4c 52 4d 50 4b 47 48 43 45 46 46 42 48 47 47 41 37 48 3e 45 4c 45 45 45 4f 4a 4c 46 49 48 41 47 4b 40 4c 44 43 49 47 4c 49 4b 4f 4b 4e 49 49 47 4b 3e 49 4b 43 4c 45 3e 47 48 49 46 3a 40 34 24 24 10 0c 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 17 1e 27 28 2c 30 36 38 3f 43 41 3d 3b 43 3c 35 3f 3e 41 43 40 3c 3d 40 3f 44 42 49 43 4b 4d 4c 4a 4d 3f 4b 4f 55 51 4f 49 43 40 40 42 4e 47 4c 48 46 4a 48 48 48 47 46 4a 4b 53 4b 40 3f 4d 50 4a 4e 52 4f 56 52 5b 53 56 54 4f 52 4b 51 53 50 52 4d 4c 4f 4f 54 52 52 50 58 59 55 4f 59 50 54 4f 51 49 4c 46 49 45 46 2d 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 2f 46 4d 47 4b 4a 4a 4c 4b 4a 4b 4a 54 49 4c 55 55 4f 4a 48 50 48 4f 4d 44 47 41 3f 44 46 41 41 40 41 46 46 46 40 42 47 47 41 43 47 47 49 4b 43 4a 3e 41 42 48 42 4d 41 46 49 44 47 49 50 52 4f 4b 49 4b 48 44 49 4e 47 47 49 4d 47 44 46 41 48 3e 32 2d 1e 15 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0f 26 25 2c 2a 2b 35 3e 41 41 45 38 39 44 37 38 43 40 42 3c 3d 37 36 46 45 3b 48 41 45 44 49 48 44 41 46 4c 50 47 52 46 59 42 42 4b 53 47 44 41 47 44 4a 4b 42 47 45 4a 4b 51 38 46 45 4e 50 47 49 4d 5b 52 50 52 55 5c 54 4e 54 4f 56 48 54 54 4b 4d 53 48 54 50 55 58 54 57 58 57 51 55 54 52 51 4c 4a 43 43 4d 43 24 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 2f 45 47 37 4b 41 40 4a 4c 49 4d 41 45 4b 4b 51 4c 51 51 4a 43 3e 4a 42 4a 4d 45 49 46 4c 43 50 40 45 49 44 46 43 44 43 45 4a 48 39 3b 42 3c 46 3c 4a 46 44 49 4d 4a 42 41 3e 46 44 49 4f 49 4e 4b 49 49 41 42 44 41 49 4b 48 51 3f 47 43 41 42 35 37 31 16 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1a 18 21 26 30 2e 36 3c 40 41 3f 3b 44 45 3f 3d 41 3c 44 45 3d 41 41 41 41 41 46 37 39 3c 45
 42 47 44 47 48 4e 50 5c 4d 47 50 4b 43 47 4a 4b 4a 4c 41 51 47 4e 46 3e 49 47 45 49 46 49 4d 50 4e 4a 45 52 4b 54 5a 53 56 4f 52 53 4b 52 4d 53 51 51 54 57 4d 5c 55 54 55 50 5e 56 5a 50 57 53 51 4f 55 48 52 49 41 44 2e 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 3c 3d 43 40 46 46 41 44 44 45 4e 44 44 45 48 4a 47 41 4b 46 4e 3f 44 46 42 42 49 46 45 48 46 46 43 42 45 42 41 42 48 42 43 47 48 44 44 4a 43 40 38 49 43 3f 40 41 4a 4c 48 4d 4d 49 4b 4e 48 49 4f 4c 4c 44 45 44 48 41 46 4a 48 46 49 3d 3f 3f 31 2d 28 19 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 0d 20 28 29 26 34 45 43 3e 41 3b 39 39 43 45 3b 45 46 3c 3d 3b 44 40 49 3e 41 3e 3b 44 3c 40 47 45 45 46 40 46 58 4e 50 49 4d 46 4a 4d 44 4d 46 42 45 41 49 47 47 49 41 3f 4c 4c 47 4e 47 4d 4e 4b 52 54 4d 4e 52 5a 53 55 55 49 51 4d 4d 58 52 53 54 47 57 58 5c 4d 58 5e 5a 5c 56 54 53 4a 52 4f 48 45 48 4a 45 2c 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 2a 3c 45 41 47 44 3e 3f 48 3d 49 46 47 42 45 4d 48 46 48 48 43 3d 44 45 48 46 43 43 46 47 42 40 45 45 47 44 41 41 40 41 46 43 46 41 3f 4a 46 46 43 48 41 41 45 43 43 4e 46 48 49 4b 4e 44 4c 4c 45 49 43 48 46 48 47 46 51 4b 4f 3f 3e 42 40 34 36 2d 26 0a 12 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 08 15 17 22 2b 29 39 3a 3d 4a 44 3d 44 37 3f 32 34 3f 3a 4b 43 42 39 3d 3b 3c 40 3a 3e 3a 43 37 46 3a 45 3d 3c 43 47 48 4b 4e 44 47 45 3d 4e 45 46 47 4c 41 48 44 47 47 47 3d 4e 3f 42 44 47 42 46 50 4f 57 49 4e 55 52 52 4d 49 49 4c 51 4e 58 4f 55 53 4f 57 50 52 55 57 5f 5c 58 50 54 55 53 52 4b 48 48 47 4f 38 2d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 2f 35 4f 3c 42 3c 3c 42 3e 42 45 45 3d 41 3d 3e 41 3c 4a 41 43 42 3e 47 3d 41 42 42 44 45 3e 41 3f 41 4d 45 41 49 4d 3d 41 47 49 44 43 47 42 44 42 4b 45 40 43 41 47 45 4a 55 52 4b 4c 56 49 4d 4b 48 47 3b 43 42 40 49 45 3e 4b 39 3d 44 3d 37 2f 26 23 12 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 11 19 20 29 26 31 40 44 55 4e 46 45 3c 45 33 3e 3d 3c 45 45 3d 38 48 3c 3a 3e 3b 49 42 48
 36 3c 3d 3f 45 44 3c 47 4f 4a 51 4a 48 4c 4c 49 49 43 42 47 4a 45 42 4e 4c 45 45 42 46 48 4b 3f 48 4b 45 4e 45 4b 4f 54 56 4d 4f 46 50 4f 4d 53 57 56 56 56 53 5b 5a 52 57 5e 5a 58 56 5b 5a 56 4c 4f 4e 50 50 4c 4a 45 31 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 2d 3f 42 40 43 45 44 41 41 47 44 49 43 3b 46 3b 3f 3e 41 3d 41 3f 47 3f 41 3d 3e 4a 47 3e 44 43 3d 46 49 45 3d 45 47 51 4b 49 46 44 44 4d 50 48 46 3e 45 46 43 41 4a 48 49 51 48 46 4f 4b 43 45 4f 3f 49 49 4f 48 48 48 4d 42 4b 42 40 45 38 37 32 25 22 0d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 17 1b 29 2e 2c 36 41 50 58 53 49 32 33 3b 3e 3c 3e 34 3e 3e 44 3c 49 40 44 44 44 41 3a 3e 42 3d 3f 46 3e 3b 44 41 44 44 4b 4a 42 48 48 48 45 4e 41 42 49 4a 49 47 47 45 45 42 3e 4a 45 4f 49 43 44 48 4c 54 4e 51 4f 53 4f 4f 50 4f 50 57 4f 57 61 57 57 56 58 56 58 5d 61 54 55 53 4e 55 4c 4b 4c 51 47 43 4a 2c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 25 3a 41 41 41 48 39 3d 40 37 49 42 3c 39 45 3e 3f 3c 3e 40 40 3a 3d 3e 44 3e 3c 48 46 42 45 40 46 44 4e 45 49 40 4b 4a 40 42 49 46 3b 42 45 41 40 4c 4b 48 42 44 49 45 46 55 4e 41 40 4c 48 4a 44 47 4a 3c 49 44 44 49 50 49 4e 3e 41 31 2e 39 23 1b 0f 09 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0e 0c 1e 24 2f 2e 33 43 58 5a 49 4a 3f 3c 33 41 3e 37 3a 42 45 3c 3d 45 49 3c 3f 3d 38 3e 3b 3d 40 3a 3a 45 3d 47 46 45 44 49 49 44 4a 4a 4b 4a 45 3c 4b 4b 46 51 4d 43 44 45 48 49 50 4c 3c 44 49 4a 40 47 48 47 50 53 4e 4e 50 43 52 56 52 55 56 5b 59 55 5c 51 5c 53 54 50 50 4f 52 4d 55 54 54 54 4e 46 45 27 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 1f 38 36 3d 3d 3e 3e 3f 3a 43 38 41 42 3e 3b 3c 3b 3e 38 42 39 3d 46 43 48 40 44 44 38 48 43 39 40 42 41 3e 46 41 42 45 42 44 44 46 4a 48 3a 46 49 48 40 47 4c 3f 52 4e 4f 50 54 4d 47 48 42 4a 44 48 46 3f 47 49 4a 45 45 44 43 45 36 3a 2f 2a 22 19 14 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0c 21 22 29 30 2b 36 49 4f 56 48 3e 3e 36 36 2e 38 38 3b 43 47 40 41 43 49 3f 44 44
 39 41 46 35 3e 3a 41 45 46 3e 48 49 4a 46 42 46 47 4a 4c 4b 43 45 48 41 48 42 44 43 45 44 51 38 23 32 4e 4b 45 41 40 47 4b 50 4d 49 45 49 47 4c 55 51 5a 56 51 51 53 4f 5c 56 55 53 54 5a 4c 4e 5c 57 59 59 4e 54 41 47 30 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 1c 3e 42 40 39 41 3c 39 3d 38 41 39 3e 43 42 33 42 45 3b 3b 41 3e 40 39 42 47 40 40 42 3c 3e 47 3f 4a 43 3e 39 3c 47 4b 42 41 4d 43 45 4a 49 48 4a 48 46 45 46 47 51 47 4d 50 50 50 46 47 44 40 41 4d 47 49 49 49 4f 46 3d 49 3f 3d 38 37 2e 29 1f 16 10 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 08 15 1d 25 2b 30 30 41 40 4b 4b 40 3a 3c 33 3d 3a 3e 3f 3f 40 42 3c 40 44 3f 41 3d 3c 3e 3e 40 40 41 41 43 40 44 4a 43 4e 45 3d 46 4a 42 4f 47 4c 4b 45 3e 4c 41 41 4b 41 48 44 44 48 4a 4d 44 40 46 48 47 4f 48 49 4d 49 4c 4a 45 47 4d 50 5a 5e 5d 56 5e 55 5b 59 57 4c 54 55 56 58 5a 5e 5d 50 4e 49 3c 33 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 35 3e 39 3f 40 32 3e 3b 38 40 3b 44 41 3a 3d 38 39 35 39 3f 44 3d 42 45 44 3d 3e 46 4c 45 3b 44 49 45 44 46 4d 4e 48 47 48 41 3c 4b 4b 46 41 46 3d 51 41 44 4c 57 46 50 50 4c 4f 47 4e 48 40 44 3f 4f 3e 49 39 4a 44 47 50 43 3b 38 37 25 24 1c 14 06 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 19 20 30 30 2a 38 3c 38 42 3c 3b 38 3c 3c 3c 35 3d 3a 3e 32 41 43 3d 44 3d 3f 3d 3b 3c 3a 3e 49 3c 40 42 40 3d 39 45 4c 40 43 4b 4b 4b 45 49 4b 44 45 49 4a 41 46 44 40 4f 46 42 3e 40 48 3b 42 46 3e 4d 4e 4c 4f 45 4d 4a 4e 55 51 53 53 59 58 53 5a 52 52 55 50 56 5e 4f 5a 5c 5a 5f 54 49 4f 3d 3b 29 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 15 35 46 39 3e 36 3b 37 3b 39 41 35 3f 3a 3a 3b 3d 3e 3b 3a 42 34 40 42 41 42 41 38 41 3f 44 43 41 4a 40 44 42 42 40 48 4d 3f 46 39 46 4a 49 44 44 46 47 43 44 45 51 46 4d 45 49 44 4e 3e 4a 3c 46 49 42 44 45 43 44 43 48 47 44 33 33 2c 25 1f 0f 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 0f 10 1f 28 28 30 2d 30 30 3b 34 3a 33 37 30 2f 38 3c 44 3c 41 3d 3b 3d 37 44 43
 3a 3d 49 3b 44 3d 40 3d 3d 43 3f 3f 3b 49 46 49 44 48 49 51 3f 45 3e 41 46 4c 40 3c 46 3d 44 46 46 3f 42 48 40 3f 40 44 3f 4a 53 51 4a 4a 43 49 50 57 57 5a 54 5b 52 5a 5b 54 59 60 59 59 5d 54 55 52 4d 59 52 43 53 3a 2f 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 35 3b 36 3f 3c 40 3b 3b 35 36 3d 3e 3e 3a 3c 41 40 3a 39 39 35 3a 3d 3e 37 41 42 47 46 44 44 46 47 44 3f 44 46 44 3b 48 49 47 41 46 41 40 46 4c 43 45 4f 4e 54 4b 4d 4f 4c 4a 42 3e 49 4a 44 44 4a 47 3b 47 43 44 45 4a 46 44 3c 2d 2b 1f 1e 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 11 17 25 24 2d 27 2f 36 30 30 37 34 33 33 31 3d 39 3f 34 3f 3c 3c 41 3b 42 43 42 3c 45 40 3f 3c 40 45 43 40 40 46 41 44 41 47 45 51 45 48 47 44 45 47 45 39 44 48 43 44 45 44 46 45 50 47 40 4a 44 4d 53 46 4c 4c 4b 4a 55 49 48 4a 57 59 5f 5e 5d 5b 5b 59 5a 5c 4e 55 5a 55 54 59 4d 53 4f 47 43 43 2f 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 18 29 3c 3a 42 35 44 3a 3b 3b 4c 39 38 3e 41 35 3c 38 3d 3f 43 3f 44 38 42 47 41 47 43 3f 43 45 46 42 42 43 3a 47 44 42 4e 44 42 44 4b 3d 45 4a 46 51 48 44 4d 4c 50 45 4b 4b 49 46 49 4a 44 4a 4b 4e 4a 40 49 3e 46 41 47 3d 39 36 33 2c 26 1c 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 14 1e 20 1b 2a 22 2e 3a 33 3a 33 3b 31 3a 35 3b 37 3b 38 3f 41 3e 40 3a 45 44 3a 3b 41 3e 42 43 44 39 43 45 43 41 42 3e 3f 49 42 50 48 45 49 47 44 43 48 4a 4f 3e 39 40 3f 47 46 45 43 41 43 45 46 51 44 40 46 4b 54 51 53 4f 55 58 53 50 51 56 52 55 5a 60 63 58 5b 4f 53 52 51 46 52 4e 48 4a 3e 2e 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 28 38 3b 45 37 37 38 35 39 3d 3a 3a 35 43 36 38 3d 43 3e 41 3d 3b 35 40 36 44 4b 46 4b 48 3e 4b 44 3e 46 45 49 47 48 46 42 49 49 44 4d 48 41 44 47 4c 40 46 44 50 49 47 48 44 42 48 41 45 43 43 43 4d 41 44 44 3f 49 43 3a 3f 2e 2f 24 20 17 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 18 1c 27 31 28 31 2d 30 34 34 34 36 37 2e 3d 37 44 36 3a 3d 3d 3b 39 39
 3b 3f 44 37 43 40 3f 40 43 3f 42 44 3a 41 41 42 52 46 40 4a 44 47 4d 44 50 40 3f 43 42 40 40 40 4c 3f 43 48 49 3f 44 4c 49 41 4d 44 44 50 49 53 51 4d 55 59 5d 58 5b 59 5e 56 56 55 55 55 4b 51 50 55 52 49 40 36 39 37 32 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 2c 41 35 46 44 40 37 3b 3d 3c 44 3b 3f 3c 3b 46 3a 40 3d 3a 3c 3e 3f 40 43 3c 47 41 3b 43 44 4b 4e 48 39 43 50 43 48 46 3c 4a 45 3f 4c 42 4b 48 49 4c 41 4e 4c 4f 4d 4b 4f 46 45 44 40 43 46 4b 3b 45 3f 41 42 3e 3c 3d 46 3a 32 26 26 15 0f 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 14 22 1c 24 2b 34 2c 35 34 41 30 30 39 30 3b 3b 42 40 40 40 3c 3e 3d 39 43 45 3f 46 42 42 42 41 3d 3f 42 3d 3f 47 40 44 41 42 49 4b 43 4e 52 48 48 42 45 44 48 3f 42 40 44 41 41 45 43 44 44 47 48 43 48 4f 4c 50 50 5a 52 57 51 57 51 62 59 56 52 5b 59 59 55 53 4f 50 4a 47 48 49 4a 3e 3c 3a 27 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 2d 3b 38 39 38 38 3e 3f 3f 39 3c 43 3d 43 39 48 43 4c 38 38 41 41 3d 45 45 4b 46 3f 47 46 46 4b 45 4e 43 4e 43 4c 4f 49 49 46 4f 48 48 48 4e 49 4e 46 44 4e 42 53 4c 48 55 47 3a 40 42 51 4d 4c 43 41 39 45 42 44 45 3b 39 38 2d 26 27 17 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 14 1a 28 2a 2d 2f 2a 3c 3b 39 3a 33 3d 39 3e 3e 39 41 3d 3d 3c 45 38 3b 4c 42 44 47 46 42 43 46 43 3f 48 48 45 41 47 42 3e 40 41 3d 47 45 4b 43 43 4a 45 43 43 3d 43 4a 49 49 4a 4f 41 3f 42 43 42 4f 47 4e 4a 4f 51 4e 52 56 55 50 59 4e 56 51 52 53 53 51 4d 4d 4f 50 4e 4a 40 3f 3e 44 3f 30 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 2e 40 3c 3b 3c 3b 42 37 3d 3f 3b 45 41 45 3a 45 41 45 40 36 42 3f 3e 3e 40 48 3d 4f 47 4e 49 4e 4d 49 4c 4a 40 48 4a 4d 4b 4c 43 3f 50 4c 4c 51 4c 46 49 4b 4a 49 49 41 3d 47 43 52 41 48 46 44 3e 48 3f 3b 3f 42 4d 3a 39 3c 2b 1e 16 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 11 11 21 24 2b 2d 32 2e 42 3a 40 39 40 3a 35 3e 39 42 41 41 3d 37 3f
 48 43 40 43 40 49 43 44 3f 3c 45 48 3c 3d 46 4e 41 48 45 49 3f 47 45 45 47 42 44 47 44 41 42 43 41 45 44 47 42 42 44 46 42 44 4a 48 48 4a 4d 53 52 4a 4f 4d 4a 51 5a 4e 4f 50 55 55 50 53 41 4a 47 50 4d 43 3a 3f 36 39 34 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 2d 39 3b 37 37 3a 39 43 38 48 33 3e 41 40 40 3c 3e 3c 3b 43 3e 3c 40 44 3f 3f 3d 40 4d 46 48 4a 4c 48 51 4a 4d 52 4c 4d 4b 4b 4b 47 4b 4c 4a 47 43 44 41 4d 47 4a 50 49 49 49 40 3e 3a 41 42 47 43 45 44 44 42 4b 43 37 35 27 25 1f 11 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0b 13 1a 27 29 2c 32 33 3c 3e 44 44 3f 3c 3c 38 35 3e 3e 3c 3d 40 48 3f 3d 40 3d 3e 45 43 43 43 4a 44 3d 3a 49 4d 4a 4a 40 44 50 44 3e 4a 43 44 49 45 4b 44 46 43 4f 48 47 40 40 45 45 44 48 47 44 4a 48 48 53 44 52 4f 48 48 4f 4d 51 52 49 46 51 4b 54 4e 4f 4f 4e 52 52 47 46 3e 40 3b 36 2e 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 30 41 36 35 38 38 3c 3e 3c 3e 39 41 38 41 41 41 47 3a 3e 45 42 48 44 53 3f 45 47 4c 54 54 52 50 58 53 59 60 63 64 62 62 52 5a 54 54 57 4f 4e 52 50 54 4a 48 45 4f 4e 41 43 43 41 47 41 45 49 4a 44 51 47 49 50 3f 33 39 30 31 1e 1d 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 06 0b 18 16 24 25 2e 2c 2e 3f 45 40 3b 3d 3d 35 3c 3b 3a 3d 37 39 45 4a 4b 3b 3f 45 46 41 42 44 49 40 49 48 49 4a 49 4a 46 45 4b 41 48 47 42 46 44 41 49 45 4c 4e 4b 47 47 49 40 42 40 44 49 46 42 4a 51 4d 57 45 4f 4e 47 45 46 3a 4e 45 4c 46 50 52 4e 54 4b 46 43 4c 46 44 40 3f 40 38 3d 34 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 29 3a 39 38 3e 3e 36 3a 33 3d 3b 3f 43 40 3e 3b 43 48 3f 40 48 44 42 50 4a 4f 4d 5a 58 67 5d 6d 71 6a 72 72 72 7b 76 78 78 6d 68 5e 60 58 4a 4f 4f 4c 4b 4a 47 43 4b 47 44 42 3d 4b 46 3f 49 49 41 4e 4d 50 47 46 38 30 31 29 19 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 14 1b 1d 27 27 2b 2f 32 3e 36 3a 38 3b 38 34 39 3f 3f 3d 3e 3c
 37 43 39 3f 3c 41 42 45 47 4f 47 45 49 49 46 44 41 41 4f 4d 47 48 48 40 3d 42 39 41 3d 46 40 45 46 43 43 44 41 49 44 4c 45 44 4a 50 49 4f 4c 4d 48 40 44 3e 42 43 3e 42 46 4c 54 4a 4d 4f 51 49 51 43 4d 38 37 3b 3b 31 2c 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 1e 3a 31 39 36 3d 39 35 3b 3d 44 42 3d 44 44 40 40 40 3d 41 42 43 4c 50 49 60 61 66 6b 78 78 7e 84 84 7f 81 8a 84 87 83 85 82 7a 71 63 6e 56 4e 50 51 45 47 45 49 4c 46 41 3c 3e 3a 46 44 46 4d 4d 51 45 49 42 3a 32 27 26 28 15 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 17 19 25 1e 24 2e 33 35 42 3b 3e 42 3d 3b 40 42 37 3a 3b 35 3e 41 3a 3d 3b 3d 44 3e 49 44 4a 4c 49 4c 4a 43 45 42 4d 4a 4c 46 45 40 43 41 47 44 42 43 48 40 4a 4b 4a 4c 3c 46 47 47 4a 4a 52 50 48 4f 56 4b 52 40 44 44 44 41 3d 3a 43 51 51 50 52 4b 4b 53 4a 43 4a 3e 3f 42 3c 39 2a 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 2d 38 35 36 45 3d 3d 40 42 40 43 3d 3e 46 3e 40 42 42 40 46 40 4a 4d 58 69 67 79 78 89 8a 7f 86 85 8f 84 86 8e 88 90 89 90 8e 8d 85 79 72 68 5d 55 50 49 53 48 4a 43 3c 45 3b 3d 45 41 41 4f 57 56 56 48 44 40 36 2f 31 21 24 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 19 1e 31 29 2f 31 2c 30 3d 41 49 3c 38 43 39 40 43 38 3d 3c 45 38 45 3f 40 41 44 49 55 4a 56 56 58 56 54 4d 47 4a 45 44 4d 42 41 45 40 49 41 40 3d 42 4d 45 48 50 44 49 45 41 43 47 52 4b 54 4c 4e 51 48 46 4a 40 43 41 4b 41 42 41 3d 4d 47 47 4d 4a 55 50 4e 44 3d 3b 3f 38 3a 29 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 2b 35 35 3d 36 3e 3f 41 3e 39 34 43 3a 44 42 4b 49 4c 48 4f 51 5f 61 76 7b 80 88 8a 8d 86 8f 90 86 8b 8d 8e 96 8c 8a 8f 8a 89 84 80 81 7d 76 6c 61 5c 46 49 4a 43 3e 3a 41 41 43 4b 44 42 45 5d 59 54 47 3e 31 2f 29 25 1b 12 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0c 13 22 20 1a 20 21 2d 27 33 30 3a 45 3f 3e 35 3a 33 34 3a 3b
 43 3b 45 3f 43 45 3d 42 3f 40 55 64 63 61 5b 55 5c 46 4f 47 4a 41 41 47 41 46 46 3f 3d 3d 3e 40 47 3f 45 45 42 44 42 44 47 51 53 51 4f 4a 4a 46 3f 3a 40 3d 3f 48 3b 3c 3c 40 3b 50 4b 47 44 4c 4d 4b 45 40 42 3b 34 3a 38 26 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 2a 3d 41 40 39 40 3e 3d 35 41 43 39 44 42 47 4a 44 4a 4e 5f 6e 6f 7d 86 85 84 89 8a 8a 8f 83 81 8a 88 8b 84 8e 8f 91 80 8a 87 7f 84 81 7b 7a 7d 6b 61 54 4a 3b 45 3b 46 43 3c 46 46 3f 44 3a 49 4f 46 3e 3b 38 31 2a 25 10 12 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 1b 1a 26 2f 29 2c 29 33 3a 42 3b 3d 40 39 41 3f 39 38 3f 3a 43 41 3d 3f 43 3f 3d 4f 4e 52 64 6c 69 64 5a 51 50 47 42 4f 47 47 48 41 47 4b 3b 41 4b 43 48 44 47 48 47 44 52 50 46 49 4f 4b 54 53 4c 4e 41 45 43 3c 41 47 3e 42 44 44 43 4b 46 49 50 49 50 49 42 39 36 3c 45 3b 33 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 24 31 32 42 3d 3a 3c 3a 3e 41 46 4b 40 4b 4e 4e 58 5f 6a 7a 7b 84 88 8e 89 8a 8c 90 8c 86 7e 89 85 83 8c 86 91 8e 8b 8c 7e 82 83 7b 81 84 7f 7b 76 62 58 52 45 4a 3f 39 49 48 45 3f 3f 42 51 46 42 3d 3a 35 31 30 23 1f 15 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0d 13 17 1e 27 20 24 25 2e 32 35 3d 3e 36 37 37 3b 3c 3c 3f 41 3c 44 3c 45 3c 42 3c 4a 4e 4d 58 63 60 6c 5a 4f 4a 53 3e 40 51 45 48 51 3f 4d 45 41 3b 43 4c 41 4d 49 42 46 44 49 4e 4c 51 4e 4c 4f 4a 50 41 42 43 36 42 45 3f 3a 41 41 43 4e 42 51 4f 48 48 42 40 35 37 32 40 38 35 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 22 35 38 3b 44 3f 3f 3d 3f 42 43 4a 4f 59 5c 60 69 77 76 86 84 89 88 8b 8c 87 91 8e 88 8d 82 82 8a 84 7e 7c 84 7f 7f 80 7e 78 87 80 81 82 7c 73 76 67 48 53 44 45 47 3e 40 45 3f 42 45 48 49 41 3e 34 36 2d 2c 23 1d 17 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 1a 26 1b 2a 25 2d 2c 29 36 30 35 31 30 30 37 3c 3a
 41 38 38 3a 44 44 40 3b 41 44 48 4d 4e 58 60 5f 5b 52 49 48 3d 51 47 46 41 46 4b 45 43 41 49 42 3b 42 42 44 4c 45 45 4a 49 4d 4b 54 4f 4c 52 4b 47 3b 3d 42 3b 3d 3e 3f 3f 3b 40 43 44 4a 45 46 44 3e 3c 3e 3f 37 3e 35 2e 26 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 22 39 38 3b 48 39 3c 47 3e 46 52 54 66 67 6e 7a 81 85 79 81 87 8b 7e 8a 84 81 85 7f 82 83 7e 7d 80 80 83 7c 7e 84 7b 84 7c 7c 76 80 84 81 82 76 6f 64 52 48 4a 45 46 41 48 3e 3c 48 47 44 40 39 3e 30 2c 2c 29 1a 1a 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 1d 28 23 28 22 29 2c 31 34 36 39 3a 38 34 32 39 3f 42 3e 34 38 3e 3f 42 41 43 46 41 4c 4b 56 56 4f 4e 42 4f 43 52 47 41 40 40 3b 43 41 43 3b 43 42 3e 45 43 48 47 49 49 4a 3f 53 46 54 57 52 49 46 43 39 3d 3f 35 3c 3a 43 41 40 42 3f 42 45 42 41 3c 4a 44 3e 38 3a 36 35 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 23 3c 32 39 3d 41 46 47 4c 60 60 69 6e 7a 80 85 7f 87 85 8a 7f 84 7e 83 81 84 85 84 82 84 7b 79 84 7f 7f 77 7e 78 75 78 76 7c 75 74 7d 7d 82 74 6d 65 54 46 45 45 44 42 49 40 3d 45 43 3f 47 3e 35 2d 2f 2b 28 15 0c 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 13 19 1c 23 25 23 26 2d 2e 33 35 3b 36 34 37 3e 3b 3b 39 43 42 3b 3a 3f 40 43 45 43 47 50 46 4b 4e 53 49 4a 47 4a 49 4c 45 40 46 3f 47 41 41 41 42 48 3e 40 47 47 40 42 45 4b 4e 4d 4a 57 4f 48 4e 48 47 3d 40 40 3f 35 3a 43 3f 41 43 3c 45 40 3d 40 41 3b 38 35 3c 34 38 37 2a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 1b 3f 38 3f 3e 43 4f 5c 5e 70 72 75 86 89 91 84 8d 8b 7e 7e 7b 86 85 85 81 7e 7d 7d 81 81 7a 78 82 7d 73 7a 72 78 78 75 79 75 71 7d 78 84 7d 78 67 5c 50 4f 4c 4b 4a 4f 42 43 3d 42 3f 40 33 38 30 2e 2a 2f 1e 19 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 19 11 1e 25 21 26 25 27 2f 3e 39 33 3c 34 35 3e
 3f 38 3e 41 39 3e 44 3f 48 47 47 45 49 47 45 4d 52 4b 45 4c 4a 4b 40 3c 4d 42 45 40 3b 46 41 3e 43 45 3e 43 3d 42 3e 44 4b 3f 42 46 46 4b 4c 4d 3f 46 41 3c 46 38 41 48 3e 42 3b 40 45 43 40 3d 3d 42 3e 3e 3e 30 3c 37 2e 29 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 3b 48 4c 59 5d 60 72 76 82 7c 83 87 86 8a 83 89 7e 80 84 7b 7c 7a 81 80 78 81 78 78 78 72 71 6e 71 77 78 70 75 71 6b 71 71 77 79 7b 81 76 75 67 58 4d 4d 3f 46 40 3c 41 39 3a 38 39 33 31 2e 28 24 20 17 1b 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 08 15 1f 1e 1f 20 23 2b 33 33 30 3e 2e 2e 3a 2d 3b 39 36 39 3f 36 42 45 40 45 42 4a 3e 4c 4d 4f 46 4b 50 46 47 47 49 42 46 41 38 41 3d 41 41 41 40 3e 41 42 3e 3e 3e 3f 43 3e 4d 49 4b 56 4d 4d 41 41 38 3f 40 41 3f 3e 42 3b 41 43 3b 3a 3e 38 40 33 3b 32 36 35 32 32 28 2c 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 3e 50 5c 6b 72 74 7b 85 81 87 86 8e 83 7f 80 7a 7c 82 7f 75 73 75 78 76 74 76 7e 75 6e 74 6f 79 70 6f 69 6f 73 6e 6e 78 78 77 6f 79 74 71 75 6a 5e 51 49 3f 49 3b 40 3a 39 37 39 33 30 30 2f 26 26 12 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0d 1a 1c 21 20 29 29 28 34 35 3b 39 39 34 37 38 3e 3d 3d 3d 40 43 44 41 47 4b 4a 40 52 4a 52 4d 46 51 4b 42 4a 46 42 4a 3f 42 4b 37 40 45 40 46 47 43 3c 3e 36 45 41 41 43 46 43 40 51 52 4c 50 49 40 46 37 44 47 3c 3f 45 4a 3d 3e 44 40 3e 3d 41 3f 3d 39 31 37 38 31 30 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 2f 5b 61 76 7d 7c 85 80 8f 8c 89 83 79 79 82 76 7e 7e 75 73 6c 6f 73 78 7c 73 76 73 73 71 72 6d 6d 69 69 6c 76 71 75 6d 6d 73 73 76 7e 79 75 72 68 51 4e 43 40 40 3d 3d 3d 3e 35 38 34 2e 2c 32 2a 24 13 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 15 18 1b 1d 22 21 36 2a 2c 35 32 2b 32 3e
 35 3d 30 35 36 3e 37 44 46 42 47 44 4a 4e 4e 45 47 4b 43 45 4a 47 49 44 41 3e 3b 43 41 43 44 44 3a 46 43 43 3b 3e 41 3d 3f 38 46 3e 43 4c 49 48 4a 45 41 45 42 45 45 43 4a 42 45 3b 37 3d 3e 3d 3e 38 34 3b 35 30 38 34 31 28 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2e 71 78 86 86 83 88 82 85 79 82 7c 77 7a 7a 7d 71 6f 6c 71 6f 73 7b 69 72 70 7a 6f 6d 72 66 70 6d 64 68 73 6a 72 6e 6b 71 7a 74 76 7a 7e 77 71 5d 58 45 3b 40 3f 47 40 40 34 35 36 2f 28 31 22 21 15 14 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0c 14 14 1f 19 21 2f 29 29 32 30 3a 35 2e 39 39 3b 3b 37 42 37 3f 43 42 40 42 47 4b 44 40 41 41 41 4b 48 47 49 39 43 42 42 42 40 40 3d 43 42 3e 43 42 3b 3f 44 3c 3f 44 4a 44 41 42 48 4a 41 43 42 45 44 49 49 46 50 4c 4b 47 44 36 39 39 3a 36 36 2d 36 2c 34 35 37 2c 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 30 74 80 8b 8a 81 79 7e 85 7d 7e 76 71 78 6e 7a 6e 71 6b 6a 73 71 6e 72 65 6c 6c 67 62 6e 6e 6b 66 66 6c 6a 6b 65 69 6e 6d 76 74 74 79 76 76 6b 62 56 44 3e 37 41 43 44 40 3b 30 29 33 28 25 2a 17 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0b 0f 0a 19 22 1c 23 2f 2b 35 2f 32 38 34 41 3d 39 38 36 40 40 42 3e 44 41 44 44 4e 47 42 49 41 4a 47 42 47 44 44 47 4f 3a 44 44 3c 42 41 3d 3b 3a 44 3a 39 3c 3d 3e 3d 37 38 48 3f 47 4a 4c 44 43 42 45 49 49 45 50 4f 5c 4d 47 3a 36 3a 33 37 36 34 2c 32 35 2e 2c 2a 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2e 70 7b 82 83 75 78 7a 76 7a 75 75 7c 6f 72 72 68 6e 6b 66 72 68 6f 6e 68 6d 73 6f 75 73 6e 63 6f 6d 68 63 68 66 6d 70 70 74 79 78 80 76 72 67 61 50 48 3c 3a 43 44 3b 3d 35 31 31 2c 28 2c 25 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 10 19 20 24 27 26 2b 29 34 39 32 42
 3b 43 32 34 33 42 3a 44 3e 47 39 42 3d 49 4d 42 48 49 44 50 4a 41 44 44 47 40 44 44 3d 45 40 49 4b 3e 45 42 3a 4a 40 43 42 3f 39 44 48 42 38 3b 42 41 44 44 41 42 43 3d 53 4a 4e 49 42 44 3b 37 2d 35 35 35 34 30 2e 2c 31 2c 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2a 73 78 82 80 7e 7c 74 78 78 72 71 6d 6e 6e 71 6d 76 67 70 65 64 61 6f 62 62 67 65 6a 64 68 66 6f 6a 69 66 66 6e 64 6b 74 54 81 7c 74 7a 6b 5f 56 54 46 45 41 44 3c 3c 3a 35 28 2c 26 25 25 1c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 15 1b 17 23 27 2e 2d 2d 31 36 3f 34 30 38 33 3b 36 35 3e 42 44 4a 43 41 46 43 4d 4b 45 46 4c 44 47 39 43 41 47 45 3f 3f 42 3d 41 3e 3e 46 41 3a 37 3d 3e 41 39 3c 40 3b 3a 43 44 41 37 41 3a 40 40 3b 46 51 50 4e 41 36 36 34 34 30 34 35 35 2d 2c 2c 2b 2c 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2a 64 70 79 7b 6a 70 6f 73 72 6e 6e 6e 72 70 6c 6c 62 63 67 66 63 66 69 66 6a 5c 68 66 69 61 64 6b 61 65 6f 66 69 72 6c 76 7c 6e 75 76 6e 60 61 4f 4f 4a 44 3d 45 3e 38 3b 3a 2d 2c 25 1f 15 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 02 15 17 26 26 22 24 2e 2b 35 38 34 39 3d 35 34 41 37 3e 39 43 41 42 3c 44 40 46 4b 4e 44 42 44 4a 46 44 40 44 44 3c 42 44 48 3e 3f 3f 40 44 3f 3e 43 3d 3b 3e 33 44 41 39 37 3a 40 39 3c 3f 41 43 3e 47 43 4a 47 44 3a 3f 38 37 32 2d 2f 39 2d 2e 38 38 33 28 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 24 63 70 6d 79 66 75 6b 64 71 6a 6e 6f 69 6c 64 6b 6a 64 6a 5f 68 5f 68 5d 61 62 67 62 69 6b 68 6b 67 63 6a 6e 68 6e 67 75 73 6e 78 74 75 6a 58 59 4b 47 4d 40 3f 39 2f 2d 2d 2b 20 1c 17 17 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 12 1f 1e 25 24 2c 31 2e 35 32
 35 3c 3a 35 35 3c 33 37 39 3f 3c 44 44 3f 3e 42 47 44 42 47 3e 44 47 43 4c 3f 41 41 42 47 4b 47 41 43 40 4a 3d 3c 38 42 3b 36 3b 43 43 44 35 3c 3d 3c 36 41 42 3b 45 4c 4b 4a 57 46 47 43 3e 34 33 35 2c 30 2a 38 31 34 23 30 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 65 6f 6e 74 65 67 6c 68 69 6c 6d 66 67 65 65 68 6a 63 64 60 63 61 62 69 57 65 6c 67 65 62 66 67 64 6e 6c 68 68 67 6f 70 7c 77 7b 74 64 62 5d 51 48 46 45 3f 39 3d 2c 29 26 21 25 1f 14 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 19 18 28 23 26 29 29 2c 37 35 3f 35 3c 35 2f 3c 3f 3d 37 42 37 39 3f 40 3e 41 42 4d 3c 43 48 3a 42 3e 40 3b 40 3b 3e 45 4a 3d 3b 44 3d 38 41 3d 3d 34 42 3a 3a 41 35 43 3d 3c 33 36 3e 43 45 4b 56 54 54 4f 48 42 3b 44 37 36 2c 35 33 30 32 35 2d 28 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 56 64 6f 73 69 5f 68 65 66 65 67 65 5f 6a 62 61 66 68 64 63 62 60 60 5a 63 5d 5f 62 5b 66 64 62 66 62 64 6e 71 73 6f 70 75 74 6d 6c 5f 60 51 4d 41 42 3c 32 33 33 2f 35 2c 20 20 0d 0a 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 1b 1c 25 2e 1f 2f 2c 33 36 3b 3c 3b 43 37 3a 30 31 49 40 3f 3e 3e 40 41 40 3e 47 42 47 37 42 42 45 3d 4a 4b 49 3d 42 40 41 3c 42 47 35 3e 39 37 38 3e 38 41 37 40 38 42 38 38 43 3e 3c 4a 51 53 52 50 59 53 50 46 3a 3c 33 30 36 36 30 32 39 30 31 33 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 55 65 6f 6d 6f 63 67 6b 70 62 6c 5f 65 6a 62 67 5f 63 5e 5a 66 65 6b 5d 64 66 5d 63 67 61 6b 5f 6f 68 67 70 72 77 64 74 6f 72 70 6f 5d 52 55 49 49 43 3c 33 37 2f 2b 26 27 19 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 15 16 23 24 20 27 2e
 32 32 3d 37 3b 3f 35 3d 33 32 39 3a 34 41 3f 3f 40 41 46 48 3f 45 45 45 3d 47 3f 40 3d 38 44 3f 41 42 44 42 40 42 3d 43 47 42 43 3c 3f 44 33 3e 3e 3e 3a 44 41 4a 51 50 54 50 46 4e 47 45 45 42 3c 32 35 2b 31 34 31 32 2b 2b 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 54 64 73 66 6b 69 67 67 66 63 68 6c 65 6e 61 66 6a 60 64 63 5d 61 65 59 65 64 5e 66 62 62 63 68 71 6d 6d 6e 69 6c 6b 72 6e 6f 70 5b 54 55 43 47 4c 43 33 3c 35 2e 26 26 23 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 15 1c 1b 21 28 26 28 2f 2d 3c 3d 36 37 32 38 32 31 2e 34 3e 3e 36 3e 41 3e 3d 42 34 43 46 49 47 45 48 3e 42 41 40 3f 48 45 3c 3b 3e 40 42 42 39 3a 3a 40 3e 3f 3d 39 38 38 44 48 4a 51 4d 48 51 41 4e 44 46 42 3e 39 33 37 32 2b 2e 37 28 2b 25 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 46 54 6d 6d 5f 5e 62 67 68 5d 5b 5c 64 68 63 5e 64 64 64 61 65 5b 5a 60 5a 5e 58 62 6b 62 65 67 6d 6b 6d 68 6e 74 74 74 6d 67 60 5e 4f 45 46 44 45 39 33 35 34 2c 2f 1d 18 0e 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 10 1a 18 1a 25 22 28 2f 2b 36 37 3e 36 42 38 3d 39 3f 35 37 39 39 3a 3e 4a 38 3d 3c 30 42 3e 40 3e 3f 40 44 44 49 40 46 40 41 41 46 3e 42 43 3a 40 45 3a 3e 43 3b 3e 37 38 43 47 50 4d 4c 4f 4e 50 50 42 4e 3f 40 3d 30 2e 32 35 2c 31 2f 35 2c 23 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 10 44 67 67 68 5c 5a 5e 6a 63 61 5f 64 5c 5f 60 5e 5e 5d 64 61 65 62 5c 60 52 5a 60 67 64 66 6d 69 68 6a 6f 79 76 7b 6c 6a 6c 5b 55 4d 50 3e 3e 48 3e 3b 36 2c 29 26 1b 18 0e 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0a 18 18 19 26 27
 26 2c 2d 31 36 36 40 41 3f 42 35 3a 37 3d 3c 39 41 40 3c 40 45 39 38 3f 3b 3e 49 43 41 44 40 3a 41 41 42 48 40 42 3e 3c 46 42 42 43 38 49 37 3f 4a 40 43 51 57 54 4e 52 47 4f 47 45 46 48 4a 41 46 39 39 31 2e 30 2e 2e 30 2d 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0c 4b 69 6a 6b 60 66 66 69 63 60 62 62 64 60 68 5b 63 5c 58 53 58 5d 5b 61 5c 5e 6c 66 65 71 66 6f 6d 69 74 6c 6d 75 70 6a 69 5a 53 48 49 43 48 46 36 34 2c 2a 2f 25 1a 13 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 0f 1b 21 27 1e 26 2d 2c 38 39 36 3b 40 3f 3b 3a 35 3f 39 33 3c 39 3e 3d 34 3b 38 3b 39 43 39 3f 42 49 42 3d 3d 45 41 3b 3c 3c 42 41 46 3e 41 3f 3e 46 3a 3e 45 43 42 50 45 4f 59 48 4a 4b 49 4a 42 4d 43 3b 3b 32 2d 35 30 2e 33 32 2d 2b 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 45 5d 61 6e 68 66 64 62 48 60 5d 5e 65 5c 62 5b 59 61 64 59 65 5c 5f 5b 5f 67 67 6b 6a 69 6a 64 69 71 74 76 69 6a 66 69 61 52 4a 49 3e 43 3e 3d 35 2f 2f 24 22 1c 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 10 19 1c 21 2b 29 26 2f 31 35 36 46 3d 3f 46 3e 39 34 38 3b 38 3d 3d 3a 34 3e 3f 3a 32 37 3b 3c 3e 3e 3b 3e 3b 3a 42 3c 3b 3b 3f 42 3d 3e 40 45 49 40 45 41 40 43 42 4a 4d 4b 48 4c 41 4a 4d 45 46 43 35 30 2f 34 33 2d 36 32 2b 2d 2e 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 43 61 68 66 66 56 5a 58 61 5b 5b 62 5d 62 5d 56 60 61 5a 5c 59 52 5a 61 5b 60 6c 69 5e 68 68 6e 67 6e 70 66 6f 6f 66 5c 51 4a 47 42 41 3c 36 34 2a 29 24 1f 1e 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 0e 1f
 1d 24 27 24 27 2f 34 34 3b 44 4d 4f 42 44 37 34 42 3b 3e 3e 38 3e 38 35 41 3d 41 3e 3c 3b 3e 45 49 46 4a 42 44 3f 3d 45 3d 3e 47 42 4d 4b 46 4c 51 50 4f 4f 4b 49 44 4b 40 4a 4b 4a 41 48 44 3b 32 33 39 31 2f 2f 34 38 32 2b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3b 53 5f 6d 61 61 61 67 64 5b 5e 5e 62 5c 60 61 5f 5a 5b 54 62 5b 57 57 5a 68 60 65 67 6e 6a 69 66 74 69 6f 6b 61 53 57 51 44 45 3a 38 3f 35 2d 27 23 1d 21 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 09 11 16 1c 1f 26 26 31 35 39 3b 40 40 4a 46 45 3c 3c 32 33 36 3c 35 34 43 35 3f 3b 39 36 36 41 3f 42 47 3e 3b 44 3a 3d 3f 3f 44 41 4d 4b 4e 51 55 56 4f 53 51 45 4e 4e 51 44 49 49 45 4d 44 4d 41 3a 38 34 35 2c 34 2a 3b 35 2f 25 24 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3c 52 5d 61 5c 62 62 5a 62 60 5b 5b 62 4f 5b 5c 5a 5c 50 59 5d 5c 60 63 5d 6a 64 68 6a 69 6b 6a 74 6b 5d 70 64 68 57 49 48 46 36 43 35 38 36 28 28 20 1b 0a 07 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 11 19 1b 1d 28 29 26 26 37 36 45 42 41 3f 3e 43 39 34 31 37 3c 3e 3b 34 35 33 33 3c 3c 38 3e 3f 43 44 42 42 3a 37 40 44 44 4d 52 56 5e 59 55 51 57 4d 48 44 40 44 49 4c 4c 43 46 44 42 4b 42 45 39 31 2f 32 30 28 33 34 2b 30 23 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 38 58 66 60 57 5e 5d 54 60 5e 60 5d 60 5d 5a 5c 58 52 54 56 5a 61 60 57 65 5b 67 64 63 71 66 6d 61 68 63 62 5a 58 55 4e 45 33 3a 36 2b 2f 28 28 1f 11 12 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 07 12 14 1d 1e 2b 27 31 2d 37 3e 41 3b 3d 36 3e 38 39 39 39 3a 3d 35 3a 38 35 3a 3a 37 3d 3b 43 45 43 48 48 3c 3f 43 42 54 4b 5e 5f 5e 60 5b 5f 61 58 54 49 48 48 47 4c 46 42 49 47 42 50 41 41 35 2d 36 34 32 33 38 31 38 2e 1a 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3b 50 5a 68 62 5c 5a 5e 5b 60 5a 55 5c 59 62 5a 5a 57 54 5d 56 5c 62 5c 65 65 6a 6a 6f 6f 6c 69 65 65 62 61 56 5b 4f 4d 42 3f 3a 34 34 26 20 1f 18 09 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 15 14 16 24 2a 2b 2e 3a 35 37 3a 33 43 38 36 3d 32 38 34 3f 3b 37 33 3b 3b 3d 35 3c 3b 3f 48 48 41 46 46 43 44 4c 50 56 5f 59 61 69 67 64 5f 5d 5b 56 49 4c 42 43 4a 4f 41 42 47 49 3b 3c 3f 3d 35 30 33 32 30 35 2d 2d 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 33 50 56 66 5b 5d 63 5b 5f 52 5a 5b 5c 5d 5e 5c 4f 53 54 56 57 56 60 63 62 66 60 68 65 6e 67 68 65 67 66 63 53 54 4c 41 42 34 2e 32 2b 22 1e 15 07 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 0d 19 1f 24 23 2d 29 2c 35 34 3d 3d 34 37 31 3c 37 39 34 2a 37 39 3e 36 30 3c 36 3b 3c 41 44 42 3d 47 42 3f 4a 4f 5b 5c 65 67 5f 66 65 68 60 5a 57 4d 4a 49 42 37 3f 46 48 3c 48 49 3c 3f 3e 3a 3a 32 33 2e 33 30 27 22 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2b 51 60 61 5d 4e 59 5c 57 57 55 58 55 51 59 55 57 56 57 58 5d 5a 60 61 64 61 6c 67 68 69 65 69 63 61 54 4f 51 50 4c 45 41 35 34 23 24 25 16 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 10 19 16 1c 27 31 31 31 37 3a 36 37 35 38 3d 35 34 35 35 36 3f 36 37 34 2d 3a 38 3f 44 3e 43 44 46 45 47 55 47 4f 55 57 59 5d 5e 62 6b 66 6b 5e 5d 54 49 49 3f 3d 45 42 42 47 42 44 3f 43 3e 38 3b 2f 35 35 31 2f 2a 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2f 54 60 63 5d 59 55 60 57 5a 58 56 57 5a 5b 56 50 56 56 52 60 5e 60 61 66 63 69 67 68 6a 5d 5d 4e 4e 53 51 51 4b 3d 3f 2e 30 22 1f 1a 1a 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 09 14 1d 1a 25 28 2c 2c 30 32 34 2f 3d 33 36 33 36 37 3a 39 34 3c 35 3b 39 3b 3f 3e 3e 46 4c 3c 4b 4b 47 49 53 54 59 56 65 5a 64 62 62 69 64 59 5e 4a 44 44 3e 41 41 44 3e 3d 49 39 42 41 44 3a 3d 3d 35 2c 32 2a 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 24 50 59 63 55 57 5c 56 5a 56 5b 59 5b 59 5a 56 5b 5b 54 54 57 5b 68 65 62 62 63 62 6b 5d 55 4f 4f 50 4f 4f 46 3a 38 2e 2a 24 20 1b 15 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 15 1f 1a 25 2c 2c 39 2e 2e 39 38 3b 36 40 38 33 40 3b 3e 38 38 39 33 41 3b 49 40 47 51 47 49 51 4b 50 55 55 5b 5c 5b 60 61 5f 61 5d 5e 53 4e 44 40 3a 44 45 40 45 3e 40 40 3e 43 3e 3e 39 39 39 34 3b 2b 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 26 4e 5d 5c 5a 5d 5c 56 57 54 57 55 54 59 54 56 58 56 5c 57 59 5f 5e 62 5a 60 62 56 5d 55 4a 44 42 44 41 3c 3b 36 2e 29 24 18 11 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 02 06 0a 11 1e 19 23 28 2e 2d 37 34 34 38 3e 36 38 33 37 3c 40 39 37 36 3a 38 3f 37 3c 45 51 4a 52 5a 5a 63 58 5b 57 52 5c 58 5b 62 58 60 59 52 50 4c 48 41 39 45 47 4f 42 40 40 3f 45 3d 3f 38 41 38 45 3d 32 2a 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 23 45 57 62 5b 51 59 51 54 52 5a 5a 5f 54 5e 56 56 5f 60 52 5a 53 60 5b 5e 5d 56 55 53 4b 48 42 3d 3b 40 34 2c 30 28 21 18 11 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0f 12 16 26 29 25 37 30 34 39 38 36 37 3d 3a 43 3b 3e 35 37 3c 38 40 45 47 4a 4a 56 5f 64 60 67 64 64 64 62 5e 55 4f 55 54 4d 51 55 47 48 3e 44 41 3f 48 48 4d 40 40 43 40 3a 3f 40 40 45 41 3b 32 33 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 20 46 50 54 56 54 4e 5f 58 4c 52 5d 54 5a 5d 5a 60 5f 57 56 5c 59 57 5c 51 53 5b 45 43 3c 42 31 39 37 31 32 35 29 20 0e 10 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0f 14 22 20 26 23 30 2e 37 38 33 3a 3c 3c 43 35 39 3a 34 38 3d 3f 43 46 4e 60 66 67 73 6e 66 63 6b 62 62 5f 58 51 48 42 45 45 4d 3d 3a 46 3a 3c 3b 45 45 42 40 3e 3c 39 3f 3e 34 42 3c 38 3a 30 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1d 42 53 55 51 50 53 56 56 50 4d 54 5a 58 59 51 59 58 58 52 53 55 59 4d 47 42 4a 41 3f 39 39 2d 38 2b 25 25 21 1d 10 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 09 15 1e 24 24 2a 38 30 36 39 34 38 40 3c 36 34 33 3b 41 3f 3f 41 47 52 66 71 6c 6a 71 6f 71 77 6c 69 55 5a 55 4d 4e 4d 3e 45 3b 3f 41 44 3b 3c 3e 41 43 43 3f 3e 3b 45 36 38 45 35 34 30 2b 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1e 47 54 5d 54 53 4d 52 4b 54 58 55 52 5a 50 4a 4c 59 58 4e 4c 47 51 48 3f 3e 41 3d 3c 39 35 36 30 22 1f 21 1d 0d 03 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0a 08 11 22 1f 22 2f 2d 35 30 3a 3a 36 38 3a 42 41 3e 3b 3b 4b 4c 59 5c 6d 71 70 7d 73 79 72 6d 73 6e 62 60 4e 46 44 3f 3e 41 3e 3c 45 45 49 44 46 43 35 3f 3b 3d 3c 3d 38 46 47 36 3e 36 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 41 4e 59 57 4b 58 4f 54 53 50 52 55 51 52 54 4e 4b 4a 50 4c 41 3d 3c 40 3a 38 39 32 28 29 23 18 25 1f 12 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 11 0f 21 20 22 23 27 30 2c 35 42 3a 3f 38 3a 39 3f 3b 44 49 49 4c 67 64 6d 6f 6d 76 75 76 6f 70 63 60 55 4d 4c 41 44 43 37 3f 39 38 40 42 3d 31 34 3c 39 44 39 3c 34 3f 42 33 3a 38 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 32 59 58 48 4c 4a 4c 55 59 51 4d 4f 4e 4d 49 4c 4f 44 40 45 38 3b 3e 32 38 35 2b 2a 25 1e 27 16 13 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 12 1d 28 2d 2d 29 2a 2f 35 3a 39 3c 38 3c 3b 44 4a 51 53 54 5e 67 6d 74 6c 68 6e 69 73 6b 65 59 55 45 44 44 41 35 3d 41 44 48 3d 39 3b 37 36 39 38 35 31 3a 3a 31 35 2c 2a 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 39 44 43 4c 42 42 4a 44 47 50 43 43 4b 42 4a 4c 42 3e 33 3a 2e 38 30 2a 2a 2e 26 22 28 1b 1c 17 0b 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 18 17 22 24 28 2f 31 38 33 2f 35 37 43 3d 3e 45 48 4f 54 5e 62 67 61 6e 6f 6c 71 73 68 64 5e 59 4c 46 44 3d 32 3c 3e 45 43 38 3c 33 38 34 36 33 34 38 3b 3a 30 32 2f 33 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2f 43 44 40 41 42 42 43 42 3e 45 42 45 30 42 3d 3a 3b 3b 32 3b 2f 1e 2d 25 2d 20 1d 1a 14 0e 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 0b 19 12 1e 2a 27 30 29 2f 2d 33 36 3d 3d 45 45 40 4c 50 5b 65 62 61 6b 68 63 68 69 6a 65 5a 50 47 42 43 3e 3c 3a 41 3d 35 41 34 31 35 2f 2b 2f 26 33 2e 35 2f 3b 33 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 25 39 3f 34 3a 3e 39 3e 3a 3a 36 3c 3c 39 38 36 2c 31 35 2c 2a 25 24 25 1f 21 1b 18 10 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 0f 14 0e 1d 1d 20 28 2e 22 28 3b 35 37 3a 44 47 48 44 4d 56 58 59 62 65 6a 5f 65 5e 5f 57 4b 46 44 3d 3b 3f 3d 36 3e 3b 3d 32 39 2c 2a 2d 2e 32 2e 26 32 27 2d 29 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1c 37 36 28 37 38 30 3e 36 2e 2f 32 34 2d 31 3a 20 29 29 27 1b 21 16 11 15 0f 11 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0c 0c 11 17 18 23 30 2d 32 25 2b 2d 3a 3b 38 3a 45 4c 4c 50 56 55 51 5d 5b 61 5d 57 51 4d 48 44 3e 38 41 35 41 3c 31 37 30 36 2a 2e 28 2c 2e 25 2c 28 27 25 26 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 20 31 35 32 2d 32 35 3a 2d 33 26 2a 2c 2e 2e 26 23 24 1f 1c 1d 1c 15 12 0c 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 09 09 18 1e 1a 25 2b 32 28 2c 30 35 3a 3b 38 3c 3c 45 47 49 49 40 46 50 4a 41 46 3f 44 3c 3b 3e 3d 2f 3a 30 31 32 27 28 25 2d 29 20 29 1d 24 23 20 24 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 22 20 18 1e 1b 2a 21 20 23 28 1e 17 1d 1e 1f 1a 1e 12 18 13 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 14 0b 14 1e 29 1e 22 2b 22 27 2b 2a 36 32 34 37 2e 2f 28 33 2f 2e 32 36 3a 3b 3a 34 36 2a 2e 30 21 2a 2b 28 24 1f 1e 24 1c 1b 20 1c 1b 15 16 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 14 0e 0f 13 10 10 11 10 0e 0a 1d 14 0c 13 0d 0a 06 08 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 09 16 16 15 23 1f 2d 27 21 27 2a 26 23 24 16 1a 15 20 20 20 22 30 38 30 32 32 27 2f 26 27 23 25 29 23 1a 1a 17 14 19 17 16 19 15 0d 11 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 05 0e 06 11 0a 0d 05 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 04 13 17 1d 1d 1f 1c 1c 1c 14 0f 10 09 07 0a 15 0f 19 16 24 25 26 23 17 17 1a 16 0d 19 12 0e 18 11 10 0f 11 09 0b 0f 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 04 06 06 05 0c 0b 06 05 03 00 06 05 06 04 0d 0b 10 11 08 0c 0b 02 06 0d 0a 10 06 06 09 00 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
