 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 05 05 05 05 05 05 06 06 06 06 06 06 06 06 06 05 05 05 04 04 04 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 07 07 07 09 09 09 0d 0d 0d 0c 0c 0c 0f 0f 0f 0f 0f 0f 15 15 15 11 11 11 0c 0c 0c 0b 0b 0b 05 05 05 04 04 04 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 05 05 05 06 06 06 09 09 09 0d 0d 0d 12 12 12 1a 1a 1a 1c 1c 1c 23 23 23 27 27 27 27 27 27 27 27 27 1e 1e 1e 14 14 14 0b 0b 0b 09 09 09 07 07 07 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 0d 0d 0d 10 10 10 12 12 12 22 22 22 2d 2d 2d 46 46 46 5b 5b 5b 87 87 87 87 87 87 b4 b4 b4 ad ad ad 66 66 66 39 39 39 28 28 28 1e 1e 1e 18 18 18 10 10 10 0c 0c 0c 08 08 08 07 07 07 04 04 04 04 04 04 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 03 03 03 04 04 04 07 07 07 09 09 09 10 10 10 16 16 16 28 28 28 32 32 32 79 79 79 a6 a6 a6 e1 e1 e1 f2 f2 f2 fe fe fe fe fe fe ff ff ff fe fe fe de de de b2 b2 b2 79 79 79 44 44 44 45 45 45 3f 3f 3f 2e 2e 2e 23 23 23 17 17 17 0f 0f 0f 09 09 09 09 09 09 07 07 07 05 05 05 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 06 06 06 0c 0c 0c 11 11 11 18 18 18 2e 2e 2e 66 66 66 5e 5e 5e 80 80 80 a5 a5 a5 f7 f7 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 f2 f2 a9 a9 a9 97 97 97 8b 8b 8b 81 81 81 7a 7a 7a 68 68 68 57 57 57 4c 4c 4c 3e 3e 3e 35 35 35 1b 1b 1b 0b 0b 0b 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 0a 0a 0a 15 15 15 21 21 21 33 33 33 52 52 52 97 97 97 ac ac ac ad ad ad c5 c5 c5 da da da fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f4 f4 d5 d5 d5 c6 c6 c6 b6 b6 b6 ac ac ac a2 a2 a2 90 90 90 7e 7e 7e 75 75 75 6f 6f 6f 6c 6c 6c 69 69 69 45 45 45 24 24 24 14 14 14 09 09 09 05 05 05 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 08 08 08 10 10 10 25 25 25 44 44 44 73 73 73 9e 9e 9e b4 b4 b4 b7 b7 b7 c0 c0 c0 cf cf cf e4 e4 e4 f6 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe f8 f8 f8 ec ec ec dc dc dc d1 d1 d1 bb bb bb ab ab ab 9e 9e 9e 92 92 92 87 87 87 79 79 79 73 73 73 67 67 67 4e 4e 4e 2f 2f 2f 16 16 16 09 09 09 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 0c 0c 0c 1b 1b 1b 3d 3d 3d 73 73 73 9c 9c 9c a3 a3 a3 b2 b2 b2 c4 c4 c4 d5 d5 d5 e1 e1 e1 ef ef ef fc fc fc fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f8 f8 f8 ee ee ee e0 e0 e0 d7 d7 d7 d0 d0 d0 c9 c9 c9 bc bc bc 9f 9f 9f 83 83 83 76 76 76 6b 6b 6b 6c 6c 6c 52 52 52 2a 2a 2a 0e 0e 0e 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 14 14 14 31 31 31 5f 5f 5f b2 b2 b2 c6 c6 c6 9b 9b 9b ac ac ac c4 c4 c4 df df df fa fa fa fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe fd fd fd fc fc fc f5 f5 f5 e5 e5 e5 ca ca ca ad ad ad 98 98 98 83 83 83 76 76 76 73 73 73 70 70 70 5e 5e 5e 3d 3d 3d 15 15 15 08 08 08 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 06 06 06 16 16 16 35 35 35 6f 6f 6f a3 a3 a3 cf cf cf cf cf cf d7 d7 d7 de de de e1 e1 e1 f1 f1 f1 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f6 da da da c5 c5 c5 b3 b3 b3 a4 a4 a4 96 96 96 86 86 86 7c 7c 7c 72 72 72 6b 6b 6b 78 78 78 43 43 43 1c 1c 1c 0b 0b 0b 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 07 07 07 18 18 18 39 39 39 68 68 68 87 87 87 99 99 99 b1 b1 b1 bb bb bb bb bb bb d2 d2 d2 f7 f7 f7 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd ed ed ed da da da c4 c4 c4 b0 b0 b0 a1 a1 a1 99 99 99 8f 8f 8f 82 82 82 78 78 78 71 71 71 9c 9c 9c 8c 8c 8c 4f 4f 4f 23 23 23 07 07 07 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 11 11 11 38 38 38 72 72 72 6c 6c 6c 72 72 72 80 80 80 8c 8c 8c 9d 9d 9d b8 b8 b8 d8 d8 d8 fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f2 f2 f2 ea ea ea db db db c4 c4 c4 af af af a7 a7 a7 9b 9b 9b 90 90 90 7d 7d 7d 72 72 72 79 79 79 82 82 82 96 96 96 53 53 53 1c 1c 1c 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0a 0a 0a 22 22 22 58 58 58 7c 7c 7c 68 68 68 73 73 73 82 82 82 92 92 92 ab ab ab cd cd cd ed ed ed fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fd fd fd fa fa fa ec ec ec d7 d7 d7 c4 c4 c4 b7 b7 b7 a4 a4 a4 91 91 91 87 87 87 7c 7c 7c 6e 6e 6e 70 70 70 9b 9b 9b 77 77 77 2d 2d 2d 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 16 16 16 3e 3e 3e 61 61 61 73 73 73 74 74 74 83 83 83 90 90 90 a5 a5 a5 c1 c1 c1 e0 e0 e0 f9 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fb fb fb ef ef ef db db db c8 c8 c8 b8 b8 b8 ab ab ab 9d 9d 9d 8c 8c 8c 76 76 76 6f 6f 6f 70 70 70 6e 6e 6e 82 82 82 43 43 43 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 3e 3e 3e 7e 7e 7e 80 80 80 6b 6b 6b 7d 7d 7d 90 90 90 a3 a3 a3 b9 b9 b9 cf cf cf ec ec ec fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fa fa fa fc fc fc f2 f2 f2 e6 e6 e6 d8 d8 d8 c6 c6 c6 b5 b5 b5 a4 a4 a4 92 92 92 84 84 84 7e 7e 7e 7d 7d 7d 72 72 72 61 61 61 73 73 73 51 51 51 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 10 10 10 61 61 61 9c 9c 9c 74 74 74 75 75 75 8c 8c 8c a1 a1 a1 b3 b3 b3 c0 c0 c0 d2 d2 d2 e9 e9 e9 fa fa fa fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 ef ef ef ed ed ed e9 e9 e9 d8 d8 d8 cc cc cc bf bf bf ad ad ad 9d 9d 9d 96 96 96 90 90 90 88 88 88 81 81 81 75 75 75 64 64 64 70 70 70 4e 4e 4e 08 08 08 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 05 05 05 17 17 17 78 78 78 a5 a5 a5 71 71 71 84 84 84 99 99 99 aa aa aa b6 b6 b6 bf bf bf d0 d0 d0 e2 e2 e2 f5 f5 f5 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fb fb fb f2 f2 f2 e7 e7 e7 e2 e2 e2 dc dc dc d4 d4 d4 c9 c9 c9 bc bc bc b8 b8 b8 af af af a8 a8 a8 a3 a3 a3 96 96 96 84 84 84 7a 7a 7a 77 77 77 69 69 69 79 79 79 4a 4a 4a 05 05 05 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 14 14 14 83 83 83 a3 a3 a3 80 80 80 90 90 90 9e 9e 9e ad ad ad be be be c5 c5 c5 cf cf cf dd dd dd ea ea ea f4 f4 f4 fa fa fa fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f6 f6 f6 e7 e7 e7 db db db d2 d2 d2 cb cb cb c5 c5 c5 bd bd bd ba ba ba b1 b1 b1 aa aa aa a3 a3 a3 9a 9a 9a 96 96 96 8c 8c 8c 7e 7e 7e 79 79 79 75 75 75 6c 6c 6c 83 83 83 3b 3b 3b 04 04 04 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 14 14 14 85 85 85 9b 9b 9b 88 88 88 94 94 94 9d 9d 9d a9 a9 a9 b7 b7 b7 c2 c2 c2 ca ca ca d3 d3 d3 da da da e3 e3 e3 ed ed ed fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f2 f2 f2 e4 e4 e4 d4 d4 d4 ca ca ca c5 c5 c5 bd bd bd b5 b5 b5 af af af aa aa aa a5 a5 a5 9e 9e 9e 99 99 99 95 95 95 94 94 94 8a 8a 8a 82 82 82 80 80 80 7e 7e 7e 70 70 70 8c 8c 8c 39 39 39 05 05 05 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 05 05 05 19 19 19 8e 8e 8e 9a 9a 9a 8b 8b 8b 94 94 94 9c 9c 9c a7 a7 a7 ac ac ac b8 b8 b8 c4 c4 c4 c8 c8 c8 cb cb cb d3 d3 d3 dc dc dc ed ed ed fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f9 f9 fd fd fd fd fd fd f2 f2 f2 de de de d0 d0 d0 c4 c4 c4 bc bc bc b2 b2 b2 a5 a5 a5 9b 9b 9b 95 95 95 97 97 97 99 99 99 97 97 97 8d 8d 8d 8c 8c 8c 8f 8f 8f 8a 8a 8a 83 83 83 85 85 85 80 80 80 6e 6e 6e 92 92 92 50 50 50 08 08 08 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 06 06 06 27 27 27 9d 9d 9d 95 95 95 90 90 90 96 96 96 98 98 98 9e 9e 9e a7 a7 a7 af af af b8 b8 b8 c1 c1 c1 c8 c8 c8 c5 c5 c5 cb cb cb dc dc dc ea ea ea fc fc fc ff ff ff ff ff ff fe fe fe e2 e2 e2 af af af b7 b7 b7 b0 b0 b0 94 94 94 7f 7f 7f b5 b5 b5 e5 e5 e5 d6 d6 d6 c8 c8 c8 bb bb bb b3 b3 b3 a8 a8 a8 9e 9e 9e 93 93 93 87 87 87 7e 7e 7e 7a 7a 7a 7f 7f 7f 8d 8d 8d 81 81 81 80 80 80 83 83 83 81 81 81 7d 7d 7d 80 80 80 77 77 77 6f 6f 6f 90 90 90 6a 6a 6a 15 15 15 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0b 0b 0b 38 38 38 a6 a6 a6 90 90 90 8f 8f 8f 91 91 91 92 92 92 9a 9a 9a a3 a3 a3 aa aa aa ab ab ab b1 b1 b1 c3 c3 c3 bf bf bf be be be cb cb cb d5 d5 d5 ed ed ed fe fe fe fe fe fe fa fa fa 76 76 76 4b 4b 4b 68 68 68 8a 8a 8a 52 52 52 3b 3b 3b 7c 7c 7c c9 c9 c9 be be be b4 b4 b4 ab ab ab a2 a2 a2 98 98 98 8d 8d 8d 82 82 82 76 76 76 71 71 71 6e 6e 6e 6f 6f 6f 7a 7a 7a 75 75 75 74 74 74 74 74 74 76 76 76 78 78 78 77 77 77 72 72 72 71 71 71 7c 7c 7c 83 83 83 2a 2a 2a 05 05 05 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 0e 0e 0e 45 45 45 b0 b0 b0 8b 8b 8b 86 86 86 8a 8a 8a 8a 8a 8a 93 93 93 9d 9d 9d a3 a3 a3 a2 a2 a2 a0 a0 a0 ab ab ab b6 b6 b6 b4 b4 b4 bc bc bc c3 c3 c3 d2 d2 d2 ed ed ed f1 f1 f1 de de de 60 60 60 2e 2e 2e 4c 4c 4c 73 73 73 38 38 38 26 26 26 5c 5c 5c b4 b4 b4 ab ab ab a4 a4 a4 a1 a1 a1 94 94 94 8a 8a 8a 7f 7f 7f 75 75 75 6c 6c 6c 67 67 67 66 66 66 69 69 69 6f 6f 6f 6c 6c 6c 6a 6a 6a 6d 6d 6d 70 70 70 73 73 73 73 73 73 73 73 73 6f 6f 6f 70 70 70 8b 8b 8b 41 41 41 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 03 03 03 0f 0f 0f 4f 4f 4f b2 b2 b2 86 86 86 7e 7e 7e 82 82 82 86 86 86 91 91 91 98 98 98 99 99 99 96 96 96 93 93 93 95 95 95 a9 a9 a9 a6 a6 a6 ac ac ac b4 b4 b4 bd bd bd d6 d6 d6 d4 d4 d4 c5 c5 c5 52 52 52 1f 1f 1f 35 35 35 58 58 58 22 22 22 1c 1c 1c 45 45 45 a1 a1 a1 9a 9a 9a 94 94 94 94 94 94 87 87 87 7d 7d 7d 74 74 74 6b 6b 6b 65 65 65 60 60 60 61 61 61 64 64 64 6a 6a 6a 65 65 65 62 62 62 66 66 66 6a 6a 6a 6b 6b 6b 6c 6c 6c 6d 6d 6d 6a 6a 6a 68 68 68 83 83 83 52 52 52 09 09 09 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 13 13 13 55 55 55 af af af 83 83 83 79 79 79 7e 7e 7e 86 86 86 8f 8f 8f 8f 8f 8f 8e 8e 8e 8c 8c 8c 88 88 88 88 88 88 9c 9c 9c 96 96 96 a4 a4 a4 a9 a9 a9 b1 b1 b1 be be be b5 b5 b5 b0 b0 b0 55 55 55 15 15 15 25 25 25 40 40 40 15 15 15 13 13 13 30 30 30 8d 8d 8d 8a 8a 8a 8b 8b 8b 8a 8a 8a 7f 7f 7f 75 75 75 6f 6f 6f 69 69 69 62 62 62 60 60 60 62 62 62 65 65 65 65 65 65 60 60 60 5f 5f 5f 60 60 60 65 65 65 65 65 65 64 64 64 67 67 67 65 65 65 66 66 66 77 77 77 5f 5f 5f 0c 0c 0c 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 13 13 13 57 57 57 a6 a6 a6 82 82 82 72 72 72 76 76 76 7c 7c 7c 86 86 86 88 88 88 83 83 83 82 82 82 7f 7f 7f 7c 7c 7c 8e 8e 8e 83 83 83 91 91 91 97 97 97 9f 9f 9f a5 a5 a5 a0 a0 a0 9d 9d 9d 56 56 56 0c 0c 0c 16 16 16 2e 2e 2e 0b 0b 0b 0a 0a 0a 21 21 21 7c 7c 7c 80 80 80 83 83 83 83 83 83 75 75 75 6f 6f 6f 6b 6b 6b 67 67 67 63 63 63 5f 5f 5f 61 61 61 68 68 68 5e 5e 5e 5c 5c 5c 5c 5c 5c 5e 5e 5e 5f 5f 5f 5e 5e 5e 5f 5f 5f 60 60 60 60 60 60 63 63 63 6b 6b 6b 61 61 61 0c 0c 0c 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 12 12 12 56 56 56 98 98 98 77 77 77 6d 6d 6d 6f 6f 6f 74 74 74 7f 7f 7f 7e 7e 7e 7b 7b 7b 79 79 79 75 75 75 74 74 74 7f 7f 7f 79 79 79 7e 7e 7e 83 83 83 89 89 89 92 92 92 91 91 91 90 90 90 53 53 53 08 08 08 0b 0b 0b 1d 1d 1d 06 06 06 07 07 07 15 15 15 70 70 70 77 77 77 7c 7c 7c 80 80 80 6f 6f 6f 6c 6c 6c 68 68 68 65 65 65 61 61 61 61 61 61 6a 6a 6a 62 62 62 5d 5d 5d 5c 5c 5c 5a 5a 5a 5a 5a 5a 5c 5c 5c 5a 5a 5a 5a 5a 5a 5d 5d 5d 5e 5e 5e 5d 5d 5d 5f 5f 5f 61 61 61 10 10 10 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0d 0d 0d 55 55 55 8c 8c 8c 69 69 69 6a 6a 6a 70 70 70 70 70 70 76 76 76 76 76 76 73 73 73 72 72 72 6e 6e 6e 6d 6d 6d 73 73 73 75 75 75 71 71 71 77 77 77 7c 7c 7c 81 81 81 87 87 87 8e 8e 8e 58 58 58 05 05 05 06 06 06 0d 0d 0d 05 05 05 05 05 05 0e 0e 0e 68 68 68 74 74 74 76 76 76 7c 7c 7c 74 74 74 6b 6b 6b 66 66 66 66 66 66 64 64 64 68 68 68 6a 6a 6a 60 60 60 5a 5a 5a 5a 5a 5a 5a 5a 5a 5e 5e 5e 5f 5f 5f 59 59 59 56 56 56 59 59 59 58 58 58 5c 5c 5c 5c 5c 5c 5b 5b 5b 0e 0e 0e 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 07 07 07 47 47 47 81 81 81 60 60 60 66 66 66 6e 6e 6e 70 70 70 6f 6f 6f 6d 6d 6d 6b 6b 6b 69 69 69 67 67 67 66 66 66 69 69 69 6f 6f 6f 6e 6e 6e 6d 6d 6d 72 72 72 75 75 75 7f 7f 7f 8f 8f 8f 5c 5c 5c 04 04 04 04 04 04 05 05 05 03 03 03 03 03 03 08 08 08 63 63 63 75 75 75 74 74 74 77 77 77 79 79 79 6e 6e 6e 66 66 66 67 67 67 6b 6b 6b 69 69 69 68 68 68 61 61 61 5c 5c 5c 59 59 59 5a 5a 5a 5c 5c 5c 5f 5f 5f 58 58 58 53 53 53 54 54 54 53 53 53 58 58 58 5a 5a 5a 4f 4f 4f 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 05 05 05 2f 2f 2f 7a 7a 7a 5d 5d 5d 60 60 60 67 67 67 69 69 69 69 69 69 66 66 66 61 61 61 61 61 61 62 62 62 5f 5f 5f 61 61 61 77 77 77 75 75 75 67 67 67 6a 6a 6a 72 72 72 73 73 73 7c 7c 7c 5c 5c 5c 04 04 04 03 03 03 04 04 04 03 03 03 03 03 03 05 05 05 57 57 57 6e 6e 6e 6f 6f 6f 76 76 76 7d 7d 7d 79 79 79 75 75 75 71 71 71 72 72 72 6f 6f 6f 6e 6e 6e 69 69 69 5e 5e 5e 57 57 57 5a 5a 5a 5c 5c 5c 5c 5c 5c 5a 5a 5a 55 55 55 54 54 54 50 50 50 59 59 59 55 55 55 32 32 32 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 16 16 16 6a 6a 6a 5c 5c 5c 5a 5a 5a 5d 5d 5d 64 64 64 64 64 64 62 62 62 5e 5e 5e 5c 5c 5c 5e 5e 5e 5d 5d 5d 5b 5b 5b 6c 6c 6c 6a 6a 6a 6a 6a 6a 6a 6a 6a 6d 6d 6d 69 69 69 72 72 72 5c 5c 5c 04 04 04 04 04 04 03 03 03 03 03 03 03 03 03 04 04 04 4a 4a 4a 65 65 65 6c 6c 6c 6f 6f 6f 71 71 71 6f 6f 6f 6d 6d 6d 6d 6d 6d 70 70 70 6c 6c 6c 64 64 64 66 66 66 69 69 69 5c 5c 5c 57 57 57 59 59 59 5b 5b 5b 5b 5b 5b 57 57 57 54 54 54 55 55 55 5b 5b 5b 4e 4e 4e 16 16 16 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 0d 0d 0d 44 44 44 5b 5b 5b 56 56 56 58 58 58 5e 5e 5e 62 62 62 5e 5e 5e 5a 5a 5a 58 58 58 59 59 59 5a 5a 5a 5e 5e 5e 5b 5b 5b 56 56 56 5b 5b 5b 62 62 62 63 63 63 65 65 65 68 68 68 57 57 57 04 04 04 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 42 42 42 5f 5f 5f 62 62 62 64 64 64 64 64 64 68 68 68 68 68 68 66 66 66 66 66 66 63 63 63 62 62 62 61 61 61 65 65 65 62 62 62 58 58 58 58 58 58 5a 5a 5a 5a 5a 5a 58 58 58 56 56 56 54 54 54 56 56 56 41 41 41 09 09 09 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 0d 0d 0d 2b 2b 2b 54 54 54 56 56 56 56 56 56 59 59 59 5d 5d 5d 5b 5b 5b 59 59 59 57 57 57 58 58 58 5d 5d 5d 5f 5f 5f 55 55 55 53 53 53 53 53 53 55 55 55 5b 5b 5b 5e 5e 5e 60 60 60 52 52 52 06 06 06 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 34 34 34 55 55 55 56 56 56 58 58 58 5d 5d 5d 5f 5f 5f 62 62 62 63 63 63 60 60 60 5e 5e 5e 5d 5d 5d 5c 5c 5c 5c 5c 5c 62 62 62 58 58 58 5a 5a 5a 5c 5c 5c 5c 5c 5c 59 59 59 58 58 58 52 52 52 52 52 52 29 29 29 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 1f 1f 1f 46 46 46 52 52 52 55 55 55 55 55 55 5b 5b 5b 5a 5a 5a 57 57 57 58 58 58 5b 5b 5b 5d 5d 5d 59 59 59 53 53 53 4e 4e 4e 4e 4e 4e 50 50 50 51 51 51 56 56 56 57 57 57 4f 4f 4f 08 08 08 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 2b 2b 2b 4e 4e 4e 4f 4f 4f 53 53 53 58 58 58 58 58 58 5e 5e 5e 5d 5d 5d 5a 5a 5a 57 57 57 58 58 58 59 59 59 59 59 59 61 61 61 58 58 58 5a 5a 5a 5d 5d 5d 5a 5a 5a 56 56 56 56 56 56 4f 4f 4f 47 47 47 11 11 11 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 18 18 18 3b 3b 3b 4e 4e 4e 52 52 52 56 56 56 58 58 58 58 58 58 58 58 58 5c 5c 5c 5d 5d 5d 5b 5b 5b 56 56 56 4f 4f 4f 4e 4e 4e 4c 4c 4c 4e 4e 4e 4e 4e 4e 52 52 52 52 52 52 4b 4b 4b 0a 0a 0a 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 24 24 24 49 49 49 4b 4b 4b 4f 4f 4f 54 54 54 55 55 55 57 57 57 57 57 57 55 55 55 52 52 52 55 55 55 56 56 56 57 57 57 5b 5b 5b 57 57 57 5c 5c 5c 5c 5c 5c 59 59 59 55 55 55 50 50 50 4d 4d 4d 35 35 35 06 06 06 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 12 12 12 35 35 35 4d 4d 4d 50 50 50 55 55 55 5b 5b 5b 58 58 58 59 59 59 5e 5e 5e 5e 5e 5e 5b 5b 5b 57 57 57 4f 4f 4f 4d 4d 4d 4c 4c 4c 4b 4b 4b 4c 4c 4c 50 50 50 4e 4e 4e 4a 4a 4a 0c 0c 0c 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 1e 1e 1e 49 49 49 4b 4b 4b 4e 4e 4e 52 52 52 55 55 55 54 54 54 52 52 52 55 55 55 54 54 54 54 54 54 59 59 59 54 54 54 58 58 58 58 58 58 5b 5b 5b 5b 5b 5b 57 57 57 51 51 51 51 51 51 49 49 49 24 24 24 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 2d 2d 2d 46 46 46 4b 4b 4b 4e 4e 4e 56 56 56 59 59 59 60 60 60 64 64 64 5f 5f 5f 5d 5d 5d 54 54 54 4f 4f 4f 4d 4d 4d 4a 4a 4a 4a 4a 4a 4a 4a 4a 4b 4b 4b 4b 4b 4b 45 45 45 0f 0f 0f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 19 19 19 45 45 45 47 47 47 4b 4b 4b 4e 4e 4e 51 51 51 50 50 50 4f 4f 4f 53 53 53 53 53 53 55 55 55 56 56 56 55 55 55 57 57 57 57 57 57 5a 5a 5a 59 59 59 55 55 55 51 51 51 4d 4d 4d 41 41 41 12 12 12 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 22 22 22 4a 4a 4a 45 45 45 47 47 47 4b 4b 4b 55 55 55 5f 5f 5f 5b 5b 5b 5d 5d 5d 5c 5c 5c 56 56 56 50 50 50 4d 4d 4d 4c 4c 4c 4a 4a 4a 4a 4a 4a 49 49 49 49 49 49 42 42 42 11 11 11 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 12 12 12 43 43 43 45 45 45 49 49 49 4d 4d 4d 4d 4d 4d 4f 4f 4f 52 52 52 57 57 57 54 54 54 51 51 51 57 57 57 58 58 58 56 56 56 56 56 56 59 59 59 5b 5b 5b 5c 5c 5c 50 50 50 48 48 48 30 30 30 06 06 06 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 14 14 14 3a 3a 3a 40 40 40 44 44 44 49 49 49 4d 4d 4d 56 56 56 57 57 57 58 58 58 59 59 59 55 55 55 4e 4e 4e 4d 4d 4d 4a 4a 4a 48 48 48 49 49 49 47 47 47 47 47 47 41 41 41 15 15 15 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 0f 0f 0f 41 41 41 41 41 41 47 47 47 4b 4b 4b 4f 4f 4f 50 50 50 55 55 55 55 55 55 51 51 51 52 52 52 58 58 58 54 54 54 53 53 53 55 55 55 5a 5a 5a 55 55 55 4e 4e 4e 49 49 49 45 45 45 1b 1b 1b 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 2e 2e 2e 3d 3d 3d 40 40 40 47 47 47 46 46 46 4b 4b 4b 4e 4e 4e 4f 4f 4f 4f 4f 4f 50 50 50 4c 4c 4c 4c 4c 4c 4a 4a 4a 4a 4a 4a 49 49 49 47 47 47 45 45 45 3f 3f 3f 16 16 16 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 0c 0c 0c 43 43 43 46 46 46 4a 4a 4a 4d 4d 4d 4f 4f 4f 4f 4f 4f 4e 4e 4e 51 51 51 4e 4e 4e 50 50 50 55 55 55 4f 4f 4f 51 51 51 50 50 50 54 54 54 4a 4a 4a 46 46 46 45 45 45 39 39 39 09 09 09 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 22 22 22 3a 3a 3a 3c 3c 3c 45 45 45 45 45 45 45 45 45 46 46 46 47 47 47 4a 4a 4a 4a 4a 4a 49 49 49 49 49 49 45 45 45 48 48 48 48 48 48 48 48 48 45 45 45 40 40 40 18 18 18 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 09 09 09 45 45 45 4b 4b 4b 4a 4a 4a 4d 4d 4d 4b 4b 4b 49 49 49 46 46 46 48 48 48 47 47 47 4b 4b 4b 4e 4e 4e 4c 4c 4c 4d 4d 4d 4c 4c 4c 49 49 49 46 46 46 46 46 46 43 43 43 24 24 24 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 15 15 15 31 31 31 38 38 38 3e 3e 3e 40 40 40 41 41 41 3f 3f 3f 42 42 42 45 45 45 43 43 43 46 46 46 46 46 46 46 46 46 45 45 45 44 44 44 46 46 46 44 44 44 40 40 40 1c 1c 1c 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 06 06 06 42 42 42 45 45 45 45 45 45 45 45 45 45 45 45 44 44 44 40 40 40 44 44 44 46 46 46 4a 4a 4a 49 49 49 4c 4c 4c 4e 4e 4e 4b 4b 4b 47 47 47 4b 4b 4b 49 49 49 37 37 37 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 28 28 28 36 36 36 3b 3b 3b 3c 3c 3c 3d 3d 3d 3f 3f 3f 41 41 41 40 40 40 40 40 40 42 42 42 44 44 44 47 47 47 44 44 44 40 40 40 3d 3d 3d 3f 3f 3f 3e 3e 3e 1e 1e 1e 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 39 39 39 3f 3f 3f 3f 3f 3f 3e 3e 3e 3f 3f 3f 3f 3f 3f 3f 3f 3f 45 45 45 48 48 48 4b 4b 4b 4b 4b 4b 47 47 47 50 50 50 58 58 58 63 63 63 67 67 67 51 51 51 1c 1c 1c 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 2f 2f 2f 3a 3a 3a 3b 3b 3b 3f 3f 3f 3c 3c 3c 3c 3c 3c 3e 3e 3e 41 41 41 47 47 47 48 48 48 58 58 58 43 43 43 3b 3b 3b 39 39 39 39 39 39 37 37 37 1f 1f 1f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 37 37 37 3e 3e 3e 3f 3f 3f 3f 3f 3f 41 41 41 40 40 40 43 43 43 42 42 42 42 42 42 48 48 48 48 48 48 4d 4d 4d 69 69 69 7a 7a 7a 71 71 71 61 61 61 31 31 31 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 24 24 24 36 36 36 3c 3c 3c 41 41 41 3e 3e 3e 39 39 39 37 37 37 3c 3c 3c 3d 3d 3d 3e 3e 3e 44 44 44 3c 3c 3c 39 39 39 35 35 35 37 37 37 37 37 37 22 22 22 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 31 31 31 41 41 41 41 41 41 43 43 43 46 46 46 43 43 43 3d 3d 3d 3b 3b 3b 3e 3e 3e 44 44 44 4c 4c 4c 6b 6b 6b 7e 7e 7e 73 73 73 63 63 63 47 47 47 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 2d 2d 2d 38 38 38 44 44 44 41 41 41 38 38 38 37 37 37 36 36 36 35 35 35 36 36 36 35 35 35 39 39 39 36 36 36 35 35 35 32 32 32 31 31 31 21 21 21 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 27 27 27 41 41 41 3d 3d 3d 3d 3d 3d 3d 3d 3d 3c 3c 3c 3a 3a 3a 3c 3c 3c 41 41 41 59 59 59 76 76 76 7a 7a 7a 6c 6c 6c 5f 5f 5f 4b 4b 4b 1a 1a 1a 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 1b 1b 1b 2d 2d 2d 3e 3e 3e 3d 3d 3d 3a 3a 3a 39 39 39 38 38 38 35 35 35 37 37 37 32 32 32 31 31 31 2f 2f 2f 2e 2e 2e 2f 2f 2f 2d 2d 2d 21 21 21 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 1d 1d 1d 38 38 38 30 30 30 30 30 30 31 31 31 33 33 33 34 34 34 42 42 42 5f 5f 5f 6f 6f 6f 6b 6b 6b 5f 5f 5f 56 56 56 47 47 47 21 21 21 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 1e 1e 1e 2c 2c 2c 32 32 32 34 34 34 35 35 35 35 35 35 35 35 35 40 40 40 2e 2e 2e 1e 1e 1e 10 10 10 1b 1b 1b 1b 1b 1b 17 17 17 0f 0f 0f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 08 08 08 0f 0f 0f 0e 0e 0e 0e 0e 0e 0f 0f 0f 13 13 13 19 19 19 27 27 27 27 27 27 28 28 28 23 23 23 21 21 21 1d 1d 1d 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 15 15 15 1d 1d 1d 1d 1d 1d 17 17 17 16 16 16 0d 0d 0d 14 14 14 0f 0f 0f 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
