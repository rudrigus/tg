 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 06 05 03 0c 08 05 05 06 07 05 05 09 13 11 14 12 08 10 15 13 0d 1f 33 3a 2e 12 0c 10 10 1a 1f 22 1e 12 0c 0c 12 05 0c 09 0c 0e 0a 0d 14 13 19 1e 16 17 13 1e 14 21 28 1d 15 12 0d 0d 06 05 05 01 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 0b 00 06 05 03 0f 0c 0a 0e 10 0f 09 11 1b 17 10 13 0f 19 1c 2d 42 3e 32 35 24 2f 38 30 2e 26 35 3b 47 39 2e 21 20 2c 2d 32 33 25 27 1e 26 1d 20 25 26 26 29 23 2d 34 36 31 39 35 1f 1f 2b 30 2a 2c 31 31 25 15 14 15 11 0c 12 06 05 03 00 07 0a 07 0c 06 06 08 08 06 05 03 00 06 05 03 05 06 05 03 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 03 06 05 03 01 06 05 04 03 08 10 0e 00 06 08 07 0a 0e 0a 19 13 14 13 10 20 22 19 12 14 1e 38 42 62 7a 64 3b 34 2b 36 3a 35 40 51 54 58 54 44 3e 4e 4c 48 3e 41 44 3e 35 3b 37 2e 3a 3b 3a 46 41 3f 4d 4d 4b 48 33 36 2f 31 2f 34 34 39 2f 34 27 27 1b 24 1c 17 1d 11 10 0a 0a 0f 08 0a 06 05 0a 0d 06 06 03 05 06 05 03 00 06 05 08 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 08 09 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 03 06 07 03 07 06 05 0e 0a 08 0c 03 0c 14 1d 15 18 20 11 14 20 1e 1e 22 32 48 60 83 ac b3 84 59 39 36 34 3d 56 6e 84 84 7e 73 68 6d 76 6a 63 61 60 69 5c 5b 56 59 59 58 61 6b 6f 6a 64 6e 6d 69 64 4b 46 3b 35 3b 3d 36 39 39 42 40 38 39 37 36 37 2b 22 1f 20 19 1f 12 1b 16 14 2b 20 0c 0d 06 0a 0f 05 08 01 06 06 03 07 06 08 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 11 09 07 07 0c 03 06 05 09 0d 17 10 09 10 10 10 13 18 16 17 29 42 43 39 47 4f 61 73 99 a6 9a 88 73 50 48 50 5d 6c 7f 84 81 75 64 74 6f 85 87 87 8b 89 82 84 89 7b 86 8e 89 99 9b 9f 9f 8d 95 8f 9b a0 84 4e 44 3e 42 3f 3f 46 42 48 56 59 56 56 52 55 49 4f 3c 3a 35 33 2c 26 1e 26 36 31 1f 1c 0b 0f 0d 05 03 06 06 09 0b 0e 06 06 06 06 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 0e 0f 0c 07 0c 1f 13 20 13 15 1b 18 20 2f 35 39 3a 45 58 64 6a 53 59 6b 70 6f 6d 6d 5c 68 57 57 5e 5a 5f 67 6e 65 69 66 66 7f a0 b6 bd c3 b8 b6 ba b8 bc b7 c2 c3 d1 d7 d3 ca c4 b6 ad ae c0 a2 84 6d 5c 50 4b 4f 51 56 64 6d 67 74 76 7a 74 71 6a 5a 69 5e 53 42 49 34 35 33 31 13 26 20 1d 1f 15 14 13 11 09 13 10 0e 06 05 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 09 03 00 06 05 04 01 06 05 03 00 06 05 04 09 06 05 0c 09 07 13 18 20 18 19 1e 1c 24 24 2b 30 41 45 50 5e 60 58 69 63 76 64 59 5d 5e 64 5f 61 67 5a 5d 61 5f 60 57 67 67 6a 67 6a 66 6f 78 92 b3 cc d9 df da d4 d2 d7 d5 db e5 e8 e6 e4 d8 d1 bc b7 b4 a4 95 96 8c 8b 7d 80 81 7a 8a 89 8a 87 87 95 94 99 9a 9a 8e 8e 85 7e 76 6b 65 52 56 4f 54 49 37 2d 37 2e 20 1f 1c 1a 14 16 19 13 11 12 0d 05 07 06 06 05 04 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 07 0e 05 07 03 06 0d 09 03 06 0d 15 12 1b 29 2a 2a 2d 29 36 3c 3d 42 4f 5b 5d 5a 5d 68 66 6c 6a 6c 62 61 64 58 64 64 64 6d 70 67 69 6c 66 6b 6d 71 6d 76 73 75 77 75 77 7b 8b 99 ad be c1 c6 c9 ca d1 df e6 df e9 d9 d7 de cb bc 9e 89 85 81 81 7f 7e 7f 7d 83 89 8d 94 8c 90 9d a1 a3 a3 ac ac b3 af ab a0 9b 8a 7c 75 74 6d 6b 68 5e 5a 54 47 3e 3a 32 2c 23 25 1b 1c 15 0d 13 17 09 0d 05 06 05 06 05 08 01 0e 17 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 09 07 06 05 0b 08 0d 0b 03 0d 0e 10 18 2d 34 34 43 43 43 50 52 55 62 63 6a 61 5d 67 52 5c 5d 63 5c 66 64 5d 5f 5a 69 6a 6b 6c 71 6d 74 72 74 78 74 75 78 83 7c 80 7d 7e 76 7b 86 8f 90 a2 aa ae c0 d0 d3 d7 e4 e6 e3 e8 d6 d2 bf a0 86 89 7c 84 79 82 7e 73 7c 7c 7c 7e 7c 7c 84 81 88 8b 95 9a ae a8 a7 b5 ad a8 a5 a0 9c 9a 92 8f 8a 87 7a 71 67 5b 62 4e 49 46 34 36 30 20 2d 1d 13 0f 12 0b 0f 06 08 0c 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 09 06 05 0e 06 11 0f 19 1b 13 10 10 1d 17 2d 43 52 55 61 5f 70 73 6e 6e 6b 65 63 61 64 5c 60 64 64 68 70 6f 69 67 6c 6f 72 6f 78 7c 74 7d 7f 84 84 75 80 83 85 8d 8a 90 91 8c 91 8e 90 97 93 9b a0 a9 bf c2 d8 da de ec e9 ee e4 db c3 a8 94 87 92 8e 8c 87 88 8a 7f 88 86 84 89 87 80 85 84 7e 80 7a 7f 80 81 8a 87 8c 93 95 8e 8a 9d 99 a4 a8 ad ac 97 92 89 7b 79 71 64 4f 54 41 45 41 38 2b 20 2e 22 17 18 11 15 14 0d 13 06 03 03 06 0d 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 0d 0b 0b 17 11 21 1f 27 28 24 28 2e 3c 4d 6d 77 79 73 76 7d 66 6b 6a 65 60 6c 6a 67 6a 65 6c 6e 6d 75 74 79 73 73 82 7b 7e 7c 7f 87 87 8a 87 8f 88 90 97 97 96 9f 9b a4 a4 a5 a3 ae aa a4 aa b3 b7 c5 d3 d6 de e9 f7 f9 ee df ce b1 9d a5 a0 9f 9d 97 8a 95 98 92 91 97 90 97 99 9a 92 91 8e 84 83 7b 80 7a 78 76 70 76 7e 75 73 78 7a 8b 91 9a a4 a8 a2 a3 9d 95 8c 6c 74 63 62 5f 5e 4f 52 4e 43 40 39 2a 2d 2e 22 21 17 0a 0d 08 0b 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 05 06 06 17 19 17 1b 1e 23 21 28 2b 31 49 50 56 5a 72 7a 7a 7a 6b 6b 6a 60 61 62 64 68 67 63 71 6e 6f 65 76 7b 74 7a 81 7e 7c 83 85 86 87 8c 8f 9a 9c 96 99 98 98 9d 9c 9f 9d a4 a6 ad ae b9 b6 bd b5 c6 c4 cc d3 d4 de e0 eb f1 f9 ee e2 d3 ba ad b3 ac ac b1 a9 ae a3 a2 a3 a2 98 98 9f a4 9f a1 9e 95 92 8d 89 86 7e 7c 7b 76 77 73 6a 70 70 73 71 6b 71 6a 73 7e 8c 8d 87 84 81 7b 70 75 73 73 7a 77 6a 69 5e 57 4d 40 3b 3a 35 2a 1a 20 0d 0d 06 0e 09 0b 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 05 09 0d 05 03 07 06 0e 0d 10 1a 15 1d 1c 25 28 2e 3d 4a 48 4d 52 63 60 5f 6a 6a 6f 6c 63 65 64 60 5c 64 64 67 6e 6e 78 6f 75 77 73 7f 84 83 83 86 8e 8e 8a 92 8a 97 90 98 9b 99 9c a0 a9 a6 a5 af ac b7 b4 c0 c3 c5 c8 d5 d5 d6 d9 d6 de e2 ea e9 f2 f9 fa f4 ee d9 cb bf b6 b0 bf b6 bd b6 b9 a7 af af af b0 a6 af aa ac 9f a5 a0 99 99 96 95 7f 86 7e 75 79 78 70 76 6d 77 6d 6b 6a 6d 70 6c 69 69 6b 69 6f 67 67 68 60 65 6e 79 81 83 76 71 65 67 54 4a 49 42 33 26 1c 0a 0f 0a 10 0c 09 07 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0a 0a 05 08 15 0c 15 1b 22 2b 2f 32 2f 3c 43 52 64 6e 64 58 52 56 55 5a 64 60 5d 62 65 6f 68 63 6f 6e 76 71 79 77 72 7a 73 7b 7e 89 87 90 91 95 99 94 9c 9f 9d 9f 98 9c 9b ac ab b3 b1 b6 bc bf c1 c9 c5 d6 d1 e1 eb e7 ec e8 f1 f4 ff fa f7 fd ff f8 ff f5 ea df c4 c0 c3 c5 bf c6 c4 b7 c0 b5 b8 c0 b3 b6 b4 b5 b3 b0 a9 aa a3 a4 ab a0 99 8d 85 87 80 84 7f 71 7f 72 74 74 73 69 6d 71 65 6c 6b 6a 66 6f 63 5c 5e 61 61 67 68 6a 75 86 7e 78 7f 6d 6c 67 51 47 31 29 21 11 1c 12 0b 0c 10 07 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 05 0e 0c 12 17 1c 18 1c 25 2b 39 3e 4a 4d 45 54 5b 65 6c 60 56 56 53 57 5a 5d 5c 5a 69 6d 72 71 6c 6f 73 71 75 79 7c 7e 78 7e 7e 84 8e 91 92 94 a7 9c 9d 9f 9e a1 ac ac af b1 b4 bd bb ba bb c7 c8 ce dc e7 e8 f1 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 da d8 c8 cd cb c9 d0 cf c9 c8 c8 c9 bf c0 bf bd b3 b8 af b4 b8 ac aa aa a3 a0 9c 8e 8f 97 87 87 85 80 7c 75 7c 7f 74 7a 76 73 75 77 71 75 72 68 64 72 60 66 5f 5c 5d 5e 6b 77 7b 84 8b 7d 75 6a 4c 42 38 2e 2a 30 2a 1b 1a 15 0c 11 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 09 06 05 03 00 06 05 07 07 07 0c 0e 14 14 1b 28 2c 34 34 3b 46 5a 51 52 53 5a 60 61 63 5e 59 61 5d 62 66 6b 63 6a 71 73 6e 79 75 7f 7e 75 80 85 87 8a 84 87 91 95 92 98 8f 91 a4 9c 9e a6 b0 af aa b3 af c0 bd ca c6 c1 c9 d7 df e4 ea f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd e7 e4 d0 db dd da e1 dc d0 d0 cd cf c9 c1 ce c7 c2 c2 be b4 b6 bb b2 b2 a4 a5 a3 a5 98 99 97 92 96 84 92 8e 80 86 85 88 8b 85 88 7d 7b 82 85 72 76 70 78 6f 6e 61 65 65 65 63 69 76 80 7a 86 73 65 59 46 35 3b 3f 33 2f 29 21 0e 0e 0a 0a 06 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 02 06 05 03 02 0a 0e 08 14 0d 1b 1a 21 2c 2a 37 47 47 52 56 5c 68 67 67 58 5f 62 5f 6b 58 64 5e 66 64 78 6b 7b 75 84 7f 7a 85 7f 88 84 8e 90 8a 8a 8f 8a 99 8d 9c 93 98 a6 a4 aa b3 af b5 b2 b8 ba bb c0 c8 c9 cf d6 e3 e0 e9 f3 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ed e4 ec e6 e6 e3 e0 db e5 da d9 d3 d3 cc cc cd c4 c9 c2 c3 b8 c2 b6 b4 b7 b2 a9 ae a6 a4 a4 9c 9d 9d 9c 96 9a 8f 91 8b 98 91 8e 94 8c 8f 89 85 79 7a 80 78 6e 64 68 64 5d 61 56 54 6c 6d 67 64 5b 4f 56 51 58 59 46 30 20 1f 24 18 16 0b 07 09 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 09 0b 09 14 0d 14 22 1f 2c 32 3a 45 46 52 5e 6b 69 65 67 79 73 64 6b 66 62 60 60 64 6e 6e 70 75 77 74 7b 82 87 89 8c 88 87 93 8f 8f 94 8d 96 93 96 92 a0 95 a4 a4 9f ae a8 be bc c0 c3 c1 bf ca d5 d1 db e1 e7 e7 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f2 ef f0 eb e6 e6 e2 e5 e0 de d6 d7 d2 d1 d0 ce ca d2 cc cb c5 c2 b9 bc b7 b5 bc b6 b2 b0 af b0 ae a2 a6 a8 a9 9f a4 a1 94 9e 95 96 9b 93 8a 8b 81 7a 79 7b 76 69 61 5f 5b 5f 56 60 5e 5f 5c 54 58 55 54 65 61 58 4b 41 3a 38 2b 26 17 1a 0a 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 01 06 05
 03 07 06 05 0c 13 15 20 26 2e 3a 4f 51 5f 64 70 77 73 77 6f 74 70 6a 5c 5e 63 68 6d 6a 6c 70 71 77 7e 86 7d 7c 82 8a 8c 8e 93 94 95 96 94 95 98 99 96 9c a1 a2 a7 a7 ab b2 af b7 b9 bd c4 cb cf d5 d3 d4 d6 e0 e4 e8 f9 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f2 f8 f2 ec e7 eb e1 e0 e1 db e1 d5 e2 d6 de db cf d2 ca cd d0 c9 c5 c4 c8 cb c5 c5 c4 b8 bb b9 b9 ae b9 b2 aa b4 a0 ab a2 a8 a2 a8 94 94 91 90 88 82 79 77 6e 6c 64 5d 5e 5b 60 5b 58 57 5c 55 50 5d 5f 5c 5d 55 4e 4a 4c 41 34 2a 20 18 13 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 09 10 10 0d 18 14 24 27 36 3d 4b 57 63 6b 75 81 82 81 7f 75 72 6d 69 69 67 6c 6f 73 6c 71 75 7e 7a 7f 80 86 88 8b 92 93 8a 98 8f 9e a1 9b 9f 9e 9f 9e a1 a6 b0 a5 ae b3 b6 bd b6 b6 c5 c5 ce dc d4 e4 dc e0 ec f3 ed fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 f2 f1 e4 e8 e4 e1 dc e4 ec e5 e5 e0 d8 d5 d1 d7 d8 d4 d1 d4 d3 cf d2 d8 d0 d0 c9 c5 c8 c7 c2 bb c0 af b8 b1 ac ac a8 a8 a0 a2 9d 9d 8e 86 8c 85 7b 7a 74 6d 68 6c 5d 65 6f 68 68 62 60 5d 5e 5c 5f 57 65 5c 57 6c 67 48 40 2c 1f 20 0f 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 07 03 0a 07 16 18 22 25 35 38 49 57 66 6c 76 72 76 78 84 75 72 63 62 66 63 68 6a 6f 72 76 76 80 80 7c 83 81 7f 84 8e 92 9a 94 96 98 97 9f 9e 9d 9f a1 a8 a8 aa ae af a8 bb b6 b6 be be bf ca cd d0 d8 d8 de e4 df f1 ef f6 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 ec ef e6 e6 e9 e3 e8 e9 ee ef e4 e1 dc df da d4 db d2 d7 d9 d5 d9 d1 dc d3 d4 d2 d6 d3 c6 cc ca c7 c4 c2 b6 b7 af b3 ae a9 a0 9b a2 94 94 91 87 7e 7e 77 75 70 6f 6f 6a 6e 6b 68 69 6b 65 5c 60 64 67 60 5b 64 74 79 69 4a 3f 29 28 1f 0e 08 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 06 0f 0d 14 19 1e
 23 30 39 41 4a 66 71 79 7b 86 86 80 7b 74 6d 6b 6a 62 6d 6f 71 74 77 7b 7e 84 7d 85 85 82 85 92 93 97 97 a1 99 9f 9c a7 a9 a6 a4 a5 a1 a9 a7 a8 b2 ad b6 b4 bb c0 c4 c3 c6 d3 d6 d4 dd dd e4 e4 eb f2 f4 ed f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ef f2 ef ec e7 ea ec e7 f2 ec e5 db dc d9 e2 e0 e1 df df e5 e3 e2 de e2 e1 dd dd d4 d9 d6 cc cc c4 c8 c0 bd bf b7 b3 b2 b0 ac a3 a2 9a 95 8f 91 85 7a 7b 7c 6c 79 79 74 76 78 77 77 6e 71 66 68 63 69 69 64 60 6b 7a 75 6f 5e 46 3a 2b 21 0d 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0c 0d 0e 13 17 1b 25 2e 36 44 52 65 72 80 8d 9a 93 8d 7d 6d 6b 67 6c 76 6d 6b 6f 6c 70 80 82 84 91 95 95 92 94 96 94 97 9c 9c a4 a5 9d a2 a5 b0 b2 ae ba ad b3 af ba ab bc bb c1 c6 c0 c5 c1 d3 cd d2 e4 e0 e4 d9 e5 e4 e7 ef f7 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ef f1 ee f4 f1 f1 e2 ed ed e6 e1 df eb e7 e2 ec e5 e4 e8 eb f0 e7 e8 eb e2 e1 e3 d5 d8 d1 d4 d2 cc c1 b9 bd b6 b7 b4 b1 a2 a2 a0 a1 96 93 8e 8f 88 84 7f 84 7c 80 7e 79 7d 6e 77 72 6e 72 71 64 5f 61 56 69 63 68 71 79 5d 43 32 27 23 0e 0f 06 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0f 0d 17 16 24 24 2b 41 3b 56 63 6d 8c 92 94 96 8b 7b 79 6c 63 6c 6a 77 78 72 78 74 7c 73 86 89 8d 94 95 91 9a 96 99 a1 99 a4 a4 a9 a8 aa a9 af b1 aa b1 ba b6 bb b7 b8 c0 bd c2 c9 cb c7 d6 cf d6 de db e4 e3 e2 e4 e6 ec f0 f3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f6 fb f5 fa f4 f3 f1 f0 ee f1 e9 e9 e7 e5 ea f4 f6 ed ea ee f4 ef f0 ef e1 e0 df ea e6 de e2 ce d5 cb c4 b9 c1 b1 b8 ad ad ab a2 a4 95 95 91 95 90 8e 95 84 87 87 85 82 80 81 73 76 71 65 6e 69 66 60 5c 5e 5e 62 68 81 68 5b 3d 2e 22 18 1c 0c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0f 05 08 0f 12 20 25 29 28 36 45 50 53 6b
 79 88 97 98 91 8a 81 72 6a 72 6f 75 74 75 7b 77 76 79 7a 86 87 8b 87 93 95 9a 9c 9d a1 a2 9a a4 a7 a4 a4 ae b2 ae b7 b8 c0 c1 be c3 ba c5 c7 c4 c8 c3 ca cd cb d8 de da e1 e2 e1 e4 e9 ec ea ef eb f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fc fe ef f8 f8 f0 ec f3 ec eb f5 f2 f2 ed e9 f7 f4 f6 f5 ef f0 e8 e2 ec ea ea df d9 d9 d7 d0 cb cc c7 bb c0 b6 a2 a8 a3 a0 a4 9b 9a 9a 8c 90 8f 90 93 87 80 82 7a 80 75 6f 65 60 67 6b 67 5d 60 5f 57 65 5a 73 80 6a 4e 39 2f 24 15 0f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 08 0d 0d 12 16 1d 20 2e 2d 36 3d 43 59 6d 6c 85 90 93 99 96 89 86 7d 72 7e 79 82 82 7e 85 8b 83 85 8c 89 8b 90 88 94 9b 9f a0 a0 a3 aa ab a6 ab ac ad a9 ab b9 b7 b2 ad be c5 cc cf ce cd cd cd cd cd d3 d5 d6 d7 dd dd db e3 e5 e4 e9 e9 ef f5 f1 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fe fb f9 fe f8 f5 f4 fb fe fe ff ff f6 f6 f7 f6 ed f5 f4 ed f4 ee e1 e1 d9 d2 cd cd c4 c2 9d b4 ab ae aa a4 a5 a3 a3 a2 94 8f 9a 9b 8f 8c 8b 79 7f 77 73 77 74 67 6a 6a 65 64 53 55 5a 61 61 74 8a 7d 62 50 43 2c 25 1c 0f 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 06 08 09 08 16 1e 24 2a 32 38 43 4d 51 58 65 7b 80 8b 9d 97 91 89 7e 79 79 7c 81 84 86 89 8f 8b 93 8c 8e 8f 92 93 94 a2 94 9b 9f 99 b1 a2 ad aa ab b2 ac b1 b1 b8 b4 c1 bf ba c6 ca ca c5 cb d0 d8 d9 d1 d7 db da d6 df d1 dd e4 dd eb e1 e7 e7 e8 ed f5 f3 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 fe ff fd ff ff ff fd ff fd fb f5 f4 f3 f4 f6 f3 eb e6 e4 de d4 cb d4 c1 bf c5 b2 b9 af aa a3 a6 a2 a7 a9 9e 9d 9b 91 8c 90 82 7c 7d 74 7a 71 75 68 69 69 64 5b 5c 5b 55 55 59 60 82 7f 74 5f 43 3a 2e 1d 0b 0b 06 03 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0d 06 0a 0a 06 15 21 22 29 3e 4b 4f 5b 57 67 76 80 96 a2 9c 90 80
 7e 76 75 82 81 83 88 8e 96 9b 93 a1 92 9a 99 9d 99 93 9e a1 9f 9d a7 a8 a7 a1 ab ad b3 b2 b3 b0 b4 b1 b9 bd b9 c0 bb c8 cc ce d9 d4 d3 d7 d5 d7 d5 d8 dd e2 d7 dc e2 e8 e3 e6 e7 e7 f1 e5 f0 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 f5 f5 f6 e9 e3 df da d7 ca ca cc bc c2 ba b6 b8 af ab 9f a7 9e 9f 99 96 90 8e 8b 90 83 81 7b 73 71 7b 71 6e 6a 67 65 5c 4c 53 51 57 58 5c 6a 81 7c 6a 52 43 31 25 20 0e 0f 00 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 0a 0d 10 0a 14 27 2f 30 41 59 68 75 7f 89 97 a6 b0 9c 85 7e 76 72 7e 81 7d 86 8f 90 97 99 a3 9d a2 9d 9f a4 a4 aa a5 a1 b0 a5 a7 a4 aa a9 a7 a9 b3 b4 c1 b9 b1 ba b6 bd c3 bb c1 cb c9 d7 d2 da db dd d5 d6 e0 e0 e0 d8 e4 e1 e1 e6 ec ee e6 f0 ed ed f5 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fa f4 f0 f3 e7 e7 e5 e0 d5 cf c6 c8 c5 bc b3 b6 b5 b1 ac a7 a0 a5 a0 9a 95 96 92 90 84 8d 88 81 89 7c 79 7c 6e 70 6b 61 5f 5f 51 59 54 51 4d 5c 6e 77 7b 65 54 39 2e 21 16 0a 06 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 0b 0e 17 14 17 1b 1f 2b 44 44 62 7f 84 98 a3 ab ad 99 84 6f 74 7d 80 88 87 93 95 9b 95 a9 a0 aa ab ab ae ad b1 a9 ad a9 af aa b0 b0 b1 a5 b5 ac ae bc b7 b4 bb c3 ba b5 c2 bf c8 cf cf d2 cb d5 d9 da de dc d6 df df e0 e3 e2 df df f0 e8 e9 ee f3 f4 f8 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa f9 f1 e9 e2 df de cd cf cf c7 c4 c0 bf b7 be ac ac a4 a5 9d 9f 9d 97 92 8d 8e 99 8e 85 85 80 81 73 7a 78 6e 66 65 5c 5a 5d 53 55 57 54 4f 57 6e 7d 71 62 42 2f 1b 19 12 09 08 0c 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0c 13 0e 19 11 1e 2f 3c 4b 60 7b 90 92 a1 9d 94 80 7e 7a 7a 7c 7d
 89 86 8e 8f 92 9c a7 a7 a3 af b1 ad b6 b7 b4 b8 af bb ae b1 b9 ac b4 af b0 b0 ae ae b7 b4 b8 be ba bd be c4 c1 c9 d4 d5 d7 e0 e1 d9 e0 df da e1 e2 df e6 e5 e4 e9 ef ea f4 f0 f6 f3 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fd f2 f6 e6 ed ea e0 e3 d0 cd cd cb cb c7 b5 bf b7 b1 ae b2 a6 a7 9f 97 9b 94 9c 93 9b 91 8f 84 81 7f 78 71 73 6d 65 65 62 58 5b 51 5a 53 52 5a 56 57 6d 68 56 46 3e 37 1c 12 11 0b 0d 06 0e 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 0b 0b 0c 1b 1d 1d 2d 3b 53 60 6b 7e 91 95 94 87 76 76 75 6b 7d 7a 81 85 83 93 9e 9f a0 a8 ad b0 b6 be b4 c1 b2 bb b8 c5 c0 c1 b5 bc b9 bb bb bb ba b0 bb b3 b6 b8 c0 c5 c0 c4 c8 cd d2 da d3 dc db e7 de d8 db da e3 e2 db de e1 e4 ed f2 ed f8 fd fd fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fd fb f2 f0 e9 e9 e5 e3 db d1 cf d2 c3 cb c3 be bd b0 b2 b2 af aa a0 a4 a2 a2 ac a0 97 9c 8c 8b 8f 82 7e 72 71 75 6a 60 61 59 5f 55 5b 55 50 56 59 50 5d 51 57 57 51 3f 27 13 06 0b 05 0c 04 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 0f 10 1e 23 31 30 47 55 65 78 84 7f 81 7e 7f 75 7a 70 75 74 7c 7b 7f 82 90 96 95 9c a2 a8 b4 af b7 bf c0 bd c2 ca c5 c8 c3 c1 bb bf c8 c2 c4 c3 bb bc be be b4 bb ba c5 c9 bf c5 cd cd d9 d2 d7 e2 e0 e5 dd e3 e1 e3 de ea ea ea e9 ea ee f0 f5 f9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f8 f3 f5 ea e8 eb e7 dd d6 cd d1 d4 d6 c9 c8 c2 ba b9 b5 bb b0 ad a8 af aa a2 a6 a3 96 94 91 88 7d 7b 7b 6c 73 71 6d 65 5f 5d 5c 5e 54 5c 53 57 52 51 58 5c 71 5c 44 2c 1e 10 08 09 0a 01 0b 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 14 19 24 36 44 54 5f 74 76 77 7a 74 6e 6e 77 75 74 76 76 7a 7c 7d 88 8e
 95 94 99 a1 a4 a5 ad b0 b4 bd bc c4 c8 be cf c6 c0 c7 cc c6 c7 c6 ca cb ca bd c7 bb c3 c0 bd ba c9 c9 ce cc d1 e0 d6 e4 dd e2 e5 e7 e0 e4 e1 e6 ed e7 ed ed ec f5 fc fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 f1 f8 ef e4 e7 e8 e3 e0 df d2 d9 d5 cd ca cc c6 c0 c4 bc b7 bd b1 b1 aa aa 9e a5 9d 94 8f 8a 7d 7e 82 79 7d 77 72 66 64 60 55 58 54 54 57 54 54 5a 59 70 7d 64 57 41 26 18 0a 08 0d 0b 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 09 11 21 23 2d 42 50 6a 73 81 6c 6e 5f 67 6f 65 6b 72 71 72 73 7e 85 83 8f 91 94 95 9a 9b a3 a8 ae b1 b2 bb b8 c4 c4 c4 c3 c6 cd cf c9 d2 cc d1 d2 c9 cc c8 c5 c9 c5 c6 ca c7 cb ce d0 da df da dd dc ec e4 e5 f4 ef e5 e9 ee ed e1 ee f4 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc ff ff f8 f8 f4 eb e7 e9 e8 e9 df d9 dd e0 d2 d2 d4 d0 c4 c9 c4 c5 c0 b9 b4 b1 ac ab a8 a2 9b 98 8f 87 84 80 82 7b 7a 72 67 63 5b 50 65 5c 5d 50 52 52 5f 63 80 86 7a 57 3b 36 2b 1a 1a 12 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 08 09 06 13 19 2a 30 3a 52 60 71 88 8a 6b 68 5e 65 69 69 6f 78 75 7f 83 84 84 90 8b 94 a0 9f 9d a3 a9 a5 ae b4 b2 ba ba bc c4 c3 ca cf cd cb d4 d7 d3 d1 db d2 d2 d0 d6 d4 d7 cf d4 d3 d5 d5 dd e0 df e3 e3 e9 eb e9 ea f6 f2 ee ef f3 f4 f4 f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff fc f9 f7 f9 f8 f6 e6 ec e5 e6 e6 e4 e1 dc d6 cd ce ce c7 c4 c7 c7 c0 bc b2 b0 ab ab a0 9c 95 8a 90 85 86 7e 78 76 6f 65 6a 5e 64 55 5c 5c 55 51 56 5c 71 84 76 69 5c 48 37 26 15 1a 10 0c 07 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 0f 12 2b 33 30 42 58 69 7b 8f 84 64 5c 62 5e 6a 6a 6a 70 76 78 81 7c 85 89 92 91
 9e 96 a1 a3 a4 a3 ad b1 b4 ba bc bc b9 cb c8 d4 ce cb d2 d3 d3 db dd d9 e1 d9 d9 d8 da d4 dd dc dc d8 de e1 e4 eb e7 f2 f3 f0 f2 ff ef f5 f5 f5 fe f6 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff fe ff fe fb f7 f3 f1 ec ee ea e7 e3 e2 e1 d3 d9 d4 cc d0 c6 c7 c1 c6 b7 b6 b1 b1 a5 a2 99 95 98 90 87 80 77 75 72 60 67 5c 60 56 58 5b 5e 4e 58 52 59 6c 75 72 68 51 40 3c 35 1b 0d 14 08 0d 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 1a 1d 34 3d 40 53 5a 7b 8b 8d 75 64 60 5b 65 61 67 68 74 70 78 7e 80 86 90 90 94 99 9d a7 9f a4 a2 a9 ac b6 bb b4 bd ba b6 c5 c5 ca cb d1 d4 d7 d7 dd d8 df da e1 e3 e2 e9 e4 e2 e0 e1 e0 e4 e9 f2 f2 f1 f7 fa f4 f3 de de fd fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fd ff ff fb ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fb ff fd ff fc f6 fb ef f0 eb ee f5 e0 e3 e4 d8 dc de d7 cf cd c9 c8 c5 c1 b9 bd af ac ad a4 98 99 84 85 82 7b 77 6a 65 5f 56 52 5b 5a 50 57 53 58 4f 54 58 5a 63 6c 5f 46 3a 34 24 18 12 0b 06 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0c 0b 0b 1b 21 23 32 4d 5c 66 77 86 95 88 66 63 65 64 63 63 70 74 7e 7b 78 75 7f 81 81 93 99 99 9c a0 9d a4 ac ad b0 b2 b7 b5 b9 be c6 c1 cd c7 ca cd cd d2 d4 d6 d7 d8 de e1 e6 e2 e2 eb ea f2 eb f1 f4 f2 f3 fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff fe ff ff ff ff fc ff f7 ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fb fb fe f7 f1 f0 ef e9 ec e4 dc e3 e4 de cd d0 d0 d3 c7 ba bf b8 c2 ad a8 a6 a5 9c 9a 91 8a 83 7a 6d 6b 62 63 64 5b 5c 5b 55 56 51 52 51 4b 4d 49 61 67 6c 55 38 29 28 16 16 0e 0c 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 07 12 11 18 1d 2d 3d 50 69 71 81 8a 91 75 6b 56 61 72 70 64 71 6c 68 7d 71 79 8b 84 8b 8c 8b
 9c 9d 9d 9b a4 a6 ac b2 b3 b5 b7 bd c4 c5 c6 cd cc c9 d7 de ca d8 d4 d3 dc db df e6 e4 e9 f0 eb f4 f6 f9 f8 f9 ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fe f8 fd f9 f9 f7 fa f9 ff ff fb ff ff fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fd fb f2 f5 f1 f5 f7 e5 ef e7 e3 e4 e3 dc d4 cd c9 cc c6 c5 b9 c0 b5 af ab a6 97 96 95 8b 81 79 71 6a 72 63 62 5d 57 55 54 59 52 57 4c 46 4f 50 55 62 62 5a 53 3e 2f 21 18 1f 12 08 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0b 0b 1a 17 1b 25 30 4c 5b 6d 76 84 8a 75 66 65 68 6d 68 64 68 67 6e 72 70 80 80 7f 84 8f 8a 8f 90 9f 9c a1 a6 9d a5 ad b1 b0 bd bb c4 c6 c2 cb d2 cf cc d8 da d0 d9 d7 d7 d8 dd dc e7 ec ea eb f3 f3 f2 fd fc ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 fa f7 f9 f8 f8 fa f9 ef f5 f7 f2 f9 f4 fb ff fa ff ff fd fc ff ff fd ff fc ff fc ff ff ff ff ff ff ff fd fc fd f6 fa f9 f8 ef f4 ee ea e9 e6 df e1 dd d3 d2 cd cb cb c5 c3 be b3 b6 af a5 a2 98 92 89 87 84 7f 72 69 6c 6e 69 5c 55 5d 5a 4f 51 5a 49 4d 50 51 4a 56 53 55 56 41 35 26 21 24 21 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 0b 12 1a 1f 26 32 2f 37 45 61 6e 82 7f 7d 6b 70 60 6a 64 6d 68 6d 6b 72 7b 7f 7d 80 8d 84 85 8c 82 91 9d 9b 96 9a a4 a5 ae b9 ab b7 b5 c1 c8 c9 c5 cc d0 d6 d3 d5 d9 d9 d8 d6 d2 d7 e0 d8 e0 e7 eb f0 f8 f6 f8 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ef f3 f1 f1 f0 d4 ed f0 f1 f6 fa ef fd f4 f0 f1 f6 f7 fb f6 fb ff fa ff fb ff fd fc f9 ff ff ff ff fc ff ff f9 f6 f6 f7 f3 f2 ee e8 f4 ee e9 e2 dd dc df dc d9 ca c6 c3 c6 bd c0 bd b1 ad ad a5 9b 99 8f 89 80 7f 77 71 6c 6b 5e 66 5e 66 59 60 4d 55 54 54 59 56 59 5c 5c 5d 55 54 40 30 2d 26 1a 16 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 0c 0a 1c 1f 22 29 33 36 49 4c 5d 6a 70 78 6f 6f 63 65 5c 68 68 6b 67 6a 6f 6d 77 7b 7f 8a 86 7f 8a 8f
 8c 91 91 95 9a 9d a2 a1 ad b2 b0 bd bd ce ba c9 d4 d4 dc d9 df e0 d8 df e5 db d9 e5 e1 e6 e0 ed f1 ee f5 f6 fa ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ef ef e9 ea ec eb eb f4 ea e8 e3 ec e9 ea ee f5 f5 f9 f6 f0 fb f8 fe fc fb fc ff f7 f7 ff ff f6 f9 f6 fd fa fc f6 f9 f4 f8 f0 f1 f7 ee f0 ec e6 e2 dc de d9 d6 dc d1 cb ca c9 c6 c1 bc b9 b5 b1 a5 a3 9d 99 91 8e 83 80 7d 70 70 6b 6c 65 61 5a 60 59 5f 55 5b 52 61 5c 60 5c 5e 5f 64 5b 4b 3a 39 23 21 12 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0d 16 22 26 29 2b 30 4c 4c 58 64 63 69 69 6c 62 64 5a 62 6d 68 64 66 64 6c 67 6f 6e 77 84 7a 82 84 87 8c 90 8e 92 9d 96 a4 a2 a5 ae b5 ac bb c2 c9 c7 d1 d5 cf d3 da e4 e5 e4 e0 e3 e2 e1 dd df df eb ec e5 f1 ed fb f5 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb eb e2 eb e5 e2 ed e4 ec e6 e0 e6 e2 e9 e8 e1 ea f4 f5 f4 f3 f3 f8 f4 f6 f0 fb fb fa fc f9 fe f8 f5 f8 f8 fe f4 f6 f3 f3 f2 f2 e7 e6 e2 e9 e9 ec dd e5 d8 d7 ce d9 c9 cd c6 c0 c3 b7 b0 b3 b4 b2 ab b2 9e 9c 98 8e 91 8e 86 82 75 71 6b 70 67 65 5c 5e 64 5f 5d 5a 62 60 5a 5f 63 60 5c 68 68 59 53 3d 2a 16 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 0c 19 28 33 3f 3b 45 51 5a 5d 5e 60 67 5d 62 69 5b 61 61 61 63 69 68 69 6d 6f 71 6f 70 81 7f 7d 8b 84 8c 91 8e 92 8e 96 9e a5 a7 b6 b0 b5 b9 bc c3 c8 ce cc d8 d9 da e1 ed e3 e9 e4 e6 df e9 e1 e7 ec f4 ee f0 f8 f8 f2 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ed e4 e1 dd dc dd de e4 e4 e1 e0 eb e5 e1 de e8 e8 ec ef ef de ef eb f5 fa f1 f8 fd f7 fa f3 f2 fa f8 f6 f1 f7 ef f1 eb f5 ef e4 f1 e9 e0 ea e6 e5 d8 de d3 ce ca cf c4 c4 c3 c3 c4 bc b4 b1 b3 a9 a6 a1 a5 9c 9d 93 8b 8c 89 7d 81 74 74 6d 6e 6c 66 69 70 66 65 68 67 63 66 5d 6d 6a 62 63 6f 72 52 49 36 22 16 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0d 19 1e 27 41 51 50 54 56 5b 57 5a 60 61 64 60 67 60 64 64 6b 63 68 61 66 70 6e 6e 73 73 7b 7e 83 84 89
 8a 87 88 95 97 9d a5 a5 a5 a9 a5 b8 ba b9 c7 c2 c8 cd d4 d5 dd e2 de e7 ea e5 e6 e7 ed e3 ec f3 ec f6 f6 ff fa f7 fd fa ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 e3 df db dd d4 dd d7 db e0 db d3 da d9 df e2 de db e0 e2 e6 ec e6 ef ef ee f1 f7 f1 fa ee ef fa f1 ed f1 ef f5 f4 f1 e9 e7 e8 eb e5 e8 e1 e4 e1 e8 d8 d6 d8 cf d2 d1 cc cf b5 be c5 b8 b8 b8 ae ae ab a3 a1 a1 9c 92 9a 8c 8d 81 76 77 80 72 73 74 72 75 75 67 78 71 70 6c 65 64 5c 5f 5e 67 7d 7b 62 4b 31 29 17 07 05 03 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 08 0c 1a 1b 23 38 53 66 61 60 5d 59 5d 60 64 5d 5d 67 64 60 61 61 68 64 62 67 74 6a 69 6f 73 78 73 81 7c 7b 8a 8f 8e 95 93 9b a1 a4 a1 a9 ab b2 b0 b3 b4 c0 cc c4 cb d1 d3 db d6 dd e4 e7 ea e9 e4 e8 ea f1 ef f5 f5 f7 fa f7 fa ff fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ec d6 d8 da d4 d8 d6 d6 d8 d1 d1 d2 d5 d1 d2 d5 d7 da e0 e3 e6 e7 e5 e9 e9 ee e3 f4 f1 ec f0 ec ed ea ee f4 ef f3 ec ed ec e3 ec e2 da dd df d9 d4 da d4 d5 d5 cc cd ce c6 c9 b5 b9 b0 af b8 b4 af ac a3 a6 98 91 9c 93 94 89 88 87 84 7a 77 82 7c 72 78 71 77 79 70 6d 68 66 5f 63 59 5a 63 73 83 7e 5e 3e 30 1f 15 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0c 18 13 22 28 33 4e 61 64 61 5e 56 61 60 6b 66 62 5f 64 62 64 6c 6c 64 6f 74 72 71 61 72 72 78 79 75 7e 84 87 87 8d 94 98 93 a3 a0 a2 a9 ad aa b3 b6 b9 bf c5 c1 cb c8 d1 d4 d5 da e4 de ea e7 ec e5 ed f0 e8 f0 f5 fe f5 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe e5 e5 d7 d5 d5 cf ce dc c9 cf ce cd cf d0 d2 ce d7 d7 d3 de e2 e2 e2 e5 e7 e5 e6 ed eb ee f2 eb e9 e4 e2 e6 e2 e4 e6 e4 e4 dd de e0 e0 db d7 d5 d8 d9 d3 ce d5 be c8 c7 c5 c4 bf b4 b5 b7 b8 ae b1 ab 9f a1 9d 92 99 99 95 8a 89 8a 8b 7f 81 7d 7b 84 7c 83 77 78 72 66 68 61 60 60 5b 59 66 75 96 8b 67 47 36 1d 19 0b 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 12 0f 1f 17 29 30 39 51 5c 66 5c 54 5d 5d 61 64 62 5d 6a 5e 6e 65 69 6e 68 6d 78 74 79 71 79 6e 85 87 7d 87 89
 7b 89 95 93 9b 9a 9f 95 a1 b3 af af b7 b2 b7 ba c3 cc c6 cd c8 cf df dd d5 d9 dc e4 e8 e4 ee e8 f4 ee f0 f5 fa fd ff f7 ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f4 e3 dd db d6 c9 cb d1 cb c8 cf c9 cc c6 c5 c4 cb c9 d7 cf db e3 de de dd ea e5 e7 e5 df e7 e7 f1 e2 ea e9 e3 e8 e4 e5 e3 e1 d8 d5 d4 da d6 d3 ce d5 cf c5 cb cc c7 c2 c1 be be b9 b4 b9 b5 b5 b1 a3 a0 a7 9f 99 9b 98 8b 94 8a 8a 84 85 88 88 87 86 81 77 77 70 68 67 63 5a 60 5e 60 5d 68 81 99 88 67 41 2e 25 14 12 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 0d 09 1b 26 2c 2b 2a 3c 50 5f 5f 5f 5b 58 60 5f 5f 61 60 64 69 63 6b 68 6b 75 6b 72 6e 78 72 7a 76 78 78 80 85 80 8b 8c 8b 91 95 9a 99 9f a7 a0 a4 af b0 b3 b8 b6 bc bd c7 c5 cb d6 d0 d5 dd d8 dd dc e0 de e3 e5 e4 ed ed f1 f6 ff fa ff ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 ed e3 dc ce cb cf ca cc cf c7 c9 be c3 c5 c9 c7 ce d0 d0 d2 da d9 e7 e3 de de e6 e6 de e5 e4 e9 e3 ea e5 e2 e5 df dc dd de d6 d6 d8 da d0 cf c6 d8 cd c8 c7 c3 c2 c8 bd be b8 b7 b5 b0 b2 b7 af a9 a4 a5 a5 96 95 94 94 91 8b 93 88 86 82 85 86 81 7c 78 6b 72 69 6d 64 66 5f 5f 58 62 6f 87 9a 87 63 49 32 1d 0b 07 0b 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 04 06 14 20 2d 3a 30 2d 43 4d 5e 54 62 5e 5a 5b 5e 67 5e 5e 69 64 63 63 69 6b 69 6e 68 76 7d 7f 7c 7a 84 7d 81 8b 88 90 8d 96 90 93 9f 9e 9d 9b b2 a7 ac b0 a9 ab b7 bc b8 c5 c2 c8 cf d6 ce d3 cf cf d6 de dd df e9 e3 e9 f6 ef fc f2 f6 f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e6 d2 d6 ce cb cb c8 ce c6 bf c6 c0 c5 c6 c0 bc cc cb d0 d2 d5 d6 e0 e1 df e1 e0 e1 e6 df e0 e0 df e0 d7 db e2 db d9 d2 d2 d1 c9 cd d4 cf d3 d2 cd c9 c4 c1 c5 c7 bd b8 b9 b1 bc ad ac b0 af af a3 ab a5 8f 98 8e 9a 95 89 88 8e 84 7f 85 81 7f 7c 75 71 6f 68 61 68 61 63 69 65 61 71 91 97 8f 62 44 2c 16 16 0e 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 1e 2c 3a 4c 44 44 4f 61 5b 59 5f 5c 62 60 62 61 65 5b 68 67 69 60 6f 6e 6c 6f 6d 7a 7e 7a 82 86 84 83 85 81 86
 93 8d 95 9c 95 9e 9b 9b a8 a4 a9 ad ac b6 b6 b4 c0 b4 b8 c7 c8 ca d0 d3 cd d6 d5 e1 e2 de e2 e4 e5 f0 f6 f4 d7 f0 f8 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 df cd c9 d2 c6 cc be c4 c0 c1 c6 c3 c5 c2 c4 c9 c7 c8 cc d1 d8 d0 d3 da e7 e5 de e3 d4 d9 e5 e3 de dc e2 dd d5 d8 d1 d7 cf ce cc cd d3 ca cc cb c5 c4 c9 c1 bf c2 c6 c0 b4 bb b1 b5 b7 bc b3 a8 a1 a5 9d 9f 9c 94 92 8b 94 93 8f 98 83 86 80 81 78 7c 75 6b 6f 6e 6e 66 6d 61 6a 7f 94 9e 8a 6b 43 2b 1e 0f 06 07 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0e 16 2c 3e 52 5b 62 5f 63 6b 5e 66 5f 64 64 60 62 62 63 6b 6c 67 6a 69 6c 65 6c 70 72 7e 7f 7d 7e 84 89 8b 8a 92 92 90 93 96 a2 98 9b a5 ac b0 aa ae ac ae ae b6 bb b7 b9 c5 c1 cf c5 c6 cc d0 d9 d7 d6 e1 e0 dc e3 e2 e7 ef f1 fb fa f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc e5 d0 ca d0 c4 c4 c9 c3 b8 c2 bb ba bf c1 be cb c0 ca c5 ca d8 ce e2 d3 df df db db d9 e1 e1 e4 e2 d7 d8 d8 d9 d9 d4 d2 d4 d5 ca cf ce c7 cb c7 c6 c3 c6 c1 c1 c1 c1 c1 c0 b3 b9 b5 b4 b3 ac aa ab a2 a0 9b 9a 96 96 93 92 91 8b 8d 7e 8b 7d 83 7c 82 7b 71 6d 70 65 64 6e 69 6c 76 9e a4 8a 6b 3b 29 17 11 06 08 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 08 15 28 31 43 4b 60 62 62 70 6a 65 6a 65 5e 59 5e 5f 5f 61 6b 67 69 6e 6c 70 6b 6b 6e 75 78 7e 7d 7e 80 7e 88 8e 91 95 91 90 95 99 9a a2 a6 a8 a6 a3 ae ac b0 b4 b6 b6 bb bc bb bc c5 c8 c8 ce d2 d5 cf d5 d9 e0 db e4 e5 e2 f3 ee ef fc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee dd cb cf c4 c2 c3 c1 c2 bf c1 c5 b5 c0 b5 c2 c2 c5 c6 ce c9 cd d7 d2 d7 db d9 dc db dd da da d4 d7 d6 e0 d7 d4 cc d0 ca cf d8 c5 ce c9 c5 c4 c8 c5 c1 c1 c0 c3 b4 bd bf b6 b7 bb b7 b9 b7 ad ae a6 a8 a3 a1 9a 92 9c 94 8a 8a 89 88 8d 85 8a 7d 76 80 73 7b 74 74 67 68 66 69 7d a3 a0 86 58 2e 22 0d 08 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 0a 17 23 38 41 53 68 74 78 7b 77 73 61 60 5b 61 5d 5c 57 64 63 69 67 6f 6f 70 6a 73 71 77 76 73 79 81 7e 85 88 90 89
 90 95 98 99 a1 a6 a0 a8 ac b0 ae b4 b6 b8 b8 b3 b7 af b7 bc b8 be bc c4 c5 c9 d0 d7 d7 dc de dc e6 e8 e3 e8 e5 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff de ce ca c4 c4 c1 c2 b8 c3 bd be ba b9 be bf be c4 c5 c9 c7 c8 d3 d5 d5 e2 df e4 df e0 d8 e0 d9 d7 dd da db d5 d3 d3 cd c6 d2 d0 d0 c8 cd c9 c9 c5 c3 c3 c1 c1 c2 bd be bb b8 b6 b3 b5 b4 ab ae b2 a3 a6 9e a1 90 98 97 8d 8e 8e 8d 88 81 85 75 7c 7a 79 75 78 72 69 72 6c 72 7b 9d 9e 86 5b 3a 27 24 1a 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 08 12 17 23 27 36 40 5a 68 78 75 83 77 71 63 57 54 57 5b 57 58 5c 61 62 6a 61 69 6c 79 6f 75 76 7f 80 7e 81 83 8a 8d 8f 91 93 9d 9a 9f a4 a4 a9 aa ab b2 ae aa b9 ba bb b4 ae b7 ba be c1 bf c1 c5 d2 cd d3 d6 d3 d9 d5 e1 e9 e6 ea eb f3 fa fe fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee d9 cf c2 c5 c6 c3 b4 c3 bd b8 c1 b5 bc be bc bc bd c1 c5 ce cf cf d2 d7 d4 da e1 d4 dc dd d6 dc dc d1 d0 d3 d5 d0 d6 cd ca c4 cc d2 ce cb c1 c8 cb c4 c6 c2 c7 c6 bf c0 b8 b2 b3 b5 af ae af a5 9d a1 9a 9e 9d 98 95 8a 8d 90 95 93 89 83 7d 88 80 79 7e 76 77 74 78 70 73 7c 9d a2 84 60 37 24 24 1c 0e 0b 07 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 11 21 35 30 4b 5e 77 80 7b 6d 6a 67 59 55 4c 55 51 57 5d 54 5a 60 63 63 71 6d 64 76 75 75 7c 76 83 83 8b 8d 86 90 91 9e 94 a4 a4 aa a5 a5 a5 b1 b1 b0 b7 b5 b9 ba bf be bb c2 bc c3 c6 c6 c5 c5 c8 d2 d4 d4 de d9 e0 e0 df e9 f1 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 d0 cf cc c5 c9 c0 ba bc b6 be be b7 b7 b5 b4 bc bb be c1 c5 ce d0 cf d5 d7 d8 d1 d4 da d8 d6 d7 d9 db d5 d4 d4 d4 d2 d0 cb cc cd cb cb ca c3 c5 bc c9 c3 c0 c0 b7 bc b5 ae af a7 ad a9 a5 a5 a5 a0 99 9f a1 94 9a 95 8e 88 8b 94 86 7c 84 84 80 7a 7b 78 7b 7b 7b 76 72 67 73 97 9e 8c 6b 39 32 25 2c 1a 10 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0e 1c 2a 36 42 4d 67 75 7d 71 6a 61 61 58 4b 54 56 5e 5a 57 5e 5b 60 62 65 62 6d 62 65 6c 76 7a 79 7f 7e 86 83 8c 8f 90
 9d a0 9c a4 ab ac a8 ad b0 b8 b6 b7 c0 b8 c3 bc c4 ba c7 ce cb c7 ce ce c7 cc d2 d8 ca d1 d5 d9 e1 e9 f2 f9 f8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d7 d4 c9 cf bb c0 ae ba b7 b5 be ba b9 b8 b6 b8 b4 bf c3 c7 c8 c6 c4 d1 d1 d4 d0 da dd d9 de d6 dc db d2 d3 cf d8 d0 d3 d0 cd cd d2 d5 c9 c9 c7 bf c6 cb c0 c2 b4 b6 ae b0 ac ad b0 ac a5 a0 a5 96 92 99 9c 9e 9e 94 8b 88 90 8b 84 8d 89 86 89 80 80 7d 76 7e 80 70 6e 72 67 84 9e 95 79 58 40 40 33 24 11 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0a 15 14 2c 37 46 50 6a 7d 80 6a 66 65 62 55 53 59 58 5e 55 58 58 60 62 63 62 64 62 67 67 6a 77 74 7a 7b 80 82 87 8f 8d 94 97 9e 96 9b a2 a7 ab ae af b5 bc b9 bc c4 b5 c6 c3 bc c7 cc c7 cf cb ce c9 ce d6 d3 d8 d2 dd de dc e2 eb f5 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 d3 cc c2 c8 c7 be b7 bb b1 b7 bb b5 b8 bf b6 c0 c0 bc c3 c6 c4 ca d0 ce cb d3 d3 d7 d5 dc d9 dc de d8 d4 d7 d6 d9 cc cf ce d6 cc ce bf c3 c7 c3 c3 bd bb bb b4 ac b2 b4 aa ae ab a3 a6 9a 9d 96 9f 9a 96 99 96 98 9b 90 90 95 89 87 8f 85 8d 80 81 88 7e 7f 71 72 77 6b 70 74 8b 99 83 66 5c 4c 3e 22 19 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 1f 25 3d 4a 5c 68 7f 7f 69 65 5e 59 56 54 5b 57 57 54 56 5a 60 64 61 62 63 61 69 6d 72 71 75 78 79 7c 87 8d 85 81 90 95 95 98 98 9b a7 a2 b0 b2 ab b6 b2 b3 b9 ba bd c4 be ca c4 c7 c8 ca c6 cc d5 d4 d6 d4 d7 df df e8 ed f5 f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ab ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed cf c9 be c0 bd b7 c0 b2 ba b1 bb b5 ba b2 be b6 b5 b4 b4 c3 c2 c1 c6 ca cd d2 c9 d0 cf d3 d2 db dc db d4 d4 cf d1 d3 c9 cf c7 ca d3 c4 c8 c3 c4 c3 bb c2 b5 b5 b0 b1 a9 ad 9e ac 9d a3 9a 95 95 99 9a 96 98 9a 99 99 97 92 8d 8c 8c 92 86 8a 81 84 79 82 78 79 6f 74 6f 6b 67 79 93 8e 76 6b 50 37 29 1f 0f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 13 1f 31 3a 4b 63 76 7e 7e 68 60 58 4f 5e 54 5d 67 59 60 61 56 60 55 64 6b 60 73 69 60 6f 74 79 7a 7b 82 84 86 8b 8b 90
 94 95 95 94 a9 9f a4 ab a8 b4 b5 b3 bf c1 be c9 c5 c5 ca c7 cb d1 cc c7 d4 d0 d2 db d7 da e6 eb ef f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f0 cb ea e4 dc de de e5 e9 f2 ff ff ff ff ff ff ff ff ff ff dc c8 c4 c7 c2 c9 b9 b6 b1 b9 b9 b3 b2 b9 bd b3 b0 b0 bb bd bf c6 c7 c0 c8 d2 d0 d2 da db d4 da d8 db d4 d9 cf d5 cc d3 d0 d0 d5 d9 c6 d0 c6 bf c2 c9 c5 bc bb b9 b4 ac aa af b2 9f a4 a3 a2 9c a1 a0 96 9b 9c 9d 98 96 9d 90 94 8b 8d 82 87 85 7e 7c 76 74 71 73 76 67 67 75 6d 89 92 8b 76 59 4f 38 23 18 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0e 19 18 2b 35 4b 61 6f 87 83 61 5b 57 57 58 5d 5d 5e 5b 56 60 5e 6c 61 6d 64 6c 70 64 6b 6f 77 74 74 7b 7f 84 82 8c 84 9b 9b 99 94 96 9f 9c a5 9d ad ae b4 ae be bd c1 c6 ca c9 cd cb d2 d5 d6 d3 d7 db d9 e3 e2 e1 df ee f3 f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ec de db d8 c9 cd cb c7 c9 ca c9 d1 df ef f5 ff ff ff ff ff ff ff ef c8 cc c2 c2 ba bb b5 be b5 b7 b9 b2 b5 b2 af b7 ba b9 b9 c2 c1 cb c6 c0 cb d1 d1 d6 db d3 d3 d1 d7 d4 ce d1 d2 d3 d6 d9 d2 ce db ca ce d0 c5 c2 c7 c2 c3 c3 af b0 b2 a8 ad a5 af a5 9f a3 a2 9d 9e a8 a1 94 9e 9a 99 9c 93 87 8d 91 8f 8d 82 85 7c 79 75 75 6e 71 6e 6a 67 6e 78 96 90 84 65 42 33 2b 14 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 1e 2c 43 48 63 76 7d 7a 67 53 50 54 5c 58 54 5c 61 5d 63 5f 68 62 63 6c 61 6a 65 6b 77 6f 79 76 74 7d 7b 8a 84 89 95 95 94 9e a5 a7 a1 a5 a7 aa a3 b1 b5 b7 bd bd c9 c7 c2 c3 c9 d2 d6 d3 d0 d5 de e4 d9 e3 e4 e5 ed f6 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e8 db db c9 c2 b5 b8 af b6 a8 ab b2 b6 b3 be c6 d0 d9 e6 f7 ff ff ff ff ff d6 c7 c9 be b6 b2 bb b5 b3 b8 b9 b1 b6 ba b5 b9 b1 b2 b8 bf c1 c1 c4 be c2 cd ce cf cf cd d3 d3 d3 d0 d1 d4 d2 d9 d3 ce d9 d5 ce cd ca d4 bd cb c3 bd b9 b8 b9 b5 b0 b2 ad ad ab a4 ad a4 9e 9b 9f 9e aa 9b 9a 9c 92 98 94 94 8f 90 8b 82 86 82 80 78 7c 6e 6d 71 6d 6e 67 75 75 84 90 8a 67 50 35 21 14 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 1c 22 2c 3b 4e 66 76 7f 7e 64 58 54 4d 5a 5c 58 64 58 64 61 5e 66 6a 60 62 67 70 71 6c 6f 69 79 76 76 75 70 84 81 8d 94
 9b 9c 9a a0 a9 aa aa a2 ab ae ac c3 bd b7 c4 c8 c5 c7 cb ce d3 d3 d2 d8 e3 de e5 e4 e4 e8 f0 f5 f8 fd f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e3 d1 cc bc be ae a1 9e a2 9c 9e 9e 99 a0 9f 9f a8 b1 b1 c1 c5 d6 e7 ff ff ff ff f1 d3 bb c2 b3 b4 b7 b5 b6 b2 b4 b5 af b7 aa b6 bc b9 b9 bc c3 bf c0 c1 be c9 c7 c7 c8 d1 d4 d0 d9 ce d6 d5 d1 ce d9 cf de d1 d4 cd d2 d0 c7 c9 c6 bd b5 b9 b0 b9 b0 af ae b3 b3 ae ab ae a5 a4 9d 9b a2 95 9e 90 8b 94 95 95 87 92 87 8e 86 82 7c 82 75 6f 73 6b 62 66 6f 69 74 70 91 84 73 5c 3b 34 1a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0f 1f 25 33 46 51 6c 7d 7f 72 5c 58 59 52 61 5b 56 5f 5c 5d 64 5f 61 66 65 64 6b 6d 70 74 74 72 79 7a 76 82 84 85 84 8e 83 8e 99 91 93 a5 9f a5 b0 b4 a5 b8 ba bd b7 bf bd c3 c9 c6 d7 d7 d5 dc df dd e7 e5 e3 ed ed f3 f0 f2 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f2 da cb c9 bb aa a9 9d 98 92 92 8c 90 8c 8a 7d 8d 7d 96 96 95 a6 af b6 d2 e3 ff ff ff ff d5 bd bf ad b5 b5 ae ab af b3 bd b9 b8 af b1 b4 b1 b8 b9 b7 bd c4 ba b9 c4 cb d2 cc d0 ce d5 d4 d0 d5 d8 d8 d5 d3 d4 d5 d2 d2 c8 d1 c9 c4 ce c1 c3 c3 b2 ba b0 b2 ad b5 b5 a6 af a7 a9 a4 9e a5 a8 a2 a1 99 9a 8c 93 8f 95 9b 85 89 8b 81 81 7d 7b 76 76 73 7a 63 68 6a 66 66 7e 8a 94 6e 54 46 2c 1d 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 16 1f 27 40 4f 61 7f 89 72 5d 58 4e 56 56 58 56 5f 5e 62 62 65 57 5e 5f 6a 70 69 64 6e 76 75 77 76 77 7a 83 7e 8d 8d 8c 92 90 94 97 a5 a4 a6 ad af a9 ad b7 b9 bf bc bf bd ce c8 ce d4 d5 d4 da dd db e3 ec f0 ed e9 f5 f3 f5 fa fa fb ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 db e1 cd c7 b1 a5 9a 91 84 83 7b 77 75 7a 78 76 76 72 6b 6f 81 7b 90 95 9f ab c6 d6 e7 ff ff e6 c1 bb b1 b5 b2 bb ac a7 b0 a7 b2 b2 ad b8 ad b0 b9 b0 b3 bf ba b6 bb c7 be c6 cf c9 cf ce d5 ca d2 d6 cf d1 cf d7 cd d8 d7 cd d6 cd c3 c9 c4 c5 ba b5 b5 b0 b3 b1 b2 ab ac b1 ad a6 a2 9e 9f 9b 9d 9e 97 9e 93 93 8c 91 8a 8f 89 83 7b 76 75 79 6f 75 69 69 65 67 6f 70 6b 74 8e 93 70 59 4c 26 20 0e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 08 12 1a 2d 38 52 67 77 7a 68 60 61 56 5a 60 5e 5c 55 5e 61 60 60 67 5d 62 6b 6d 6f 6b 66 70 71 7c 7a 80 81 85 86 87 92 8a
 94 90 97 a0 9c a0 a1 a8 a1 ad b1 b9 bc bd c6 be ce ca c4 d7 d5 d4 e0 d9 e2 e5 e5 e3 eb e8 ee f8 f3 f4 fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e0 d5 d4 c9 ad 9e 90 85 7c 74 68 66 50 50 5d 52 58 57 51 59 59 6c 6b 75 81 86 8f a1 b6 c8 e0 ff f0 c5 b5 b5 b0 af ac b4 af b4 ab ab b5 ad b5 b0 b7 b5 be ae c6 bd b7 bb ba c1 c1 bd c2 c4 c6 d8 ca c9 ce cf d3 d6 db d2 da cd cf d1 c9 c4 c2 c6 c0 b8 b4 b9 b4 af b1 ae a7 aa af a3 a8 a4 9f 9d a1 9f 9b 99 96 8a 8f 8d 8a 8e 87 7e 85 81 79 77 77 6d 6f 6c 6e 6d 6a 67 67 6b 6d 89 90 7a 60 41 36 1a 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 14 25 30 40 54 6a 77 7d 69 5b 5a 5b 58 5b 56 62 67 62 60 64 62 66 64 66 65 71 6f 69 67 75 77 7a 79 7e 7b 7d 82 8b 93 95 92 93 97 a3 a7 a1 a2 ab ae ad a9 b3 b8 bf ca c0 cb ce d5 d3 d2 d4 da da dd e6 e0 e4 e5 e9 f1 ef f3 f4 f9 fc fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 d2 c9 bf a8 94 89 7c 59 60 54 49 4f 4d 46 44 48 49 46 4e 4c 4f 50 5f 60 67 6b 71 8d a0 a6 be f5 f4 d0 c0 b1 b7 b0 af b6 ab af b1 a9 b0 ba b2 bc b3 b7 bc b0 bc bc b5 b6 bb bb c1 c7 bf cb c2 ce c9 cc cf d0 d7 d6 ce d9 d3 d5 ce c4 c9 c0 c3 be c3 b1 b6 b9 ae a9 ae a7 ab a3 a0 9d 9d a7 9e a3 97 96 96 94 8f 8f 8e 89 8c 8d 8e 82 86 7d 7f 78 76 6f 6e 6e 67 63 6c 6e 69 68 74 85 97 7a 68 42 35 28 0b 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0e 19 2c 42 5a 6f 7b 78 6e 5f 58 5b 58 5e 5b 63 64 69 64 5e 63 65 6b 65 68 71 6f 73 72 6c 71 7e 75 7d 85 87 88 86 85 8a 9b 90 9b 9b a7 99 a8 a7 aa b6 b7 b7 ba b8 bc cb ca cf d3 d0 d6 d5 d9 d8 e5 e3 dc e8 e6 e6 ed f1 f3 f5 f4 fc fc ff ff fa ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 c9 b5 a8 96 7c 73 60 54 46 4c 46 45 3e 3e 44 40 41 42 41 3c 3f 50 50 4a 4d 5a 62 6d 81 8e 9d ce f7 e1 c9 b6 ad af b2 b1 af b5 b6 aa b0 bd b7 ae b2 b1 bc bb bd b8 ba b6 be b8 c2 bc c4 c8 ca cc ce cc cc cb cf d0 d7 d3 d0 d1 ca c7 c5 ba be b9 b6 b0 ad ae b0 a9 af a3 ad a2 9f a5 a5 9c 9c 9b 98 93 95 95 98 93 90 8c 88 89 89 88 84 7a 7d 75 74 73 69 6d 6d 69 65 5a 60 6a 72 8a 92 73 62 3e 3a 1b 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0b 19 1d 2a 42 51 66 7a 78 62 5e 5b 59 61 65 67 68 64 66 6c 6c 6c 67 6c 6c 69 6c 6c 6d 79 75 82 80 83 80 8b 88 84 8f 90 8b
 8f 93 98 9c 97 a8 9e a6 ac af ad b6 b2 ba bd c1 c1 c4 cc d2 dc d9 d4 d5 dc df da e4 e3 e0 e2 ee f1 f0 ef f2 f9 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee bd a6 95 73 64 55 43 41 3d 45 3e 42 3e 3b 3b 41 37 43 3d 3e 36 41 43 43 44 4b 4d 54 69 72 8e b3 e1 e2 bd b5 b7 ad b0 b2 b5 b0 ac b5 b1 b1 b7 b7 b2 ba bb ac ba be b7 b9 bd b8 c2 bd c3 c1 c6 d1 d6 d0 d1 ca cd d3 ce cf c7 cd c9 c1 c3 ba b2 b2 b0 b0 a8 aa a5 a4 9f a3 a0 9f a0 a6 9f 9a 95 9e 91 95 8b 88 8c 87 8f 86 87 84 8a 86 82 71 73 72 72 74 6f 70 6c 68 68 6a 64 6a 71 89 89 7c 61 4c 36 1d 08 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 14 1a 2f 38 59 61 70 7c 67 5f 59 53 5a 62 69 6a 6b 66 67 6a 74 6f 6b 6d 6d 72 74 77 71 78 7b 84 84 83 8a 89 8b 8f 91 8f 8f 8f 9d 93 a4 9b a0 a6 af a9 af b0 b6 b0 b2 c0 c1 c9 c7 cd cd d6 dc e4 d8 d9 d9 e3 e4 e6 e3 eb ee e7 f6 fc ff ff f2 ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d5 ab 92 75 5d 45 44 51 47 3b 3f 36 36 42 37 31 3e 36 2e 31 3c 3a 38 3b 41 42 3c 43 50 57 67 79 94 cd e4 c1 c0 b0 ac b6 b3 b6 b3 ba b0 b7 b3 b2 b4 b1 b8 b7 b6 bd b8 b5 bd b9 b9 c5 b8 c5 c9 d4 d1 d0 d3 cf c7 d0 c6 cf cd c1 cc bd b6 bc b5 b0 ad ae a7 a7 a9 9c a6 9b 98 9e 9e 9c 9e 91 98 93 99 8e 94 8e 93 90 8e 8c 8d 84 82 86 78 80 79 7b 70 64 73 6f 73 6d 69 67 63 63 71 6e 84 95 7e 5f 51 3b 1e 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 15 15 26 3c 4b 5d 70 78 60 63 62 5d 61 5f 66 64 69 70 69 69 6e 75 71 6d 6d 69 6d 78 76 79 83 80 83 7f 86 8c 83 89 93 94 97 93 9a a1 a4 9f a9 a4 a7 b1 a5 a9 b3 b5 b8 bd c4 ca ca cc cb d3 d6 e0 e0 dd db e0 e6 e2 e8 ed f6 ed f0 f7 f9 fe f6 f7 fa ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 b5 8f 74 5f 53 41 40 3d 36 41 35 2e 36 30 27 25 28 2b 28 30 26 29 2c 35 37 3f 3f 44 45 4d 4e 6f 87 be e3 cf b4 b6 ac b4 b6 b1 b2 af af b7 b2 b4 b3 b4 ba b7 b8 b4 b5 c3 b9 bb bb c0 ba bf c4 ca c7 cc c7 ce cf cc c7 bf bb c1 c6 af b6 b2 aa a9 ac a6 a2 a7 9c a2 9e 9a 99 98 a0 96 9e 96 8e 8a 86 8a 8d 86 89 8a 83 8b 81 81 86 81 7f 80 6d 7c 7d 71 72 6c 6b 67 67 6a 65 6c 65 81 8a 93 82 6c 4a 30 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 11 1e 24 38 49 67 75 74 65 56 5d 56 5c 65 66 6a 6a 6b 6f 72 6e 69 74 77 6c 73 77 70 7d 74 83 80 7c 83 81 89 8b 8c 89 95
 90 91 9a 97 9f a2 9d a4 a6 a1 a7 ac ae b3 b4 b9 b9 b9 c9 c5 c7 d0 d1 d1 d6 dd d5 cf dd e0 dc e3 e8 e6 f0 ec ef f4 f7 f5 fa f8 fe ff fc f9 fd ff f9 fc fe fd ff ff fe f5 ff fa ff fa ff ff ff ff ff ff ff ff f4 c0 93 7a 5c 4b 42 35 34 39 28 33 25 2d 27 28 28 27 1b 20 15 1f 20 28 29 2d 31 38 34 37 37 47 43 5f 7f a9 da d2 c1 bb b6 b1 b1 ae b6 b1 b6 b4 b7 b1 b6 be b7 b8 ac b2 b2 b2 be b8 b7 be ba ba bd c6 be c8 c1 c6 c5 c5 c6 c1 be b0 ba ac ac ae a0 a7 a4 9b a1 9c 95 9d 97 99 96 94 9a 8c 8e 91 8f 8a 8b 8d 8c 85 83 82 80 85 8b 80 86 82 7a 76 7c 74 71 6b 6e 65 62 65 63 5a 62 6c 70 76 8b 95 83 66 44 2b 16 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 15 14 25 3b 4b 61 74 75 65 5c 5d 5e 57 5e 64 6b 68 70 6d 6a 74 73 72 77 79 7b 79 7e 7e 7f 85 79 80 82 88 89 8c 87 8f 8d 93 98 93 9a 9f 9b a0 a0 a2 a3 a8 a8 ae ac af ba bb b9 c3 c5 c3 ce d1 cc d4 ca d5 cd d9 db dc df e8 e4 ea ef e7 ef f3 f2 fd f3 f7 f7 f5 f7 f2 f8 f7 f0 ef f4 f6 fd f7 f9 fc f0 f8 fd f9 f7 fe ff ff ff ff ff e2 a4 7e 64 4d 42 3f 31 31 2c 2c 2f 25 24 1a 17 1e 1d 1b 23 1a 1f 22 24 22 23 26 2c 2d 2f 35 3f 4f 51 72 a0 d3 d3 c4 c7 b6 b3 ba b4 b0 b6 b9 b8 b8 be bb b6 b4 bd b4 b3 b2 b9 be b4 b2 c1 b9 bf c0 c4 cc c7 bf c1 c5 c1 b7 b7 b5 af a9 ae a9 a8 a1 a0 97 96 a1 9e 94 9c 94 91 90 8d 93 8c 8e 8e 8c 89 8e 81 8a 85 89 8b 84 8b 7e 80 7a 7f 7d 7a 7a 77 72 6e 6a 6a 63 64 64 5f 61 69 6f 78 85 95 7f 66 4d 3a 15 12 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0e 1c 28 35 4a 67 6f 81 61 59 63 5c 5c 62 66 63 6f 6f 69 6f 6f 71 70 73 76 77 80 79 7c 80 79 7e 84 85 86 8f 85 89 89 8b 94 97 93 98 97 9e 9c 96 9a a3 9f a5 a9 b0 af b9 b4 af bd bf bc bc c2 c4 cf cf ca d0 d4 d4 da d9 dd e7 e2 e9 de e9 f1 e6 f1 f5 f6 f6 f5 f1 fb f6 f4 ef f6 f2 f0 f0 f9 f5 f6 f8 f6 f8 f7 f8 f8 ff ff ff ff ff cc 97 76 5a 46 36 2d 28 22 24 20 25 24 1f 14 15 17 1a 19 15 16 17 17 15 1f 20 1e 25 22 2a 35 36 44 51 68 9a d1 cc c5 c5 ba b1 be af b3 b7 b1 bc bb c2 c4 bf b8 b0 b5 b6 ae b0 ae b6 ae b7 b6 b5 bd bc c2 c6 c0 c2 c0 bf b9 b3 ad ab af a5 a1 a1 9b 9c 9e 92 9b 90 8f 92 8f 8c 8e 8c 8f 88 8b 94 84 81 85 88 89 80 81 84 84 85 87 81 7d 7a 79 76 74 71 76 75 65 69 6a 67 6a 6b 5d 65 70 72 84 96 81 65 44 28 1c 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 08 1a 23 39 54 62 78 70 69 5d 53 55 5c 64 5d 65 68 69 6b 68 73 71 7a 75 71 7a 7d 7a 83 7d 7c 84 86 80 85 88 89 8b 8b 8d
 97 8f 96 8f 8e 98 94 9e a0 9f a5 a5 af a8 af b5 b0 b1 b6 b7 b7 bf be c5 c1 c7 cd cb c7 d7 d6 d6 d5 dc df de e2 e1 e7 e6 ee e3 e6 ec e8 ec ea ef e8 ed f2 ef f0 ee f3 e4 f2 f3 e8 f4 ed f4 fc fd ff ff ff fe b2 83 6a 52 41 32 25 23 26 20 1a 19 1c 1a 16 15 11 14 13 1a 05 10 14 0e 16 19 10 15 1e 1f 25 2f 35 52 64 8c c7 cf ca c0 b7 b4 bd be b9 b5 b9 b5 bb b9 b7 b9 bd b2 ae b4 af ae b0 b4 b5 b2 b7 b6 bb bc bd b9 bb b4 b8 b8 b1 a9 ae aa a3 9d 9c 96 8f 93 90 8b 99 90 86 8d 8a 89 85 89 8d 85 86 84 7f 83 7d 81 88 86 84 83 77 7d 82 7a 7f 78 78 7b 6f 77 67 6b 6c 6c 69 5b 69 68 65 5f 6c 70 82 8b 78 60 46 34 22 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0c 15 30 3d 50 65 76 74 6b 61 5a 5e 62 63 62 66 69 6a 72 69 73 76 71 77 73 74 79 75 7c 7f 7c 7f 86 80 85 8e 83 90 93 8e 91 8f 92 93 92 95 99 9c 9e 9a a3 a6 a2 a7 a3 ac b8 ac b5 b2 b4 bb c0 bd c1 bf c2 c9 d2 d0 cd cc d6 dd d4 de d8 d8 dd d9 e2 e0 dc e9 e2 e7 e6 e3 e8 ef ee f0 e2 e5 e6 e9 e3 e8 ed e8 f1 ef e5 f0 ff ff ff ea ab 81 63 47 37 32 2b 1f 20 13 19 13 0c 0d 0e 0e 03 12 0c 0d 13 0c 0c 13 13 1f 20 1b 16 1b 1a 23 33 52 6f 8b c8 ce cd c5 bc c6 bb bd ba be ba c5 c1 c5 c3 bc bc b4 ae ab aa b7 af b2 ae b0 ab ba bf b9 b9 b9 b1 b1 b3 aa b0 a0 96 a5 a2 95 9e 92 92 89 91 94 87 8d 87 82 85 87 86 84 89 77 81 84 7a 82 82 7c 83 7b 83 81 7b 7f 7c 7b 7a 75 73 75 6f 6b 71 68 6e 64 61 6e 62 65 65 6b 70 6a 85 8c 78 64 4b 2f 24 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 16 2c 38 50 64 74 79 65 60 60 5b 61 61 65 65 6f 70 71 69 72 74 74 73 76 79 7a 81 7f 83 77 7b 77 7c 82 88 8b 8a 8a 8d 94 8f 8f 90 92 90 92 96 9b 9d 9c a2 a2 ab a7 a4 a7 a4 ad b0 b0 b1 b7 b7 b3 ba c4 b7 c1 ca c0 d3 d4 d1 d1 da d6 da da d9 e1 de e4 e3 db e0 de e9 e1 db e5 e0 e7 e9 e5 db e5 e1 e6 e4 ea e7 e9 e8 fe ff ff da 93 77 59 48 36 2a 1e 0d 16 0e 14 0f 09 0d 0a 13 0e 0b 0a 10 05 12 10 15 0c 13 15 18 16 1d 21 2c 2b 48 68 8e c8 d1 d2 d1 c5 be c3 b9 bb c7 c3 c1 c1 c1 c5 b7 b6 ae aa b1 ae b6 be bb a6 b4 a7 a4 ad b0 af b5 b2 b5 ad ac a5 a2 a0 98 9d 93 90 8f 8e 8b 8e 89 88 88 85 86 83 7e 85 7e 84 87 83 8e 7f 7a 7e 84 7c 86 81 7f 7b 82 7b 7f 73 77 72 75 6c 6e 6f 60 66 6b 62 68 70 65 66 67 69 6a 7d 88 76 64 46 2e 13 0e 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 11 14 25 37 4e 66 6f 76 67 5c 62 58 5f 5e 60 6b 70 70 6f 72 6b 72 77 75 79 7f 78 7c 7b 80 80 7c 7b 81 83 81 7f 7d 86 7d
 8e 8a 87 8c 8f 90 94 92 92 9a 96 93 99 9e 9d a0 aa a7 a5 a5 b1 aa b3 b3 bc bd b3 ba b9 b9 be c0 c0 c2 ca d8 d4 d2 d7 d4 d3 d7 d6 e5 dc d3 dd e0 dd e1 e6 dc da e0 e1 db dc e1 df e4 dc e3 e6 e6 ed ff ff e5 a2 6e 55 44 37 1f 17 0f 17 16 0b 0d 07 0a 06 08 07 0d 08 0b 06 0b 0a 0e 11 04 0a 0a 12 1c 22 1b 2b 3c 6b 95 c5 cc d5 cb c5 bf c2 c5 c3 bf bc bb c0 b6 bf b0 ab b0 a8 a3 ac b3 b5 b1 ac ab aa a4 a5 ab a8 ae ae aa a3 a3 9c 9b a0 94 95 8b 89 8a 89 86 8b 80 81 83 82 84 80 7d 82 7f 7a 81 77 78 79 79 80 6d 77 75 80 7d 77 7a 77 70 72 76 77 72 6f 66 6c 68 68 6b 6b 65 5f 60 67 61 69 69 78 84 6d 57 44 1f 17 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 0b 20 22 37 4a 67 76 7d 69 5a 5a 62 62 68 67 66 6a 71 75 75 6f 79 76 77 6f 7c 75 79 72 7a 7a 7b 7b 7d 7f 80 7e 84 91 8a 8a 85 84 84 8d 8a 88 8b 8e 8d 8e 9c 96 97 9c a3 a6 a8 9c aa 9d a8 b1 ac b5 b3 ac b1 bc b9 bb bc c7 c2 ca ca cf ce d3 d1 d0 d0 d6 d3 db de d4 db d4 d1 db d6 d7 dc e1 dc dc dc da db d9 df e5 e2 de ff ff fb ac 69 56 47 27 13 0d 17 0e 08 08 0d 11 0b 06 08 08 05 06 05 0a 09 10 05 04 0c 0f 0d 12 0e 16 1e 24 3c 69 9c c9 d6 d2 d3 c9 c3 d0 c3 c8 c4 c7 c2 bc be b4 b5 b1 aa aa a3 a9 b9 b3 aa a0 af a6 a7 9e a0 a0 a0 a8 a9 a1 a6 9a 93 8c 89 90 84 84 82 84 80 7e 7a 84 7d 7e 84 7f 8a 7c 84 7d 79 7c 75 78 7a 7b 7c 81 70 77 76 72 75 71 74 77 73 70 71 76 6e 65 6c 64 68 68 68 5e 69 66 70 66 69 6b 7f 69 5e 40 26 18 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 10 12 2b 35 4b 66 79 79 63 62 5f 5a 5f 68 64 6c 6d 72 73 6b 6d 72 70 79 7c 78 7d 7d 7a 7a 84 7f 7a 7b 83 80 77 86 82 80 7e 82 87 84 89 89 8e 94 90 8d 95 94 94 96 9a 99 9c a4 a5 a5 a5 a8 b0 a7 ad a6 b1 b2 b7 b4 b5 bf b7 c4 c1 c5 cc c4 c4 ca d6 d0 d3 d9 d8 d6 d3 d1 da d3 d3 db dc db d6 d5 df d5 d6 d4 d2 d9 de db e5 f5 ff ff ba 73 55 47 22 1b 06 08 0b 0d 0f 0d 07 0c 0d 0e 0a 0d 07 06 0c 08 08 09 05 02 0a 17 17 0f 16 19 23 33 72 ac c9 d8 d5 cd cb cb cd c7 c5 ca c7 c0 bf bc b5 af a9 a9 a4 a8 ac b3 ae aa aa a5 a3 9a a2 99 9d a5 9f a4 9a 99 9d 90 85 8e 8d 84 80 87 7f 7d 77 75 76 7c 7e 7b 7d 7e 7f 7b 75 7c 81 7d 71 7f 76 75 77 7d 7b 77 7d 72 73 75 75 6f 75 6e 65 6d 6e 66 65 66 70 69 6b 6a 6e 69 68 6a 6f 7d 6f 5a 42 29 22 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 16 1b 21 37 4a 69 71 77 6f 63 5e 5a 63 60 65 5f 67 6f 70 69 73 6f 74 79 76 73 7b 79 6f 70 80 79 79 7b 7b 80 80 7b 84 82
 89 81 81 85 86 87 81 88 8a 92 93 9b 92 99 93 99 9e 99 98 a1 a5 9f a5 a9 a8 a0 a9 b2 af b1 ba b0 b7 b6 b7 c5 c5 be bf c6 c3 c7 ce c9 c9 cb cd cd cc d2 cc d0 d3 d8 d5 d3 d3 cf d6 dc d7 d6 d1 d2 d2 e7 ff ff d6 82 54 43 24 0f 08 05 03 0b 06 05 03 08 06 0a 08 00 06 09 06 07 09 05 0b 0b 0e 0f 0b 0a 0f 1a 1f 32 76 b0 c9 cf d5 d3 c8 d6 d1 cd c6 c5 c0 c5 c2 bf b3 ae a8 9f 9f ad aa b0 ac 9d a8 a6 a6 95 99 a2 95 a1 8f 95 96 94 8d 90 86 87 87 7e 81 7c 80 80 76 7a 7d 7b 7d 77 77 7d 7a 78 73 70 77 72 6e 71 78 7b 70 76 75 73 78 6e 75 6c 70 67 6f 73 69 6e 64 68 69 6f 66 6d 68 6b 68 64 67 66 62 78 6d 5a 40 26 14 03 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 12 10 2a 3b 47 65 6d 73 6d 5d 5f 63 62 69 6a 68 6f 6b 6b 74 70 6e 73 73 79 7a 77 7b 7c 76 7c 78 7b 7a 7c 8a 77 7d 83 7b 83 7e 81 83 88 83 8d 92 91 8b 96 8f 96 8f 95 9b 97 96 97 9e a2 a0 9e 98 a7 a6 9d a7 a4 a9 a7 b3 b5 b3 b5 bb be b8 b8 c5 c6 c2 c7 cb c5 ca ca c7 c9 cd c6 d1 cd cd d4 d1 d5 cc d9 d6 d2 d0 d5 cc d7 da ed ff e5 a8 64 45 23 13 07 05 03 0e 06 06 05 00 06 06 05 05 06 05 03 01 06 05 03 06 09 05 13 10 0e 0f 19 2e 70 b5 cb ce d5 d5 cc d1 d4 d0 d0 cb c6 bc c4 be b1 b4 a6 ac a0 a8 a8 ad a7 a6 a6 9c 98 9b 97 9b 95 9f 98 92 96 92 84 86 87 89 85 7b 85 71 78 7b 73 77 73 7c 77 7b 7c 7d 7a 72 75 6c 74 75 79 78 7d 77 6d 82 6e 7b 6b 73 77 74 79 6c 6e 6d 6d 6c 69 64 69 60 6a 70 6b 6b 6e 6e 5f 5f 61 68 68 5a 3a 25 15 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 06 0c 1d 25 34 4d 5f 71 79 6e 62 64 61 62 64 69 61 6c 6f 6e 6f 6f 6f 71 75 70 74 75 79 76 6f 76 75 79 78 76 84 79 76 7d 7e 7e 7e 89 89 80 86 85 92 9b 8d 8f 8e 8b 89 93 96 9b 95 96 9b 9a 94 9a a0 9c a1 a2 a2 a6 a8 a9 ac b2 b0 b3 ba bd b5 bf be c3 c4 ca bc c6 c1 c3 c7 c6 c7 c7 c8 c7 d2 d5 d2 d2 cc d0 d0 cf d1 cb cf d7 d4 de fc ee aa 71 45 21 15 0e 08 06 00 06 05 09 09 06 05 07 06 06 0b 05 03 06 08 06 0d 0e 17 0e 0f 07 14 12 2e 78 ba c9 d4 ce d2 cc d0 dc d2 cc ce c8 d2 be b9 b6 a8 a6 a4 a8 aa b1 b0 a9 a2 9f 9c 99 a0 9a 90 90 92 92 8a 87 8a 7c 7e 80 7a 86 77 75 7b 7b 73 73 7b 77 75 7a 78 74 7d 7c 78 77 70 7b 73 73 75 6f 75 77 74 7c 80 6f 7f 71 71 74 78 76 6f 65 6e 6d 6d 71 69 6f 75 75 6c 6a 6b 6c 61 61 6b 62 5f 3c 26 1a 09 0e 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0f 1a 20 40 4e 5f 73 75 68 62 64 63 64 67 67 69 6e 6d 69 6c 70 76 72 74 77 70 70 74 72 78 78 74 74 7e 78 7d 74 7a 7a 81
 7e 7a 80 82 80 8a 8d 85 8f 8e 8e 8b 8f 8c 88 8b 89 87 96 97 94 90 90 92 9a 9b a3 9b a3 a3 95 a5 ac ad a5 b2 ab b0 b3 bb c6 bc c0 ba c1 b5 c4 c6 c6 c8 ca c4 c9 c6 c9 d1 cc cb c6 c8 cb cf ce ca cf cc c6 e2 ea c2 81 48 20 0e 06 05 04 04 06 05 03 0b 08 05 07 00 06 05 03 06 06 05 03 09 06 14 0d 07 08 0e 1b 24 74 b5 c7 ce d5 ce ca d8 d2 d3 ce da cf c6 c9 be b1 ac a8 9e 9e a4 a8 ab a2 a7 9f 9c 94 96 93 93 8b 94 8e 8d 87 84 80 81 80 7f 77 7c 80 78 6e 76 75 78 7c 77 74 81 6f 7b 75 7a 84 78 74 73 72 76 75 70 77 76 78 77 77 72 75 6f 70 6e 75 69 70 69 6c 6b 74 70 72 7b 72 6a 68 60 62 61 64 69 64 56 3e 26 0d 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0f 18 22 37 46 58 76 78 6c 6a 62 64 64 64 63 63 6d 6d 66 6c 6e 6d 71 73 74 6f 77 72 6b 75 75 75 73 6f 6e 73 7c 6f 78 7d 7a 79 81 81 7f 83 8b 81 85 82 8d 8b 81 8c 8c 8a 8a 8a 8d 92 91 8d 91 93 98 89 95 98 9b 95 9a a4 9d a2 a3 b0 af af ae b6 b5 ac b2 b1 c3 b7 bb b9 c7 c0 c1 c3 bb c1 c5 c5 c5 c7 c7 ce c7 d1 cd c6 c4 c4 c8 c5 d1 bb 87 44 1b 07 09 05 03 00 06 05 03 02 06 05 03 00 06 05 03 02 06 05 06 00 06 07 0d 08 08 0b 18 34 74 b8 cd d4 d7 d7 cf d3 d5 de da dd d4 c7 bd b2 b8 a9 a5 a5 a0 a4 b0 a3 a5 9a 94 95 96 98 93 8f 8c 85 87 8e 83 85 7d 7e 7a 80 7b 74 77 7c 72 72 77 77 6f 71 7b 76 7a 75 77 7a 7c 74 7e 7e 75 74 76 73 73 71 73 6b 73 75 6e 6f 6c 71 6c 71 6f 6a 62 6a 70 6e 75 6f 62 63 61 6b 62 51 5d 5e 63 54 30 20 17 01 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 09 06 18 2b 30 4a 5b 6e 7f 6c 67 61 67 67 67 63 67 60 70 6f 70 73 74 72 73 75 73 73 77 79 74 75 75 7b 75 70 72 77 77 80 85 81 80 7a 84 87 83 7b 86 80 87 87 89 85 87 84 89 8e 90 81 87 89 8f 8d 8c 92 91 8e 91 92 8e 98 9f 9c a1 a5 b0 a8 a2 ad b1 ba b3 b3 ac ba c1 b9 be c2 ba bf be be ba bf c9 bb c5 c4 bf c3 cb c6 c5 cc ca c7 c4 bf b7 92 4d 25 04 06 05 03 00 06 0a 05 00 07 05 04 03 06 05 03 02 06 05 03 00 06 0c 10 0f 15 0a 15 24 6d b5 cc d5 db d6 d2 db d6 dc d4 d3 d9 cb b7 b4 ac ac a6 a3 9e ac 99 a0 a4 a4 99 91 96 8a 8b 90 8a 8d 85 88 7e 82 80 71 79 75 73 79 7c 76 7e 6f 6f 77 7d 78 79 7c 75 78 76 75 7f 79 7b 72 7a 78 80 81 73 78 70 76 6e 74 74 75 72 72 5f 6f 67 67 71 6e 6e 75 72 70 6a 61 60 63 5d 59 5c 65 61 54 35 22 1a 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 0e 12 21 36 4d 66 70 7d 73 6d 6b 64 62 6a 64 6e 71 6d 70 73 71 76 72 78 7b 75 7a 73 77 76 6f 78 7a 71 78 81 79 7b 7c 82
 7f 82 85 82 85 7f 7d 80 86 8a 87 83 82 84 82 83 80 86 84 89 88 87 8c 86 85 91 87 88 8f 8d 90 94 9a a0 a0 a4 9c a3 a7 a5 b2 ad b3 b5 b2 b2 b6 ae bc af ba c3 ba be c1 be c3 c8 c2 c4 c5 c2 c0 c0 c1 c2 cc bf c0 b8 94 52 22 0d 07 05 07 01 06 0a 03 00 06 05 03 0c 06 05 03 00 06 05 0a 0a 06 0f 0b 0d 0b 0e 13 22 6f b3 ce d6 da d4 da d8 de d8 d9 db cb c9 c5 b5 b9 aa a8 a0 a3 a5 a2 a1 9b a2 8d 94 90 91 93 91 8a 8c 8a 89 80 76 7b 6e 79 7f 7c 74 7c 77 7b 71 7d 70 76 71 76 6f 76 79 6e 7a 73 71 77 73 6e 77 75 77 76 7e 76 71 70 76 74 74 71 77 71 73 69 70 6e 71 75 6f 73 71 6c 6d 63 5e 61 59 58 62 5d 51 3b 34 1a 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 11 15 2e 35 49 51 6c 75 6d 6f 6e 6b 68 60 65 65 72 6d 70 7b 6e 6f 73 70 78 70 6c 74 6f 71 7b 76 76 70 6b 75 71 79 7b 7e 77 75 7a 7c 7c 7c 7d 7a 6e 76 77 80 72 7c 83 7d 80 7e 7b 83 7f 7f 82 84 88 81 8a 88 8a 8f 90 8f a0 90 94 94 97 9a a2 a8 a7 b0 aa ab ad b6 a8 b3 b5 b5 ac b8 b4 be b5 c3 be bb bc c4 bd cf c0 c1 c6 bf bf be b4 ae 96 57 24 09 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 06 0c 0b 14 14 1d 65 b2 cc d2 de de dd d9 dd d9 d6 d6 cf cb bc ba ab a6 a4 a0 a3 a4 9c 9e 9d 98 95 94 8b 92 93 94 94 84 85 80 85 7f 75 6f 75 75 78 7a 7a 7f 71 70 6c 7a 77 6e 6e 65 6d 72 71 74 6f 6d 74 65 6b 66 74 75 74 7c 75 7b 73 67 72 69 6c 72 72 70 74 6f 6e 72 6c 67 75 68 6c 5d 66 60 61 56 58 56 5b 5b 3c 30 17 0e 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 06 12 1b 1f 31 42 5e 6e 83 75 70 72 6f 67 6b 70 73 72 7c 70 73 6d 78 73 7b 70 76 74 74 73 70 72 6e 7a 75 6e 7c 74 7b 7c 78 83 7f 76 7c 79 79 7a 7b 7a 81 77 78 78 79 7d 7a 81 7e 73 80 7c 78 7e 7f 84 82 7d 8b 88 8f 8c 8d 92 8b 93 96 9c 96 9f 9e 9f ab 9d a5 a6 a1 b2 af ac b5 af b5 b2 b5 b5 b8 b6 ba c2 b6 b9 bd ba ba bf bb b5 ba b8 ae 96 66 28 0a 06 05 05 05 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 07 0e 07 13 0f 1f 65 a9 cf d9 de df d9 df de dd dc ce cb bf ba af b2 ad a4 a8 9e 97 aa 9a 9d 9d 99 9a 8b 94 99 91 8f 8b 8b 88 81 82 79 78 79 7b 87 7e 7b 7f 6f 73 76 77 71 74 75 70 6e 6f 72 6a 67 62 66 6a 67 68 6f 71 6f 72 76 75 77 74 75 6b 6d 6a 6c 71 6f 6d 6b 6c 70 6e 6c 71 6d 62 66 60 5a 56 5a 5a 5d 52 3c 2e 1d 14 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0c 1a 24 38 42 61 68 79 7e 68 67 6c 6b 79 72 73 72 73 7f 71 6e 74 7b 75 7d 74 75 7a 70 6f 71 73 79 71 7a 7d 70 7b 83 79
 83 7e 7d 7b 7c 77 7a 78 74 82 72 75 79 80 7b 7e 75 7d 76 7c 79 7d 82 7f 85 7b 7f 84 80 7e 8a 8f 83 8e 8d 94 94 95 93 99 a3 95 a3 a1 a2 a5 a1 a5 ad b1 a9 ab b4 b1 af b7 b4 b2 b8 b2 b8 c1 bd c3 b8 bc bf b7 ac ae 9b 62 33 0e 06 05 03 08 09 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 07 0b 04 08 10 16 24 68 b6 ce d6 de da db df e0 db d0 d8 c7 c5 c0 b7 ac b2 a4 ac a7 a4 a1 a1 9a 9c 98 92 8d 8f 9e 9b 96 8d 8b 86 86 83 7b 81 80 82 83 76 7d 7b 6a 70 74 72 73 74 6d 76 72 70 6f 6d 6e 6a 66 66 62 62 6e 66 6a 6f 77 84 74 6e 6e 6f 70 6f 68 6c 6c 65 66 70 70 6b 6e 65 62 62 60 5e 60 5f 5d 58 61 58 47 2a 25 07 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 11 1a 27 34 49 51 6e 76 7b 63 67 6f 68 73 71 72 7c 75 7c 74 73 71 72 79 77 74 75 6f 71 71 69 6e 69 71 74 71 76 6f 7e 77 7f 7f 83 78 72 75 7c 77 7d 7e 75 78 7c 77 79 78 73 79 76 72 6f 7a 79 80 7b 7a 80 7d 79 7c 87 84 8a 87 85 90 8e 90 92 92 92 9b 96 9b 9a 9f 9f a7 a7 a5 a5 a9 a4 ac b2 b5 b7 a7 b7 b5 b5 b9 b3 b5 b3 b8 b1 ba b0 a7 99 60 33 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 05 06 05 0a 06 0d 0a 0c 1e 5e b4 ce d9 da de d3 dd df d9 cf cb c1 ba b7 b3 a7 a2 ac a1 a4 a8 9d 9c 9d 90 92 92 8c 94 9f 9c 95 95 8f 87 86 84 84 80 82 83 75 7b 72 72 74 71 68 70 6a 70 73 73 67 63 60 73 64 67 6d 5e 5f 60 61 6a 6f 74 77 7b 6b 6c 6b 64 71 6a 69 75 64 69 6c 67 69 6d 68 67 6a 5e 6b 5f 61 5e 5d 65 57 58 4b 33 1a 0e 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 1a 23 2d 42 5b 6e 7b 73 65 5e 65 6e 68 6f 6b 76 74 75 75 73 71 72 6d 73 6f 6f 74 68 70 70 71 78 74 7b 7b 73 7a 7c 7c 7a 76 75 7a 75 80 7a 78 73 6f 76 70 72 75 74 6f 71 71 7b 7e 75 75 7d 74 86 79 7e 7f 7e 7f 7b 84 7f 81 8b 86 8d 8a 87 91 90 93 99 95 9a 96 9a 9e a0 98 a1 a3 a5 a7 a5 a5 a8 b3 af b1 aa b1 b7 b4 a9 b0 ac af ac ab 9a 69 2a 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 02 07 11 15 1f 58 b0 cf d8 db de d8 d5 d2 c9 d0 ca bb b5 ae b0 a8 ae a4 a0 98 a7 ab 9c 9c 99 92 8d 86 8f 8d 9d 99 9b 97 8e 8b 8a 89 77 7b 7d 77 70 76 6d 64 6c 75 66 73 76 6d 6b 65 6a 73 64 63 5e 5d 5e 60 61 66 67 60 6d 76 7a 7a 6e 78 65 6d 6a 6f 6a 65 6c 6d 75 6f 70 61 60 61 66 64 60 5d 57 61 5c 5c 60 44 3a 28 14 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0d 13 24 37 41 58 6d 7b 6c 6a 62 64 66 67 70 67 68 74 71 73 71 72 76 77 77 6e 74 70 6b 6f 6f 73 70 74 7e 78 81 73 7b 7f
 7a 78 7b 7c 81 70 7a 72 74 74 75 72 6e 76 69 72 71 72 7f 75 73 7e 81 73 7a 7b 77 7a 7e 85 7a 83 80 80 80 8b 86 8a 90 8e 92 8e 92 8d 90 91 98 95 9f 90 9e 9d 9e a6 a4 af ac aa af ad a1 a6 af b0 aa ae af a2 a6 a6 9c 62 2a 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 09 07 03 06 06 0d 0e 14 53 b5 cd d3 dd dc d6 cf ce c8 c6 c3 b4 ac b4 b2 a9 a5 a1 a4 a2 a7 a8 a1 9c 98 9b 8e 95 8d 92 94 9b 97 96 92 8c 87 7f 7e 7a 7c 79 7d 75 76 6d 67 72 67 70 6c 65 69 68 73 6f 6d 69 62 63 60 60 5b 61 68 5c 75 6e 74 75 74 67 6d 68 6f 67 69 66 6c 64 62 65 69 65 64 60 5a 64 56 5a 56 59 5c 60 5a 51 40 2c 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 12 20 2e 3d 51 6c 6e 6c 66 57 5c 5c 5d 62 64 62 64 67 64 5f 65 71 76 7c 72 70 6a 69 6d 6b 6c 72 6f 7d 79 72 7e 76 79 7a 7a 80 79 74 75 74 75 7d 71 79 74 6e 6b 69 76 6b 73 71 73 6e 77 7b 74 77 70 7a 77 81 79 75 7b 7f 7e 82 7d 87 7c 7a 89 86 86 8e 90 90 8a 93 95 8e 92 94 99 92 a0 9a 95 9f a1 a3 a1 a9 aa ae aa ae b1 a6 a5 a0 9f 8c 5d 32 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 04 04 08 0c 0a 19 5a af cc d6 de d7 cf c9 c2 bf b3 bb b2 aa ac a1 a6 a5 a9 a3 a2 a9 a7 a4 a0 9e 9b 98 95 88 8e 98 9b 97 8d 90 89 7e 78 7e 74 76 73 6e 68 6f 63 67 69 65 6a 6c 6d 69 69 63 71 5f 63 61 5d 5a 5b 60 5e 58 64 66 75 78 6a 73 63 6d 6b 67 71 64 60 63 65 69 67 65 67 65 61 5b 56 5e 5a 59 56 5c 5c 5d 4f 3a 2b 13 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 19 2a 32 44 52 6d 7a 6d 67 5a 5d 5f 5f 64 5f 61 65 5f 6e 62 66 6c 6c 70 6b 76 72 6d 70 77 77 75 72 7a 78 77 7c 7d 76 7a 7b 79 75 7d 7a 72 72 74 72 74 70 69 6f 6b 70 6d 70 73 74 73 77 7d 7a 73 72 76 7a 70 72 7a 83 80 7d 81 84 7f 81 7c 8b 87 88 82 8b 85 8c 8d 8d 93 8a 90 97 96 95 92 9f 9d 9f a3 a5 a3 a1 a2 9f a4 a5 9f a5 9f 9d 95 68 31 0f 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 01 06 05 03 06 06 05 0d 08 08 0a 10 1a 4d a9 cb d5 d8 d2 c1 ca bf b9 b3 ae ab b0 a5 a5 a1 a4 a2 a6 a7 ab ac a5 a6 a2 96 98 91 8b 90 90 91 9a 92 8f 91 84 80 7b 7d 7b 7a 6a 68 72 64 5f 69 67 6d 69 65 67 5d 67 61 66 61 5e 62 5c 59 5b 5e 61 64 63 66 6e 70 6f 6e 6b 70 6a 6a 64 63 61 62 63 64 69 60 63 5b 55 5e 5e 5c 54 61 57 53 60 4c 45 2b 1c 10 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 0f 1e 1d 2a 4b 54 5f 74 6f 5b 62 57 5a 5e 61 5c 61 61 5c 60 66 67 6d 71 70 6a 74 70 6e 68 76 76 73 76 77 7c 75 73 7b 7d
 78 7d 7b 76 7c 72 76 7c 6e 76 74 6f 70 71 78 76 72 6e 75 73 75 70 72 75 73 70 79 74 6b 79 73 7d 7c 72 7d 7d 78 7d 7d 80 81 81 82 86 8b 88 81 84 8a 8e 90 8e 90 8f 93 90 99 9a 9b a1 9e a4 a0 a3 a7 a0 a1 9f a1 9b 8d 64 36 0f 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 06 09 0d 08 13 19 3d a3 c5 ce cf d0 ba c1 bb a9 b3 ab a9 a2 a8 a3 a0 a5 a3 a1 aa af a5 a5 9d 9c 92 96 95 8f 88 90 92 9d 91 8f 88 85 7e 7a 7c 74 78 67 66 66 5e 6c 60 62 63 67 6a 64 62 69 63 63 5e 5f 5d 64 55 61 63 68 64 6d 68 70 68 6f 70 6b 62 62 6a 70 66 64 64 66 6a 66 61 60 66 5c 64 54 55 56 59 64 5a 61 4f 4a 37 22 15 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 0f 19 25 2e 45 52 58 6c 64 63 5e 5b 57 5a 59 59 5d 5c 57 60 61 62 67 6f 6e 64 6c 6c 6c 72 75 75 6a 68 76 72 76 7b 77 75 7b 74 81 6f 76 74 79 70 6a 6f 66 6b 72 70 6d 72 6c 69 77 74 77 6f 76 6c 6f 74 79 70 74 71 78 84 7c 80 72 80 7d 7a 76 7e 7d 82 7d 84 7b 85 86 8e 8a 8a 8e 91 8b 88 90 92 93 95 96 9d 99 a1 9b 97 a2 9f 97 9e 93 98 87 64 30 0e 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 06 0a 0f 0b 41 90 be c8 c7 c9 b9 ac ab ad a9 ad a1 a4 9c 9f a7 a3 a3 a9 a6 ad a3 a8 9e 9a 97 93 8d 90 91 8e 8a 8c 93 89 8b 84 77 76 7a 6c 68 67 69 6c 61 65 6b 65 63 67 66 61 68 62 5d 64 5e 62 61 5c 5d 5c 5f 58 61 69 69 71 68 68 60 67 5c 60 6a 61 60 65 61 64 61 60 5e 63 5c 55 5b 5a 57 54 59 5b 5e 60 56 48 32 20 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 09 25 30 3b 48 4b 57 63 5e 57 53 5f 51 59 5c 59 5e 62 59 5f 57 5e 60 64 67 67 65 65 66 67 6e 6d 71 73 69 75 73 74 76 78 74 75 78 70 75 7d 75 75 70 71 6c 68 6f 6f 6f 74 68 75 6d 78 6b 76 79 79 7d 77 6c 70 70 76 71 6f 7a 7f 76 74 72 72 7c 75 80 81 7f 7d 80 82 85 86 8e 8b 89 84 89 8c 8c 90 91 8e 93 95 97 95 a0 9d 96 98 9a 9b 98 98 8c 6a 34 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0e 3a 94 bb be c1 b8 ad a9 a4 a5 a0 a1 a7 a4 91 9b a2 a1 aa a7 a9 a1 a4 98 98 97 95 90 90 90 92 92 93 90 90 92 86 81 79 7a 78 72 6d 69 65 60 5e 67 62 62 60 5d 64 68 62 62 61 62 59 5b 56 61 56 5c 67 64 61 62 65 6a 69 6e 64 62 5f 63 63 63 60 5b 66 64 64 5b 60 5c 58 5b 56 5c 4d 59 59 58 5b 5e 5f 45 39 1c 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 19 2c 3c 4a 53 64 66 5b 52 5e 5a 5a 60 57 64 57 5e 5d 5e 64 61 64 61 65 6c 69 69 61 64 63 6a 6f 75 74 7b 78 76 76 74
 7a 76 72 78 6a 71 78 6f 72 6e 6d 70 6e 6f 6d 71 76 71 77 75 72 75 7f 77 79 71 70 70 7a 70 72 76 7b 78 7c 84 80 73 79 73 7f 79 7d 7c 7c 81 7c 82 8b 83 8a 85 8e 82 92 96 87 89 8c 94 9a 9f 94 97 94 9d 97 90 96 94 8c 65 2f 0e 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 04 06 07 0d 11 2e 88 b5 c2 be b5 a7 ab a6 a2 a3 92 99 9a a5 9c a6 a4 b0 ad a2 a6 a5 9e 97 9e 92 97 97 93 91 92 96 8d 8f 87 84 7c 7c 78 74 6c 69 6c 6c 6b 69 5f 64 5e 65 62 5b 68 61 61 56 5d 5e 60 62 5f 59 64 62 5e 63 6a 72 74 63 67 67 62 70 60 66 64 60 68 68 63 69 5e 58 5f 62 5f 61 51 52 5b 5d 55 58 60 5a 44 3d 27 14 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 14 20 25 44 42 57 5e 56 55 5d 61 5a 60 59 55 5d 5e 57 5a 5f 54 60 64 66 65 67 65 69 66 6c 63 69 66 61 6f 71 71 72 6f 73 78 74 75 72 6b 6f 6c 74 6f 72 76 6f 68 72 6c 70 78 73 79 6e 75 6f 76 6e 7a 73 70 77 6a 70 76 78 7a 78 75 74 78 70 7a 7b 7e 7d 79 79 7e 7c 7e 81 84 7f 83 82 85 8a 88 90 8b 8f 92 97 90 92 8f 94 96 9a 9b 93 99 91 92 66 33 0d 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 03 13 25 80 ae be b8 b0 a5 a2 9b 95 9c 9c 9b a0 9f a3 a9 aa ad a0 a2 a0 99 99 8a 98 8f 93 94 90 99 9b 95 96 8a 8b 85 7e 72 6f 71 6e 6b 65 69 68 65 61 63 5e 57 5e 60 66 57 5a 58 5b 55 59 5e 5b 5a 5e 61 64 68 6a 68 6a 65 5c 63 60 67 5b 59 67 58 61 68 64 5f 5e 5b 5b 55 53 55 55 58 52 5a 50 53 5f 5c 4a 40 25 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 18 24 2c 37 43 56 52 53 5f 5c 65 5d 56 5f 5b 5d 5e 5a 63 51 5c 62 61 64 65 65 64 61 5d 61 62 66 62 69 6d 6d 65 71 70 72 70 68 6f 6c 69 67 62 72 73 6d 66 6f 6a 6c 72 6f 73 71 75 76 74 77 74 7f 7c 7b 6b 76 71 70 79 78 72 76 73 7f 76 79 71 76 7d 70 7a 75 74 7f 7c 82 7a 7d 7e 84 89 88 85 91 8a 90 8a 98 98 98 99 8e 9b 93 8b 9b 87 8e 89 6a 2c 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 09 06 0f 11 28 7e ac b4 b0 a8 9b 9f 8f 92 92 9f 99 9d 9d a4 ae ad af a0 9f 9e 9e 98 92 92 8d 8d 94 91 95 90 8d 8d 8a 86 79 82 76 6b 6d 5d 69 60 66 5f 65 66 65 57 52 64 5d 5c 55 5a 5d 59 5d 52 5f 5f 5b 5f 5f 64 60 66 67 61 5c 66 60 5a 62 5f 66 5e 63 62 6a 5e 65 5b 5d 58 51 57 4e 4e 50 4e 54 5a 59 5c 5a 4e 3b 2e 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0d 10 1d 34 40 4a 55 50 51 55 57 6e 63 5c 61 55 5d 5c 64 63 5f 5f 5d 57 60 60 64 66 60 6b 61 61 5f 66 5f 63 68 62 6a 62 69
 67 65 65 6a 6c 6e 75 6d 6a 72 74 70 72 6e 71 74 6c 66 70 7a 73 76 7e 6c 78 70 75 72 74 6f 72 78 73 75 77 72 70 74 73 7a 79 72 78 7c 73 84 7a 7f 81 7a 80 84 7f 87 83 86 82 8f 90 90 93 91 8e 8f 8a 90 98 8f 8d 91 87 69 3d 0e 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 04 0a 27 70 ae ae a9 a8 9e 97 94 90 93 99 98 a4 9e a6 a5 a8 a3 a1 a5 92 99 98 90 94 8c 8f 8c 94 99 99 92 8c 83 7f 81 78 6e 6c 6e 6c 71 5e 68 6b 61 63 60 64 5f 5f 61 60 57 5d 58 5b 5e 59 60 59 56 5f 68 6a 66 65 62 68 64 61 60 5e 62 5d 5c 65 5d 5f 61 5e 61 58 56 4e 51 47 5a 50 57 50 58 53 52 60 63 4b 3e 27 13 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 1a 19 31 49 43 56 57 54 57 59 5c 63 5d 5f 5e 57 5d 60 5b 57 5c 61 5c 67 5b 5b 66 5e 5a 61 5e 61 69 66 65 65 64 60 62 6e 6a 6e 6b 64 6c 71 73 69 7f 73 69 70 77 70 74 76 69 6f 75 79 76 79 79 77 78 6f 6b 70 71 74 74 74 74 76 6f 76 74 77 70 71 78 80 77 7d 7c 7b 74 7c 7e 79 80 7b 83 85 7e 88 8a 85 8d 8c 92 90 91 94 96 8f 8c 95 87 87 88 6a 35 12 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 00 06 06 06 0f 1e 5f 9c a1 a5 a2 92 96 92 98 95 9f 99 98 a1 a4 9c a4 a0 a1 9c 9c 91 8c 96 8f 92 96 95 99 96 8c 8a 7f 7f 75 71 74 6c 70 6d 64 66 60 6b 64 56 59 65 63 61 5e 56 5e 5f 52 57 5e 5c 5d 5a 5c 5c 62 63 67 6c 61 6c 69 61 62 62 5f 5e 5e 63 5f 5f 66 67 59 5a 5e 52 5c 59 4f 5a 5a 50 53 49 58 52 5f 61 52 41 2a 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 10 2a 38 43 57 58 55 54 51 52 52 5b 58 61 56 5f 5c 51 61 61 5e 61 55 65 5b 5c 59 60 5f 5b 60 5e 55 5f 5e 63 5d 5d 63 5c 62 69 5e 68 70 6b 69 6c 6d 72 6d 71 70 70 6d 68 69 77 6d 77 77 79 7c 79 78 70 6f 70 6d 6f 74 6f 74 6f 73 79 67 73 74 71 74 73 6d 77 76 7c 78 7e 7c 80 7d 7f 78 7c 85 88 94 8a 8b 87 8e 8c 8c 86 8e 8f 8a 8c 87 8e 89 65 33 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 0c 18 5f 9b a1 a1 99 8e 94 95 8f 91 9d 9c a5 a4 a1 a8 9d 94 9b 9c 95 8f 91 8d 93 94 9b 9a 9a 91 90 89 84 81 75 6e 71 6a 65 65 64 6d 5e 66 64 5c 5c 60 5f 5e 60 56 57 5a 57 5c 60 53 54 5b 61 5f 61 66 64 61 64 66 66 5c 5f 5c 59 5e 50 5b 63 60 5d 5c 55 60 50 59 5d 53 53 51 53 48 54 4d 4a 58 56 5d 4c 34 2d 15 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 1f 20 32 43 4b 5a 53 50 54 5e 56 55 4e 5f 58 64 56 5b 5e 53 5e 5c 5c 5c 5c 59 59 59 52 54 5f 54 5a 61 5c 5a 62 5b 66 62
 62 65 62 64 6e 72 6b 77 6d 69 72 71 70 6e 6a 69 64 6e 75 6a 73 7c 7a 77 72 75 73 75 77 75 72 75 6e 76 73 6f 6d 70 6e 6e 70 74 70 77 7b 77 6e 7b 7d 7a 78 7f 76 81 83 80 85 7b 89 89 8a 87 89 88 8e 87 87 98 87 82 85 64 37 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 02 06 05 03 00 0b 05 03 07 11 51 8e 9b 9f 96 91 96 94 95 93 9c 96 a2 9a a5 9b 9d 9a 97 95 95 8d 8f 8a 92 99 9e 96 92 90 88 8e 81 7f 74 6a 6c 68 66 6a 63 6a 60 5c 6b 64 5d 5a 5b 61 56 65 62 53 56 59 64 56 5f 5f 59 5f 68 6a 62 63 69 67 64 61 5a 5d 5f 57 64 58 62 5f 59 5c 52 60 5b 5e 55 51 50 58 4c 53 50 57 52 4d 5f 5f 48 35 24 12 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 10 18 21 31 4b 57 57 4d 4f 4a 50 5e 54 54 54 4f 58 5c 58 59 4c 4f 5e 56 5b 56 50 57 53 53 58 52 53 5e 54 5e 5b 54 59 60 5f 60 66 66 69 6d 66 6b 6f 78 71 6b 71 6e 67 69 67 62 6e 69 75 70 72 76 70 76 70 77 73 6b 77 72 72 77 6e 71 74 6f 76 72 71 77 6e 6d 79 70 7a 79 74 73 70 74 80 7a 7e 85 7f 7f 83 85 84 84 86 84 8e 87 84 87 8b 7c 7d 7d 70 3f 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 08 1e 51 89 95 99 94 8e 97 8c 92 96 a4 9d a3 9a 9b a2 97 99 96 91 96 89 92 94 95 92 99 90 86 90 87 87 7d 73 70 71 6f 6f 68 6a 62 68 61 63 63 5a 5d 62 60 59 5d 5e 5c 5c 5d 5e 5d 59 58 62 64 62 60 5e 64 5e 64 5d 5f 5c 6a 58 5f 59 55 5e 61 5e 5a 59 55 59 59 4e 56 53 50 57 46 4d 4e 4b 52 54 56 5b 4d 34 24 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 1c 2a 43 4b 51 54 50 51 52 51 4e 54 4b 52 53 4b 5d 57 4e 52 4e 5a 5a 5b 59 52 59 52 4c 4f 58 60 4e 5c 59 57 4d 54 64 60 5f 66 6b 66 6b 70 72 68 72 6e 69 68 69 6c 69 62 65 62 6d 6d 6c 75 67 74 75 78 74 75 6a 64 6f 6f 72 70 6c 76 6c 6c 78 73 71 75 6f 6f 77 6c 77 7b 7a 77 7a 7a 78 7c 7c 7e 79 80 83 84 88 82 80 79 80 81 81 7c 74 79 78 65 37 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 04 0b 46 84 90 97 94 88 89 8d 98 9b 9e a0 9b 91 97 92 93 94 8e 8d 8b 8d 90 90 98 8e 90 88 86 83 88 78 75 75 6c 66 62 62 60 5e 69 5a 61 60 64 5a 5e 62 56 58 5c 55 5a 57 5a 5d 5c 5b 5c 62 58 59 61 5e 62 63 5b 5f 60 5e 64 58 5b 5a 60 5d 5e 56 56 57 57 57 5b 58 4d 4f 53 4e 52 54 51 4e 51 4e 59 5d 49 30 20 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0c 1e 28 39 49 50 54 4c 52 55 4f 50 4f 3e 49 4a 50 56 51 52 54 52 54 51 56 58 55 59 4e 4a 50 52 54 4e 50 4b 59 58 59 65 54
 58 60 62 61 74 68 75 72 70 7b 66 67 71 6c 6b 60 62 69 65 6a 6a 66 70 68 72 73 77 7c 72 77 72 6a 73 6f 73 75 71 71 76 6f 7e 79 7b 78 79 76 70 70 74 7a 79 78 79 70 75 7e 7e 7a 8b 7c 7e 7c 7a 7f 87 80 7b 76 80 77 80 64 3f 0b 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 05 06 0f 3e 88 8a 92 90 8c 8f 9a 8e 9f a0 9e 91 94 8c 90 97 90 96 8d 8d 95 8b 8c 91 90 86 8b 86 81 7d 79 77 76 6f 6c 67 6b 66 5d 64 5e 60 67 63 61 5a 5e 64 5d 56 5a 59 5c 5c 65 57 64 5c 56 5b 54 5b 58 5e 5a 5c 56 58 57 57 5e 57 5d 5b 5e 6a 5c 5b 56 4c 59 52 59 53 53 57 52 54 50 4d 52 52 51 54 56 43 2f 1f 11 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 1b 22 29 3d 48 54 50 52 4d 4e 4c 50 4a 4c 4f 4d 45 50 4d 59 59 4f 55 55 53 57 4f 4a 50 55 4c 57 53 5a 51 51 56 52 50 57 56 5b 60 60 64 64 6e 69 6e 71 6d 70 6b 68 66 65 62 64 6a 6d 65 64 68 65 6e 6d 6d 72 74 74 6f 70 6e 72 73 75 75 70 73 79 78 7a 72 7e 7a 71 76 73 72 76 66 7a 70 82 7b 79 7a 7e 7c 7b 7a 7d 80 7e 82 81 83 7d 7a 74 76 75 57 32 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 04 14 42 79 90 96 8f 86 90 98 97 9b 9d 8b 98 8a 8d 92 89 92 92 87 8f 8b 97 90 8f 8b 89 8d 87 80 7f 7a 76 6e 6b 6e 66 6d 66 5f 64 64 5e 61 65 56 55 62 5b 58 5e 58 5c 62 60 5c 68 63 60 63 5d 5b 51 59 5d 59 60 5c 55 5f 67 58 60 5f 69 5c 5b 53 58 5a 53 53 54 5e 58 50 4f 50 51 54 50 50 46 4f 54 4b 3b 2e 2d 10 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 0f 23 36 3f 4d 5d 4e 47 43 48 4d 47 41 4b 4a 4c 51 4e 4f 4a 58 4d 47 55 51 4e 57 50 4d 4d 50 4d 4c 4e 50 54 58 55 4b 53 58 54 54 59 61 60 6b 68 72 6a 6c 6f 6a 64 65 68 63 67 60 5c 64 62 6b 66 5f 68 66 67 6c 69 6f 72 73 70 6b 6f 6f 73 70 6c 71 7b 6b 76 77 6e 74 70 74 76 71 6f 77 73 72 78 75 76 74 7b 76 78 75 76 75 74 79 78 75 72 78 75 62 3b 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 15 30 7d 82 87 88 7f 90 97 9a 9a 93 90 84 88 86 88 90 89 82 85 83 90 90 8a 8c 85 82 82 81 7a 73 75 74 6c 62 6c 69 62 63 69 5b 60 5c 56 63 5b 60 5f 5e 5c 58 5a 5f 58 69 5c 5d 64 5e 60 54 4b 53 51 60 59 5b 5e 63 5d 5f 5b 5c 6a 6f 6e 5e 54 56 4e 49 4c 50 54 54 4c 50 4d 50 49 50 4d 4a 4a 4e 45 30 23 25 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 16 1f 2a 3d 50 59 4b 43 46 4d 48 56 4a 4b 4e 48 49 57 4e 51 4e 4b 4a 52 4d 5d 55 4e 4f 4f 52 4d 53 4b 4e 4a 51 4c 57 56 51
 53 59 5b 5c 67 60 6d 64 68 70 65 66 69 62 5d 66 64 61 69 5f 6c 68 63 63 66 69 69 71 68 71 76 76 70 70 6f 71 73 6d 6e 75 73 75 73 74 73 6e 6d 6d 70 79 74 6e 6f 76 6f 73 6f 72 7f 74 73 79 70 6c 6c 74 72 70 7f 6e 79 64 34 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 04 06 0d 3a 70 7d 86 90 88 9e 98 96 94 8c 8a 8c 85 7d 85 7e 8a 8c 87 90 92 8b 83 88 8a 81 87 84 73 79 79 66 6e 6b 6c 60 64 5d 60 5d 61 5c 5e 61 5e 58 5b 5b 5b 5c 56 62 64 62 5f 67 65 67 59 4e 4a 54 55 52 5a 5b 5a 5e 55 60 5b 64 71 74 69 61 53 50 4c 50 51 4b 54 54 51 51 4f 4b 4f 48 4c 47 4b 4b 3d 31 27 1e 13 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0c 23 23 33 47 59 4f 52 43 4a 4e 51 4b 4a 42 49 48 4b 54 4d 4f 52 53 48 49 54 52 50 49 4e 48 4d 5b 4f 4a 57 53 59 52 57 58 57 50 53 59 55 62 63 62 68 64 67 6c 64 66 5f 65 64 6a 61 62 63 59 65 65 61 65 66 65 6c 6c 64 69 6f 6a 63 6f 73 6b 67 6e 6f 73 76 70 76 72 78 6b 72 74 72 7a 73 71 75 6f 75 7b 6e 78 74 76 73 72 73 7c 74 6a 75 71 70 6c 68 34 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 07 06 05 0a 2e 77 8a 8e 8b 8c 99 97 8e 93 95 91 8e 87 80 84 88 83 85 87 89 89 8b 8e 84 86 86 81 82 71 76 71 70 6f 69 6d 67 62 61 61 64 61 5e 63 65 5e 60 60 64 58 5b 68 5f 62 5d 65 63 66 60 55 54 53 55 61 59 57 5e 62 5b 5a 5b 56 63 70 6d 64 5c 55 57 53 54 56 54 57 59 52 54 51 4b 4c 4d 4f 53 44 47 3b 24 21 18 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 16 10 21 36 40 54 58 50 4e 47 4e 4f 47 4b 45 51 4a 51 52 4f 50 52 4d 48 50 4b 51 53 50 48 4a 49 4f 54 4e 51 54 53 4c 51 56 51 4b 5e 54 50 5d 67 5d 65 69 68 5b 5a 61 62 5e 60 65 5d 57 62 61 60 60 67 64 61 64 67 67 6c 6d 68 69 6f 68 6e 6c 65 65 6a 69 66 65 6c 73 6a 75 73 77 71 6f 62 6c 72 6b 6f 73 6c 71 71 68 71 78 7b 6d 70 73 6a 7e 6f 6e 65 3c 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 03 00 0b 2e 6e 87 8f 96 95 9e 98 8f 90 8d 85 84 82 87 85 83 8e 8b 86 87 80 85 87 84 87 87 7e 76 7a 74 74 6d 65 6d 61 64 61 5d 64 5d 5c 54 5b 65 5e 60 61 50 57 5a 5d 65 54 5b 5e 61 53 60 49 4f 4b 4e 5b 59 5a 58 5e 5f 58 59 50 5c 5e 67 60 59 59 54 56 54 51 4e 52 55 4f 51 49 4e 4c 50 4d 52 41 3a 31 24 21 14 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0d 1a 2f 3a 47 58 49 4a 47 4c 48 4d 4e 4b 4c 4c 4b 4d 51 4e 4b 45 4b 52 54 4f 50 4d 4c 4a 50 4e 50 4f 4e 4f 53 50 51 51 4b 54
 4d 4f 54 53 55 5c 5a 5b 5d 5d 5c 56 5f 63 61 64 64 58 5c 65 5b 64 63 55 68 5b 66 5f 66 67 66 65 6e 6a 69 69 5c 62 6d 62 61 6e 6b 77 6c 72 6d 64 74 6f 71 72 74 73 73 6d 6a 6d 6c 6e 73 6b 77 76 75 74 75 72 74 70 77 66 3c 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0c 25 73 87 87 90 94 9f 8f 8a 86 85 89 84 86 7b 86 87 83 81 88 8e 83 86 77 84 7d 81 7b 76 7d 6a 6b 69 69 6b 67 6a 61 5f 5a 64 5a 5e 5f 5c 5e 55 59 59 5b 64 55 60 5d 65 60 62 56 4d 52 4f 4d 54 59 55 5c 57 53 5a 51 5e 5a 5b 5f 5f 63 54 5c 45 4c 54 4e 46 54 4c 41 4e 55 45 4d 4f 4e 4b 3f 44 30 24 1b 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0e 16 31 36 54 5e 56 48 44 4c 46 50 44 4a 4d 46 50 4b 48 4d 4b 50 45 4e 54 4d 4e 4f 4d 50 4a 50 51 4d 4e 4e 53 4f 4c 52 53 4e 50 54 55 53 5d 5f 63 57 59 5b 5c 5e 5b 5f 55 5b 5c 69 67 62 5c 5f 5d 6a 5f 64 67 5e 62 6b 67 6c 65 6b 71 6e 69 6b 68 65 66 68 72 6f 72 72 6a 6d 72 6b 6f 6e 71 74 6b 6b 6f 72 71 71 72 6f 71 77 70 73 75 72 72 73 7a 65 44 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0a 06 1d 69 87 8d 90 91 9e 97 90 8d 86 83 88 7c 80 81 82 88 84 85 80 7e 7f 7e 86 7f 7c 7d 73 73 74 70 65 64 64 60 64 62 62 61 64 62 5e 62 5c 59 5e 5d 55 60 56 67 5e 5f 66 5b 59 4e 50 54 53 55 4d 58 56 5c 60 59 5c 4e 5c 5a 5e 54 59 53 53 4c 4c 4e 53 50 52 4d 51 51 55 57 4e 50 4b 53 4c 44 38 23 20 23 14 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 17 20 2f 3a 4a 58 54 53 49 48 3f 4f 4b 54 44 4d 4b 4c 52 4f 4c 4a 49 4b 50 4f 50 4c 4e 53 51 4c 50 4c 4c 55 4e 51 50 49 4e 4e 4d 4b 55 53 51 5c 50 55 59 60 5b 56 57 5a 5e 58 5f 5c 61 5f 5b 60 63 68 5c 55 61 5f 5e 5a 64 6a 6d 6e 66 6b 67 71 5c 6b 67 63 64 68 6a 6f 70 71 73 70 74 68 6b 69 6b 70 6b 68 72 6e 70 7b 74 70 74 7a 7d 76 74 77 6e 67 3e 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 0d 22 66 7f 8c 92 8d 95 94 90 89 86 85 81 80 79 7e 84 87 86 84 86 83 84 79 84 79 84 7e 6a 74 6c 6e 6e 6a 63 61 66 61 60 62 56 63 5f 64 5c 5c 5c 5a 5c 62 5b 5b 53 59 60 58 55 4c 50 51 4e 4a 4d 4f 57 50 4d 52 50 56 51 5e 59 59 56 55 57 4b 53 53 4d 4e 50 50 4c 52 4f 50 4c 4d 4c 4c 4f 48 37 2a 22 1e 12 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0b 1e 1c 2b 3d 4d 55 4f 53 41 46 47 47 4f 46 4b 51 3f 45 4a 49 45 4d 4f 4d 43 4b 47 42 55 46 4d 48 4a 4d 4c 53 4d 4f 53 4b 48 4b
 49 58 51 53 4b 54 4f 49 53 4f 51 58 57 4b 5c 5a 56 5f 5f 66 5e 60 62 5f 5f 64 59 57 5f 5f 5e 61 65 61 6b 69 64 69 67 62 66 62 66 6e 62 6e 69 72 69 64 71 72 66 6e 72 65 6d 70 74 77 71 78 75 76 7b 76 79 78 6d 77 76 6c 40 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 1f 65 85 8f 90 92 8b 8f 90 8a 8b 84 7e 80 88 7f 88 84 89 7b 84 77 85 79 7e 76 7d 7e 73 79 6f 6a 6f 5c 65 6b 63 67 59 66 62 60 5f 65 5b 59 59 5b 60 5f 5e 55 5e 59 59 56 5b 4d 44 47 4c 4d 50 4b 49 50 50 4f 4d 4b 51 53 51 59 5c 4e 4d 48 4b 4c 50 4c 54 49 49 50 4d 4b 4d 4c 4f 43 4d 3b 39 24 1c 19 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 19 21 2f 3b 50 63 58 55 47 48 4b 51 44 45 49 43 48 4b 4a 47 4f 44 50 46 44 43 46 4e 4e 4b 4e 4e 41 54 4b 46 51 4e 49 49 4e 54 49 55 4e 4e 53 54 57 53 4b 4e 50 51 52 5f 54 56 52 5b 5b 5a 5c 58 5c 57 61 5f 58 64 5f 5f 63 65 64 6d 61 62 5e 64 64 68 6c 65 6b 72 5e 66 69 60 69 6d 70 6a 6b 66 68 70 75 6e 77 6f 7e 74 7f 7d 7b 7e 7c 7d 7a 76 72 66 3c 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 60 84 88 8d 90 90 93 8a 8a 82 80 83 78 7a 78 80 88 81 7f 86 7a 87 7f 7b 7e 7b 77 73 6a 6e 69 67 5e 63 66 61 5e 66 5a 65 68 5f 5f 5e 5d 5e 60 5a 5b 60 5c 5e 5e 57 4e 4a 4c 51 4b 51 47 49 4d 51 52 4e 52 4b 4a 4e 51 52 50 5b 49 56 4d 4d 54 4a 54 4f 48 53 50 54 4f 54 53 4c 4c 47 40 30 23 20 15 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0b 1c 3a 41 57 65 58 55 46 4d 4d 4f 4a 51 4e 4e 4f 4e 50 53 53 45 49 49 44 4e 50 4c 4c 45 4b 4e 4a 4f 52 43 45 48 52 4d 50 4a 49 4d 50 56 50 4e 52 56 50 55 4e 4f 55 50 56 54 52 5c 5a 5b 59 58 63 53 5d 5d 59 61 5d 58 62 65 61 66 68 65 5e 65 66 65 66 61 69 6b 73 69 6a 6b 68 69 6b 76 70 74 75 79 75 70 81 74 76 7f 87 83 7e 79 7c 74 73 7a 77 6d 43 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 1e 57 86 88 8d 88 8e 95 90 8d 7e 81 7a 81 83 84 88 7d 7f 7d 7e 7e 7a 7a 7a 7b 79 75 6c 6c 65 63 63 6e 64 68 64 61 5d 5f 56 61 5f 58 66 4f 5f 5b 5a 5e 5d 5b 5b 53 4d 50 50 4b 50 52 4b 49 4e 54 4c 49 4d 4e 46 47 54 4d 4a 4e 57 50 4c 4b 4f 54 47 4f 50 4c 51 4c 50 4c 50 55 4a 50 45 33 35 21 27 13 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 04 0e 10 24 26 38 51 5f 55 50 4d 4b 45 46 4e 44 42 4e 47 47 43 4f 4c 45 4c 46 47 4b 44 4d 43 45 48 41 49 48 4c 4f 49 49 50 4b 4c 48
 50 49 49 4c 4b 50 51 54 4c 52 48 57 4f 4d 4f 54 4d 4f 56 57 58 54 5c 5f 63 5e 56 5b 5c 5f 61 63 61 5c 55 69 65 5f 5d 64 71 5b 72 66 5f 6a 63 6d 66 66 6e 6e 6a 74 71 72 7c 75 7d 7d 7d 7d 75 7e 7e 7c 75 78 71 77 73 71 47 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 18 56 7b 84 86 84 8f 8f 90 8d 85 80 7a 77 82 80 85 86 87 79 81 7f 80 74 71 77 75 6f 6c 6b 6f 70 69 62 5e 63 62 5a 60 5d 61 5b 56 5b 5a 55 5a 5e 5c 56 5b 5e 54 4b 50 4e 49 4c 47 47 54 41 42 4c 4d 51 48 41 49 44 4d 48 50 4c 53 49 57 41 4e 4a 4a 4e 53 4a 51 4a 4f 50 4f 4a 46 4e 4e 32 29 1c 1c 12 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 17 23 28 3a 4d 5d 5d 5a 49 49 4a 4e 44 4b 44 4e 43 4c 45 48 4e 4d 40 4a 48 4b 4c 44 41 3e 44 45 44 4c 49 4a 46 49 4a 4e 4e 4e 47 50 40 4f 54 4b 57 52 54 4e 4d 51 4e 4f 56 50 4a 52 50 51 51 50 52 5a 57 59 62 5c 5c 5a 52 5a 60 5f 65 62 5f 5d 60 5e 68 69 69 6b 64 70 72 6f 70 70 69 79 79 6f 79 7c 75 7a 7d 7e 75 7d 7b 82 75 73 7a 79 76 7b 79 70 43 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 17 56 81 88 8b 8a 8c 8f 84 81 83 7c 80 7d 79 7f 83 80 79 78 7b 7c 80 79 7c 6f 73 6a 73 68 64 62 66 65 61 61 55 5c 64 5e 5c 60 5d 5d 5e 51 55 55 5b 5e 5d 52 53 52 4f 4c 4e 4b 49 4a 49 52 49 53 4b 4b 4a 50 52 4d 49 50 50 4b 4a 57 50 44 49 4b 50 52 4c 51 4f 47 4b 4d 47 4a 49 4e 43 3c 2e 20 11 0e 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 09 15 23 1d 33 4b 56 58 56 45 48 42 4b 4d 48 4b 4a 47 43 4a 40 47 46 41 46 43 45 48 45 46 44 3e 46 47 48 4f 4c 48 48 4a 45 49 47 4b 4c 51 48 49 50 53 4a 4a 52 4d 4d 52 57 4f 49 50 52 53 53 52 51 55 52 52 56 57 54 4f 54 5e 5a 62 5d 5f 5a 5c 5d 60 64 66 66 6e 6c 6a 70 6d 6d 74 72 78 75 73 79 7b 7d 78 7a 79 76 72 7a 77 75 71 75 77 70 6f 74 72 68 40 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0f 4b 86 82 89 80 82 88 90 8b 8a 80 80 73 75 85 83 79 7f 7c 7f 78 7a 77 76 6d 70 68 6d 6d 67 5f 65 68 63 63 5d 59 56 5d 59 5c 58 5e 53 60 5a 57 5a 56 58 54 47 4e 50 4c 4b 49 49 49 49 49 50 51 44 45 4b 4d 5a 4a 50 49 48 45 53 52 57 51 44 49 44 4d 4d 49 53 4c 51 50 4c 52 48 49 46 36 25 19 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 09 09 20 20 34 4c 54 5d 53 53 41 4a 4e 44 40 3d 43 49 48 4a 45 4c 3f 48 3c 45 40 44 4b 44 47 41 41 47 49 45 49 53 54 4f 4c 52 49
 48 45 47 47 4c 47 51 53 50 4f 4f 4a 47 50 4a 53 56 51 4a 53 4c 50 55 55 5b 55 54 4c 50 58 57 54 58 54 53 5b 59 5f 51 5d 61 60 65 6e 6b 72 6d 75 77 76 75 73 6c 74 70 72 6d 6b 76 70 79 6d 76 77 6e 70 7e 75 6c 72 71 72 44 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 4a 7c 8c 8d 85 85 89 88 8e 8d 8a 85 83 77 80 80 81 84 81 80 80 72 77 77 68 76 6b 6e 6b 66 69 68 63 61 60 62 57 58 55 56 58 55 5b 57 5a 58 58 58 55 54 4d 4b 4f 4a 43 4d 4c 4c 54 4c 48 4a 46 45 4b 4d 45 47 47 46 40 49 4f 49 4a 47 45 4a 51 43 4a 49 52 43 53 54 4a 4e 4a 4b 4c 3e 2a 1b 18 0f 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0d 13 1d 25 2d 42 4e 58 56 4e 50 49 49 49 43 48 43 44 47 43 4c 41 44 43 48 51 44 48 47 41 48 43 41 4c 47 47 4b 4c 4e 51 51 49 4e 4f 4e 50 4c 51 4e 54 59 4a 53 4c 4c 51 52 45 4e 52 4b 59 52 4b 4e 4f 50 54 5d 4f 5b 52 54 59 5b 5d 62 5e 5c 50 54 56 57 59 60 65 69 6a 6f 74 76 77 70 6f 70 6b 6c 68 63 6d 67 61 6e 6d 6b 6f 6b 70 69 76 7d 70 6d 75 63 45 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 47 79 87 88 80 89 85 83 8c 94 90 91 84 86 8d 84 8a 79 7b 78 79 7c 74 77 70 6b 6a 68 64 65 5b 5e 5a 5a 67 63 60 61 5a 60 59 5e 62 54 54 55 52 4f 55 4e 51 4b 4e 4d 4a 4a 4c 49 51 45 45 48 4a 45 4e 4b 4b 4d 44 4b 4b 4d 54 4f 4a 4c 4b 47 4f 49 50 50 4e 46 4c 4c 50 57 4e 50 4c 44 2a 20 13 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 06 14 13 22 25 3f 4c 5a 57 45 44 4c 45 41 43 46 49 4b 49 50 4b 48 3d 4c 3e 4a 3c 42 48 4c 3e 40 44 3e 46 49 4b 4a 46 46 4b 47 4e 47 4e 4b 48 50 4a 50 49 55 4e 43 4b 4c 4f 47 52 51 54 4e 55 51 55 51 51 48 4e 56 57 5a 54 57 5c 54 55 5e 58 5b 5f 55 58 62 5c 67 67 6d 6e 75 75 6a 6a 62 65 69 6c 69 68 6e 6e 78 6b 6a 70 6a 6b 6e 69 6b 6f 68 5f 6a 61 42 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 40 7f 85 91 83 89 89 86 7c 88 8d 86 86 88 8c 8e 80 87 81 7f 76 7c 73 73 6d 6e 69 6b 61 64 6a 61 5e 60 5e 55 5d 5a 5a 5a 5c 5a 57 64 5f 53 56 55 4e 4f 55 45 4a 4f 4f 53 51 53 4b 43 43 48 4f 47 48 4b 49 41 46 49 4c 46 45 52 4e 56 4d 53 4b 4f 51 4e 4a 4d 4b 4e 53 52 51 4e 40 3f 33 1f 15 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 12 19 1d 2d 2f 4c 4c 49 4d 49 4a 49 4a 41 41 45 48 49 48 41 49 37 34 3c 3e 44 45 39 43 42 3e 3c 3e 45 47 47 49 54 41 40 44 4a
 45 4e 47 48 4d 51 4c 50 4f 4e 45 52 4a 42 4e 50 4d 50 4f 50 52 48 52 4f 53 4a 4d 50 4e 52 5c 57 56 57 52 5d 53 5a 57 57 64 56 60 68 70 72 6f 6f 6b 5f 63 61 63 6a 68 65 6a 5f 67 67 64 69 6d 67 6a 67 6c 68 67 5f 69 5e 43 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 3b 74 8b 8b 7c 80 81 7e 84 84 79 85 87 81 84 80 8d 89 83 84 7e 72 71 6f 65 6f 66 67 66 61 64 63 5d 63 59 58 58 5a 52 58 51 5d 5a 58 56 50 55 5a 4f 4f 4a 4a 3d 49 48 46 48 45 44 51 44 45 50 41 49 48 48 46 4b 46 51 48 47 51 4c 49 4e 45 48 4b 52 4b 4f 47 4e 50 4d 52 4e 44 4a 35 2b 19 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0a 1a 1a 26 31 3b 4e 44 4a 4b 4b 45 41 43 4b 41 4c 45 47 3d 42 44 42 41 3e 45 49 44 3c 41 4f 43 40 49 40 49 48 4d 4e 4d 50 4d 4c 45 46 49 41 4a 45 4a 4f 4d 4a 4d 4c 51 42 4e 50 47 50 4c 4b 55 48 52 4e 56 51 53 4e 55 56 55 52 59 55 5c 53 55 5d 61 5e 65 70 69 67 6a 65 65 68 60 63 64 64 60 64 64 68 6e 6f 69 64 69 62 6e 6b 6c 6d 5c 64 61 62 63 41 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 3a 73 81 90 81 89 85 7b 82 7e 7e 81 7b 7c 83 82 88 84 7e 81 7a 7d 6b 70 72 71 66 6e 62 67 63 5d 55 60 5a 5d 5c 5d 5a 5d 5d 53 57 51 4b 49 4e 49 4f 4f 4a 45 4b 4e 4a 4e 48 42 4c 44 45 4b 48 47 4d 4b 45 3f 49 40 43 51 47 4c 4d 46 54 4e 47 46 4a 4d 49 4a 46 4c 53 4f 54 42 40 39 22 15 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0f 15 1c 20 2d 3b 45 43 4b 4b 47 53 48 47 47 4a 43 4b 47 4a 42 46 47 45 41 40 3e 4b 49 3e 44 39 40 46 48 49 4c 50 46 4a 4a 4d 4e 55 4f 48 49 46 50 4c 49 57 53 4d 4a 4d 4a 46 4a 50 4c 55 4d 52 57 53 5a 4b 4e 53 5b 53 59 59 57 5f 55 64 60 60 5a 64 61 6a 67 6e 6d 66 69 67 5b 69 68 5c 60 61 65 66 62 65 6e 6d 67 6b 69 68 66 65 65 68 64 65 61 5c 45 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 38 6f 7e 88 7d 83 83 86 77 80 84 81 7c 80 87 82 82 8c 83 7f 84 7d 75 78 73 69 79 73 69 6a 6e 6a 5e 61 5f 5c 59 5a 58 59 5b 5e 5c 5d 54 4b 56 4d 52 4f 4a 45 3f 4a 4a 4c 50 47 46 4b 44 49 4e 4d 4e 4d 4d 4b 4f 4f 58 56 49 4c 41 54 51 50 51 56 45 51 51 4f 57 4a 54 50 4a 46 3a 2e 20 0e 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 18 17 1c 2e 2f 38 48 4a 44 46 44 4b 47 43 4a 3f 40 48 44 3a 46 41 45 41 43 44 42 41 42 40 3e 40 3c 3e 41 45 50 42 42 40 48
 51 55 4b 47 4d 44 4a 4d 49 4d 41 4e 4f 49 4b 4b 43 50 48 52 47 50 4f 4d 4d 46 50 54 4c 51 58 5f 58 5a 55 55 61 63 54 64 60 68 69 65 66 66 60 50 65 5b 5f 66 62 61 65 65 66 66 58 5c 61 60 64 67 6a 61 61 59 5e 62 5c 5d 47 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0c 2a 75 83 84 81 80 7a 74 7c 76 79 7f 7b 73 7c 6e 7c 7e 82 83 7c 79 73 79 6e 74 6f 6f 6e 69 67 65 64 5b 5f 5b 61 5f 58 56 5a 52 59 53 4d 4f 51 4e 4a 49 44 43 47 3e 4a 48 4a 47 47 49 48 41 3f 45 53 4e 51 47 4a 46 48 4f 4e 4d 4c 4e 47 4a 53 43 4a 4e 52 51 53 4d 50 52 54 41 3a 26 18 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 0b 18 21 2a 34 3b 44 47 4d 4d 49 4b 42 4a 45 44 43 39 43 3e 40 45 40 46 44 44 40 4b 3f 42 44 40 39 44 3d 47 49 4c 53 49 46 4e 42 4c 4c 4d 48 4a 4c 50 46 45 46 46 4b 4d 4d 49 4e 4b 4c 44 4b 46 4e 48 4e 4f 51 52 56 54 5b 5f 5c 68 64 5f 5a 63 61 67 69 5a 5f 60 59 60 5c 56 59 63 60 62 5e 63 60 68 66 5f 5f 63 69 61 60 61 66 5c 59 54 5d 57 40 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2d 6b 77 7e 76 70 75 79 72 70 73 74 7b 74 78 79 79 7a 7e 7b 7e 74 77 74 6f 6c 76 69 67 66 65 66 63 61 69 5f 5a 56 5a 59 59 54 59 4b 49 4c 51 4b 4d 46 47 4d 49 4d 4b 48 46 45 4b 42 44 4a 50 40 42 44 4d 43 46 50 49 45 4b 49 49 51 4a 50 4a 4a 4f 44 4e 4a 4f 4f 4e 4f 45 45 2e 20 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 14 22 2f 36 3f 4a 49 4d 4c 42 4c 45 49 3f 4b 41 4b 3d 42 3c 3e 44 3e 3f 48 41 3e 3e 42 45 45 50 4a 44 47 3d 4b 54 48 50 54 50 4a 46 44 41 47 40 50 45 49 51 49 51 45 49 4d 54 50 4c 4b 49 50 4d 4e 57 51 5b 5c 4f 5c 5e 5a 5f 64 5b 5f 63 60 62 5a 5e 5f 63 5b 5e 60 5f 60 60 56 5f 67 6b 5f 67 69 65 68 69 69 63 67 57 60 62 5a 54 61 57 54 48 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 29 5f 79 74 6c 71 74 75 75 7a 6e 6e 74 7b 7d 7b 7f 7e 77 7c 74 75 70 76 74 6f 64 69 63 5f 6a 5e 5d 5f 5b 59 58 5c 5b 51 56 51 53 4b 4b 51 48 54 4f 51 4a 48 42 49 4a 4d 51 48 45 46 43 45 4c 47 49 52 50 53 45 4b 4a 48 4f 58 4e 51 48 4e 47 4f 4d 52 50 4f 4f 4c 56 50 4a 38 36 22 04 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 1c 1a 22 2e 38 4b 4b 4e 4f 4b 49 47 4c 3f 49 44 49 45 3a 3a 44 3d 46 44 47 48 44 42 46 48 47 49 40 3f 40 44 46 48 4d
 4a 53 4c 48 4e 4d 49 47 4e 41 4b 44 4d 51 47 46 52 49 4c 48 4f 4f 49 50 52 4d 49 49 55 52 53 5d 60 60 5a 61 4f 5e 60 57 61 55 5d 5f 66 59 56 5a 5d 61 5b 64 5e 5e 64 59 66 63 5d 5c 5e 6c 63 5f 62 67 5c 5f 54 59 59 55 44 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 1e 5e 75 75 69 74 76 64 78 6f 7b 76 74 76 71 78 72 6d 71 6b 6e 6d 6e 6f 65 6b 63 68 63 61 5d 54 59 5d 5a 5e 58 58 57 57 56 53 4d 4c 47 45 4d 51 49 4c 45 47 4e 4b 4f 49 4a 47 43 4f 45 4c 4d 52 49 50 4d 42 42 46 4b 44 49 51 4a 4b 47 4c 49 4b 4e 4f 4d 4c 4a 58 4f 50 44 3a 2b 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0e 14 23 24 30 3f 49 44 4d 48 4d 41 41 49 4a 48 4d 48 41 45 43 42 41 40 45 44 47 40 4c 44 40 47 3d 41 46 48 4d 4b 40 47 4e 48 40 4a 46 44 40 44 46 4b 40 44 46 41 4b 48 49 48 45 4b 48 55 45 4f 4a 4e 4b 51 52 54 61 5d 5e 63 55 5f 5e 5c 54 5c 52 5e 5f 53 55 58 5b 59 5e 54 4d 59 58 5c 5d 5c 62 5d 5f 55 63 65 65 5f 58 55 54 52 57 52 50 42 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 52 6d 6d 6a 6f 69 6c 66 71 69 71 70 75 75 6f 76 7c 73 77 70 75 6a 6a 64 5f 62 5d 55 5e 5f 5f 5b 5b 57 55 4e 5b 51 5c 50 4b 50 50 4b 47 4c 4c 47 41 42 45 4a 4c 49 4f 46 4a 42 48 47 4e 44 43 49 49 46 4b 45 4d 52 53 53 4c 4e 49 4c 50 52 4b 4e 50 4a 50 51 4b 53 45 3d 2d 1f 14 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 17 19 2a 2a 37 4a 4f 4f 47 4b 4e 44 3f 43 48 47 42 40 3c 40 45 44 43 49 43 43 3e 39 47 44 44 45 3e 41 48 4d 47 47 4e 4e 4a 4a 4a 4c 43 4e 43 47 42 45 49 4a 42 43 4c 46 4e 44 47 4e 49 52 4b 4d 4f 46 47 59 4f 57 5a 51 51 5c 58 5b 5a 48 53 5b 5d 5e 58 5f 50 58 55 50 56 5e 54 57 5f 56 5b 57 62 61 58 5e 59 59 56 5e 5c 60 59 54 58 54 44 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 20 4e 70 73 70 6b 69 6c 64 6f 6d 6f 6f 6a 6e 73 71 73 6a 65 6f 66 62 6a 5e 60 57 65 53 61 60 5a 5e 5c 57 58 4d 53 51 57 4f 50 4d 46 47 4d 50 4b 44 4a 48 4f 4f 4d 47 45 46 42 43 48 44 4f 45 49 49 4e 46 49 4c 4a 4a 46 50 50 45 51 4c 4f 4d 4e 53 4c 52 52 47 56 45 4a 3f 2a 1c 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 02 11 16 22 34 3b 3e 46 4d 4d 54 4e 48 4c 44 4a 51 42 44 46 41 40 46 47 45 43 3a 44 41 46 4d 4a 44 48 46 45 44 43 48
 47 4e 51 4d 4a 49 49 4a 43 47 47 4f 50 4b 46 3d 4d 46 44 4b 45 48 40 46 48 4c 4a 53 4a 4e 4e 52 58 55 50 56 53 4f 48 4d 57 4f 56 5f 5d 4f 59 58 56 58 56 5c 52 5a 64 5c 53 5f 5e 61 5c 5f 5b 5c 5c 63 5e 53 59 54 5c 56 47 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 17 50 69 6b 63 65 6a 6b 6a 6b 65 69 6a 67 73 6e 71 70 70 6d 64 60 63 63 55 5d 65 58 5c 54 53 5b 51 53 59 4f 5b 5b 58 56 54 50 54 50 49 42 51 4b 45 4a 42 4e 4e 4c 41 4d 4a 44 4e 45 46 46 45 45 4a 4e 47 4b 4b 53 4b 4c 4f 51 4b 49 57 4c 47 47 52 54 53 55 48 4c 4a 44 3f 2a 15 0b 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 08 09 13 14 24 35 3f 4d 56 51 4b 46 4d 43 49 41 47 3e 4a 40 47 4d 46 45 46 3d 3c 42 3c 49 48 44 34 3a 46 4a 45 43 4d 4a 4f 4a 47 4a 4e 42 41 44 46 4b 44 4f 46 54 49 43 42 50 44 4b 49 48 4f 50 52 45 51 46 4c 52 54 52 56 57 56 56 52 53 4b 53 50 57 53 51 5b 5a 51 50 5b 59 4f 57 5b 60 5d 56 56 58 5d 55 5c 58 59 5a 53 58 58 5c 52 56 50 47 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 51 5e 65 65 65 6b 6a 6c 6c 66 68 70 66 70 6f 63 6d 6b 65 63 60 5c 5f 62 57 5a 52 56 54 59 5a 57 5a 57 4c 50 53 52 51 4d 4f 4d 4b 4c 4e 47 4b 45 44 48 4b 4d 44 3f 47 47 4a 49 43 45 49 45 4a 4c 4e 44 47 4a 4f 4c 4c 45 4d 4e 4e 4f 49 45 4b 51 4b 4c 4d 47 51 4d 3e 2d 1c 08 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 0e 1b 28 2f 2f 51 51 52 50 46 46 47 4c 48 45 47 44 45 41 45 44 41 41 44 44 3d 3e 43 44 49 43 4a 4b 3e 47 44 49 56 4d 49 4b 47 4d 49 44 4b 4e 47 52 3f 52 47 46 4a 46 43 4d 45 41 4e 46 4a 4a 52 4d 4b 50 53 54 56 54 53 50 49 49 4c 52 55 53 50 50 51 55 58 4e 56 4d 55 53 55 4f 53 4f 4e 5a 59 57 59 5e 5a 55 56 58 59 50 50 56 53 4f 47 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 45 6a 69 67 6d 65 67 6e 6c 6a 68 6e 67 6c 64 6e 62 5d 60 63 5e 5c 5d 5b 5f 59 5d 60 56 58 52 52 50 4d 4b 52 4f 50 51 55 54 55 49 53 56 4e 4a 49 45 42 4d 49 40 4d 48 45 43 44 4a 42 46 46 48 4b 4c 54 4a 4b 4c 48 44 4a 5c 4a 4d 4c 55 51 4c 52 51 54 4b 49 47 47 35 31 14 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 12 1e 20 2d 33 3d 52 4e 54 48 4a 45 48 4f 4b 49 46 39 41 42 52 41 4b 48 44 3f 3d 49 44 42 42 48 44 48 44 3b 48
 4b 40 46 46 47 49 3d 42 49 48 51 54 47 43 49 40 46 47 44 51 49 46 4e 3f 4c 4b 46 4b 49 55 5b 55 56 51 56 53 4d 51 4e 51 4f 4d 4b 4f 51 4b 53 51 52 54 54 4f 52 55 4d 54 50 5e 59 5c 52 58 52 54 5b 5c 56 4a 52 53 52 54 3d 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 4f 5d 69 58 5f 63 63 64 66 69 66 66 66 66 62 61 65 64 5b 5c 58 58 5d 57 53 4e 50 55 52 57 54 4d 50 58 51 54 4a 50 4c 52 4b 4d 4d 41 50 4a 51 45 48 4b 45 4c 44 4b 4c 46 44 42 43 45 49 46 47 4b 4f 49 52 4c 4e 43 45 51 52 55 52 50 53 49 4b 4a 49 4b 54 4b 46 42 31 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0e 12 1f 26 32 3b 42 4b 4e 4a 49 4c 4b 4d 50 4e 4d 48 44 42 41 3d 46 42 42 40 39 38 48 3b 3d 45 40 40 40 47 47 43 49 44 45 40 42 40 44 41 47 41 50 48 3f 40 45 3f 48 43 4d 40 45 4c 53 4f 4c 4f 4b 48 44 54 52 50 56 4c 4a 51 49 46 49 49 48 4b 4d 4a 57 57 52 52 4e 52 52 50 4d 53 4b 50 51 56 5b 57 5b 51 54 53 57 58 51 52 4c 59 4f 42 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 3a 64 6b 68 60 69 5e 66 66 64 61 5e 61 5c 59 62 59 5b 54 52 5c 53 58 57 4f 4e 58 4d 58 50 4b 51 4f 51 4b 49 4f 52 4f 4d 43 42 4e 44 46 41 49 47 41 51 4d 42 4b 44 46 44 46 42 3e 47 4a 4b 4d 4d 43 42 4e 46 4c 4a 4a 4a 4c 42 4f 4a 54 53 4f 55 4f 53 56 4b 4a 3d 25 14 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 13 21 22 24 3e 3f 43 4f 49 49 4c 53 53 4f 42 49 44 42 45 43 45 3e 4b 3f 42 47 43 3e 3e 4a 47 46 4b 3c 49 4a 49 46 48 45 44 48 43 44 49 49 51 43 41 43 49 42 3d 45 49 4c 46 47 4c 4b 47 45 49 46 4d 4e 53 54 58 58 4e 50 4a 4f 51 4c 52 47 4a 49 48 4f 51 50 4a 4d 4f 54 49 5c 4f 4c 55 4e 51 4d 5c 52 5c 54 4e 4f 53 58 4e 57 4f 51 4c 25 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 34 5e 69 5a 65 64 62 57 5a 5f 62 5e 5c 5c 52 58 5e 56 55 4c 5b 52 52 53 53 4e 54 53 52 52 4a 4e 51 56 51 41 58 52 4d 4f 48 41 53 48 45 49 4a 42 44 4f 46 44 4a 40 47 4a 48 45 45 4c 46 48 47 45 4b 44 3f 50 53 4a 4a 4d 51 4f 4d 4f 4e 50 4e 55 4d 57 49 4d 40 38 21 13 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 09 11 1b 2c 2e 49 47 45 51 50 4a 46 51 4e 4b 48 42 43 3f 3c 4a 47 47 44 39 3c 43 40 4b 46 48 47 40 48 4c 4b
 4d 49 46 4a 50 4b 45 4b 4a 4e 47 44 48 4a 46 52 46 49 46 4a 4c 47 42 45 4b 4b 42 45 49 50 53 4b 52 4f 4a 59 47 50 45 48 4c 49 4b 4b 4b 4c 4f 4b 57 50 51 4f 52 51 48 4c 51 4f 58 55 48 57 54 51 59 54 57 51 4c 4f 52 55 45 23 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 3c 5f 66 5c 5f 5e 5b 60 5e 57 5d 62 57 55 56 54 53 50 4f 53 5a 45 5b 4c 59 51 57 53 57 56 55 50 46 4e 52 4d 4d 4b 49 49 4b 47 47 4a 4b 51 44 4e 4b 45 4d 47 49 3b 40 52 46 47 41 4a 4b 47 41 49 47 4e 4a 44 4a 4d 44 4e 56 46 50 52 4e 53 47 52 52 57 4b 47 38 32 24 0f 04 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 11 1a 25 30 39 3a 44 4d 4c 49 4b 52 4f 48 42 49 4a 42 3a 3b 43 44 45 41 3e 43 46 41 43 47 39 3f 3e 3d 45 46 4d 46 49 44 41 42 4c 51 42 4d 45 42 4c 45 49 4b 45 4e 49 3d 4e 49 49 40 43 4a 43 43 44 49 4a 54 52 53 50 47 4f 49 44 4c 46 48 50 51 4a 4d 4b 4e 4a 56 4d 4c 50 55 4f 53 4e 51 4e 56 4d 55 57 55 4b 44 54 53 52 52 4c 3f 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 30 5b 6a 5c 60 5d 5d 54 5d 5c 60 55 52 53 4c 55 57 55 5b 4b 53 4b 54 53 50 52 4d 52 54 54 51 45 4e 46 48 4e 4b 4a 4c 56 49 4a 4d 44 48 47 42 41 46 4e 50 47 42 40 41 46 47 40 46 43 46 43 44 49 44 4d 4a 43 46 4c 4e 4f 44 4f 4b 45 53 53 4d 53 50 54 4a 40 35 25 0f 15 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 1f 28 31 32 46 46 47 49 54 55 5e 5d 4d 4d 41 4b 42 3f 41 4d 43 44 43 43 46 44 40 41 41 43 40 43 44 49 44 4d 46 40 45 49 50 4b 44 4c 3a 47 45 45 50 4a 49 48 4a 46 3d 43 47 44 42 46 45 44 40 46 4f 57 5c 59 51 4d 48 45 4d 49 45 4c 49 4d 4f 4c 42 4f 52 46 52 4f 51 4b 4b 4f 50 55 55 59 53 5a 4b 52 4a 50 4e 4c 4d 53 5a 52 49 2e 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 2c 57 5b 59 62 60 55 53 4e 59 54 4f 55 4a 4f 4c 53 54 53 50 4f 4d 5a 4b 52 4b 55 50 52 4f 5b 51 4d 52 42 4d 4f 4d 53 50 4e 47 4c 4d 48 49 49 43 46 42 49 44 48 49 45 47 3e 45 4a 41 47 42 44 4a 3f 48 43 48 46 55 48 4a 4b 51 46 55 55 51 51 47 50 4a 46 3b 2d 1f 13 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 16 1d 2e 35 45 43 4b 4d 51 59 64 61 52 4f 52 48 45 4a 3f 3d 43 41 45 41 45 3e 42 45 45 40 44 43 47 46
 4a 41 45 45 4f 46 3f 4c 45 4a 4c 48 44 4c 44 3d 48 47 47 46 49 44 49 3f 49 47 4f 42 44 49 48 55 4e 50 4e 4c 44 4c 49 44 46 44 4a 4b 4e 4d 50 4c 4d 4e 51 4a 55 4c 51 53 50 53 57 50 4d 53 52 51 4a 4f 47 53 49 5d 51 51 50 2f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 36 53 57 59 59 56 4e 54 52 58 55 54 53 54 54 55 52 4d 53 52 4f 4f 50 51 57 54 4c 58 59 57 56 53 47 42 4e 4c 50 51 48 4b 4a 47 49 4b 4f 4e 46 40 45 4a 4a 4a 4f 44 46 51 4f 4b 40 3f 45 45 44 49 43 49 45 4b 5c 4a 46 48 4f 4f 55 47 55 4e 47 55 4c 53 3f 36 1f 1b 0e 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 12 18 26 2f 3e 43 3f 51 51 50 64 67 64 54 48 4e 41 42 43 49 43 43 40 40 43 44 3f 43 3e 42 39 3d 3e 4a 41 42 44 40 47 4a 44 53 4a 4a 4d 49 43 38 4b 43 42 41 43 47 48 3c 44 44 42 46 40 43 3b 48 56 54 56 54 49 45 57 4d 4e 44 47 4e 52 51 4b 47 4d 4c 51 4f 4d 51 50 4a 51 50 4e 4d 51 48 4e 4e 53 54 53 44 4b 48 49 47 56 56 42 31 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 2c 51 58 58 5c 58 4c 58 4f 50 56 50 50 53 49 47 52 4f 50 42 58 47 53 4b 4e 4c 4c 47 52 56 4f 4d 4e 4b 48 44 50 42 42 52 43 44 4e 48 49 48 4a 4e 41 47 43 48 4c 4d 45 45 4c 48 48 3f 43 41 45 48 4c 46 45 4a 41 4d 47 4a 52 50 4c 51 4e 54 4c 4c 50 4a 3f 2d 21 1c 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 13 23 2c 45 44 44 51 46 5b 60 69 5c 4d 4b 43 49 4d 3d 42 3e 3f 46 3c 43 40 3b 42 44 41 45 46 47 42 49 44 3c 47 42 45 49 44 4e 44 43 46 40 43 44 46 4c 47 48 3c 49 3c 40 47 44 42 44 3e 4b 47 4e 4f 46 54 52 4a 4a 4e 43 41 44 47 4b 53 42 49 46 4a 47 4c 50 4d 4e 49 52 4c 44 4f 4c 4c 50 4c 4d 4e 4a 52 44 44 4f 55 4d 4b 27 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 23 48 55 5b 5a 52 50 4b 56 4d 50 4b 4f 4c 4a 4c 4f 52 4b 4e 4f 4a 48 4d 4f 48 4f 46 58 50 51 4c 46 47 45 4a 3f 41 47 48 4c 41 46 43 49 46 41 4f 40 49 4d 40 4a 42 4a 44 48 42 42 44 49 41 42 44 4b 47 4b 45 43 45 49 4e 52 53 58 48 4e 47 47 4d 46 46 32 27 1d 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 19 23 2d 40 45 45 4c 4d 55 58 67 65 54 50 52 4b 3e 47 47 3e 45 45 44 4d 42 44 46 45 3c 43 42 43
 3e 45 46 4e 4b 4b 4a 4a 49 4a 45 47 49 3f 40 44 49 4b 44 47 43 46 4d 3f 4d 43 48 44 3d 44 4a 51 51 47 4b 4d 4c 52 48 49 4f 4b 47 4f 4d 45 46 4a 4f 4b 50 4d 50 4a 55 4a 49 4c 51 4f 4e 4a 4c 44 52 50 4f 50 49 4f 4f 53 49 2f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 1a 4a 54 58 56 52 45 55 4e 57 54 4b 52 53 4d 51 50 48 52 4d 4b 4f 4b 4c 4b 4e 52 4a 4a 4b 4c 48 4d 4b 4c 46 3d 4c 42 47 4e 49 45 44 4d 48 4d 47 4b 49 43 48 4b 42 4c 44 43 49 47 4a 46 46 4a 46 49 46 49 48 4e 43 4e 53 4f 5b 57 4f 54 53 54 4e 43 43 34 21 1f 0a 09 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 1a 22 2e 34 3c 45 4b 4b 56 5c 5e 5c 54 54 49 41 47 44 45 47 44 3e 3f 44 41 46 43 47 41 48 45 44 43 47 3a 46 44 49 45 48 49 44 3f 3e 3e 49 41 45 44 41 44 44 45 44 44 44 45 46 4d 45 3b 3a 48 4c 45 4a 4d 49 4d 48 52 49 4e 4e 49 4a 45 4b 4d 49 4d 49 4b 4c 4b 4f 49 48 46 4f 4f 4c 46 53 4c 4f 4c 4d 44 49 44 4c 4a 52 48 2d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 4a 5b 53 59 55 53 53 4f 4c 49 49 52 47 48 52 51 4d 49 46 50 47 4e 4d 45 4d 49 48 4a 49 44 46 46 45 49 4a 4b 44 44 49 49 43 44 47 45 4a 4d 44 4c 3e 43 43 49 44 4f 40 46 46 43 45 44 4a 4c 49 46 48 4c 4a 48 50 55 54 56 5b 60 57 52 53 49 4f 44 35 2a 19 0f 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 13 2c 2f 3b 3c 41 4b 56 5d 5e 60 51 49 50 43 42 4d 48 46 40 43 3a 3a 48 47 3c 4a 42 44 42 45 45 42 3a 41 45 47 3a 49 42 57 3f 40 47 4f 42 3f 3b 43 3f 47 47 3d 42 40 44 46 4b 34 42 41 49 4d 44 45 44 52 45 46 47 4c 53 4c 48 4f 4a 50 42 4e 4d 47 49 4f 40 4d 45 49 4c 4a 49 4d 4c 45 4d 4b 4b 4d 46 46 45 47 54 4e 41 30 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 47 53 45 57 4c 48 50 50 4b 4d 42 47 4b 4c 4f 49 4f 50 4c 45 40 4b 45 4e 53 50 52 4c 50 44 52 42 49 4c 48 4a 46 46 44 45 4c 4b 39 3b 41 3c 48 3d 4a 47 44 49 4d 48 42 3f 3b 45 41 47 4a 46 49 48 48 4d 45 48 4d 4a 58 5d 5c 61 4f 56 51 49 45 38 37 2d 12 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 1d 1d 28 33 43 43 4f 56 5a 5f 5a 4f 54 50 4d 4c 4f 47 4a 4a 42 45 44 43 42 43 48 3a 3b 3d 45
 40 47 44 44 45 47 46 54 46 43 4c 48 3f 43 44 48 44 47 3e 4c 45 4a 42 3b 45 42 42 45 42 45 4a 4d 4b 48 3f 49 3f 4a 4f 4b 4d 46 4b 49 44 4a 45 4b 48 4b 4d 4f 44 51 48 44 47 44 4f 47 4d 43 4a 45 47 47 4e 46 52 4b 49 4e 46 36 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 23 3d 4b 4b 51 4f 48 4a 4a 4a 4f 46 46 47 4b 4c 47 41 4c 4a 51 45 49 4a 49 4b 53 50 4d 4b 48 48 47 45 47 45 45 45 4b 44 44 47 49 44 43 4b 41 41 39 48 41 3e 40 40 4a 4a 46 4c 48 45 47 4b 44 45 4f 4d 50 49 4d 51 56 55 5b 5d 5a 54 57 47 45 44 34 29 24 13 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 14 13 26 34 39 3a 4a 5d 59 56 5b 52 49 47 52 5c 50 54 4f 42 41 3e 47 44 4b 41 43 3e 3e 45 3f 42 49 46 44 44 3f 41 50 46 4b 45 49 42 45 48 41 48 42 3f 42 3f 47 44 45 45 3e 3d 49 49 45 4b 45 4c 4d 48 4c 4c 41 45 48 4f 49 4b 4d 3f 49 44 44 4e 48 49 49 3b 49 49 4c 3c 48 4d 47 4a 44 44 46 40 4b 47 45 44 47 4e 4d 44 36 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 37 4e 4b 52 4c 46 44 4e 41 4d 49 4b 48 47 50 4b 4a 4d 4d 4a 43 4a 4b 50 50 4e 4d 4f 4a 44 43 46 47 48 46 43 41 42 43 45 43 45 40 3e 4c 47 45 42 46 40 41 44 42 42 4d 45 44 44 46 4a 41 4c 4c 49 4f 4b 51 50 56 58 5a 64 5d 5c 4b 49 4a 44 39 38 2b 22 06 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0b 1a 1d 2b 38 3b 4c 4d 4e 55 54 50 50 44 4e 49 51 55 46 52 49 47 3e 40 3f 3d 44 3c 41 3f 45 3c 4d 3e 46 3e 3d 41 44 44 44 4b 40 44 3f 38 4c 40 44 45 48 3d 45 43 47 46 44 3a 4b 3d 3f 42 48 46 45 4f 4a 51 41 45 4a 47 49 42 41 40 44 47 44 4e 43 49 44 40 47 40 41 43 46 4c 4a 46 3e 41 48 46 48 45 44 45 44 52 41 44 38 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 30 54 45 4c 45 42 47 45 47 49 49 42 48 43 45 48 44 51 4b 4b 4a 47 52 47 4b 4b 4d 4e 4b 42 44 42 43 50 48 42 49 4d 3d 41 48 48 43 44 45 41 41 3f 4a 45 40 42 40 47 43 46 4f 4a 45 48 57 4b 51 50 52 54 48 51 54 54 5d 58 4a 55 42 45 4b 44 3c 30 22 1d 0f 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 15 20 2a 37 35 42 4c 49 52 4b 4b 4f 48 54 46 55 54 4c 4e 4b 41 3e 4c 42 3c 40 3e 4c 45 4c
 3b 42 42 45 4a 46 40 49 4d 49 4d 46 45 47 47 45 46 40 41 44 49 44 41 4c 4b 43 44 3f 46 47 4c 40 4a 4b 45 4c 41 45 49 4a 4e 44 44 3f 47 44 43 46 4d 4a 49 45 42 4d 4c 42 45 4d 48 45 44 4c 4e 4c 40 44 46 44 47 46 4a 4b 48 36 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 37 46 49 4e 4d 4a 47 46 4d 4a 50 49 43 4d 42 48 46 49 47 4c 4a 52 49 4a 46 46 51 4e 42 47 46 3f 47 4c 45 3d 45 47 50 4a 48 45 43 42 4a 4e 45 44 3d 44 44 43 41 4b 48 46 4c 43 45 51 52 48 4f 5c 50 5b 58 5e 59 59 5a 5d 4f 54 4a 48 4b 3f 3b 30 23 1b 09 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 1b 22 33 3c 3b 41 44 47 48 49 46 3b 43 4e 53 51 4e 40 48 44 4a 41 4f 43 47 45 46 47 3e 44 45 40 45 4b 43 40 47 42 43 42 48 46 3d 44 45 43 40 4a 3e 40 46 49 47 47 46 44 44 42 41 4a 4a 51 4b 43 41 45 47 4d 46 4a 44 49 47 45 46 44 42 4a 3f 46 4f 46 45 44 46 43 46 48 4f 45 49 48 44 49 3f 3e 41 43 3e 41 4d 3d 31 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 32 47 4a 4a 51 42 46 47 3f 53 49 45 42 4e 47 49 47 47 4a 4d 46 46 48 4e 45 42 4c 4b 45 48 41 47 46 4d 47 46 3c 4b 49 3d 41 47 44 3a 3f 43 3f 3e 4b 49 46 40 43 49 43 44 52 4b 46 49 5a 57 5a 55 5b 60 4c 56 52 54 57 5c 52 54 44 47 39 35 3b 21 17 0c 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 12 13 25 31 3d 3c 3a 42 47 47 41 4d 4e 56 51 58 50 45 46 4f 53 49 45 4b 4c 40 43 41 3c 42 40 42 46 3f 40 4c 42 4d 48 43 43 46 46 41 45 46 46 45 42 3a 49 4a 45 50 4c 42 44 46 49 4c 53 51 40 45 4a 4a 3e 43 43 3f 49 49 44 46 45 39 46 4b 45 47 44 47 46 45 4b 3f 47 3f 44 44 45 40 43 3e 44 43 42 44 43 42 46 37 2e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 2e 3d 48 4a 48 45 46 42 4c 41 49 4d 4a 46 47 44 49 43 4d 45 49 50 4c 4f 46 49 49 3a 47 44 3b 3f 41 3f 3b 41 3f 3f 42 3f 42 41 43 47 44 38 45 47 47 3d 45 4b 3e 54 4e 4e 51 5b 5a 5b 5e 57 5e 58 5b 56 4b 51 54 55 4f 4e 49 48 4a 3e 42 35 2c 20 15 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 13 2a 2c 37 40 37 3b 44 3f 48 46 4b 58 5a 58 46 48 47 4b 54 57 4f 4c 4c 50 45 4a 49
 3e 49 4f 3c 45 41 47 4a 4a 42 4a 4a 4b 46 41 43 44 46 44 47 3e 42 48 41 49 44 45 43 47 46 55 3e 26 35 51 4e 46 41 3e 44 47 4a 46 40 3c 3e 3e 44 4b 44 4c 43 3e 41 44 40 49 43 41 43 48 4c 3b 40 48 41 45 44 3d 49 3a 49 3e 30 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 33 4a 4a 46 4c 43 43 45 41 4a 42 4a 52 4c 3e 4d 50 45 46 4b 49 4a 43 48 4c 43 42 45 3d 3e 44 3e 48 40 3d 36 38 44 48 3d 3c 48 3f 42 48 45 47 49 47 45 45 44 48 53 4b 52 58 61 66 5f 61 59 53 51 5b 54 52 54 54 5a 4f 44 4a 46 43 43 3e 32 2a 1b 13 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0e 1e 28 32 3b 41 3d 45 3c 41 48 48 4f 5d 5d 5c 50 4e 4d 4f 53 53 4b 4d 51 4b 4a 43 43 46 46 49 49 48 48 4a 46 48 4e 45 4f 47 3c 45 47 3c 47 42 49 4b 44 3e 4c 43 43 4e 44 4f 4c 49 4f 4f 51 45 42 47 45 46 49 43 42 45 41 42 42 3d 3e 3e 40 47 4b 4a 47 4f 43 48 48 46 3d 46 43 45 42 43 45 45 3e 41 43 3f 42 30 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 2a 44 43 4b 4b 3a 48 45 40 4b 47 50 51 47 49 42 42 3e 43 49 4c 44 49 4c 49 41 41 47 4d 46 3a 43 47 43 41 41 49 4a 44 44 44 3e 3b 49 48 45 41 46 3e 53 44 47 53 60 51 5d 63 66 6c 61 65 5a 4f 50 4d 5b 4a 57 48 58 4b 4b 51 49 43 43 3e 28 23 19 10 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 19 23 2d 3e 41 3e 45 44 39 42 44 4a 4f 5f 60 54 46 4b 46 4f 41 50 55 52 56 49 47 43 41 43 42 46 4f 43 45 49 44 40 3e 48 4d 42 44 47 45 45 40 44 49 41 46 49 4b 43 4c 48 45 56 4e 49 42 44 4b 3c 44 45 3b 49 47 46 47 3d 45 40 45 49 43 42 40 45 47 3f 48 3e 40 42 3e 43 48 39 44 44 42 45 3e 37 41 3a 3d 37 2c 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 29 4e 43 49 43 46 41 46 3f 49 41 4a 46 47 47 46 47 44 41 4a 3d 47 49 46 45 43 38 41 3e 41 41 3d 45 3b 40 3d 3e 3b 44 49 3c 44 37 44 48 49 46 47 4a 4c 49 4e 55 64 5a 60 5f 63 5c 64 4f 54 44 4f 52 4b 52 59 55 50 4a 4d 49 46 3c 3a 30 26 1d 0c 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 12 17 27 35 38 40 3e 3d 3b 43 3f 47 43 4f 4c 48 49 48 4d 46 4e 4e 52 5a 50 56 4d
 41 46 4f 43 4d 44 48 44 43 48 43 43 3e 4a 49 47 40 42 43 4c 3b 42 3a 41 46 4f 43 41 4c 45 4b 4e 4b 45 44 4a 42 41 41 44 3e 45 4d 49 43 41 39 3f 44 49 45 46 41 47 3f 45 46 3e 42 47 45 41 45 3d 3e 3b 35 42 41 38 4e 3b 3a 38 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 28 43 40 4a 48 49 45 44 3d 3e 47 4a 48 44 46 47 46 3f 3f 3e 39 40 41 41 3b 41 42 45 42 40 3f 42 42 3e 39 3b 3f 3d 35 44 44 43 40 45 41 43 49 52 49 4d 5a 5e 68 63 65 64 61 5d 52 4b 4f 4e 47 4b 51 52 4d 5b 51 4c 4a 4c 4b 4a 42 30 2c 1c 1b 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0f 16 1e 30 34 3e 3b 3f 46 3e 3a 44 42 44 45 44 4a 43 48 3e 49 49 4f 59 55 57 50 4c 46 4e 48 49 45 4a 4d 49 45 44 4a 45 46 43 48 43 4a 40 44 45 42 44 46 47 3d 4a 4f 4c 4d 4e 4b 4c 49 53 4b 42 4d 45 4f 52 43 48 45 42 41 4b 3f 39 3a 45 48 4c 4a 47 44 45 40 41 44 38 3d 42 41 3f 42 39 42 42 3d 3f 44 38 32 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 1c 42 44 4b 40 4c 43 44 42 53 43 40 45 46 3d 41 3e 40 43 47 45 48 3c 43 48 42 45 40 3d 40 41 42 3d 3f 3e 36 40 3e 3d 48 3e 3f 43 4b 42 4b 53 4e 5b 53 54 64 66 67 59 5b 56 52 4c 4d 4e 48 4e 4e 55 55 50 57 49 4e 47 4c 42 41 39 38 2b 23 18 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 0f 19 27 2b 2c 3c 33 3e 48 42 47 41 49 3e 47 3f 43 3e 43 40 47 4d 4f 55 4f 59 55 4c 48 4b 48 4b 4c 4b 41 49 4b 45 44 46 41 41 48 3f 4d 47 45 49 47 44 46 4d 51 58 47 42 4a 45 4b 4a 47 46 43 44 44 45 52 42 3d 42 40 49 45 46 40 45 47 40 3c 3b 3e 3a 3e 40 45 4c 44 44 38 42 41 3e 35 43 44 42 49 42 37 2f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 3e 44 4d 41 40 42 3e 40 41 41 41 3b 46 3b 3e 40 45 42 46 41 3f 38 43 36 44 49 42 46 43 38 45 3d 37 40 3e 43 44 42 42 3e 49 4d 4a 54 53 4b 4f 51 56 4f 5b 5b 61 55 4f 4e 47 47 4c 47 47 46 47 4a 56 4e 4d 4e 44 4e 48 40 44 32 2f 22 1e 14 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 17 1f 25 35 41 38 44 3b 3f 41 41 41 44 42 38 44 3d 4b 3d 3f 44 47 49 4d 52
 56 5b 59 44 4e 48 47 45 48 46 47 45 3f 43 41 44 53 45 41 4b 45 46 4c 46 52 44 45 4c 4c 47 47 45 4f 42 45 4a 4b 41 47 4c 4a 40 4b 3d 3c 45 3b 46 40 3c 43 47 4a 40 42 41 47 3c 3b 40 41 41 37 42 40 45 43 3c 37 33 3a 3a 39 2e 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 44 3a 4c 4b 45 3d 41 42 41 48 41 41 3f 3e 49 3c 43 40 3f 40 41 40 40 43 3a 45 3d 36 3c 3d 44 47 41 34 3c 4a 3b 41 42 3b 4c 4d 45 54 4a 54 50 50 53 4b 5c 58 56 51 4f 52 49 47 49 44 45 48 4f 40 4b 49 4a 49 43 41 42 4a 41 34 26 22 12 0a 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 1a 28 28 33 3d 48 3a 43 3f 4b 39 3c 43 3b 43 43 4b 47 45 45 45 47 4d 52 64 69 60 5b 4e 4c 49 47 44 45 49 41 41 4a 42 45 43 40 47 4d 45 4f 52 4a 4b 4a 4d 4b 50 46 47 43 47 41 42 46 46 45 44 47 47 42 45 48 43 43 41 4a 43 48 3f 45 3e 4e 42 40 3c 44 42 43 44 42 40 43 3b 38 3b 42 47 3d 3e 3d 30 2f 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 1a 3c 3b 3d 3d 3d 43 44 44 3b 3e 46 40 44 3b 4a 45 4f 3a 3a 43 41 3d 43 42 45 41 3a 41 41 40 43 3e 47 3b 47 3b 45 47 44 49 4b 59 51 4c 4e 52 48 4d 45 48 53 48 55 4f 49 59 49 3f 43 44 54 50 50 4a 47 42 4c 45 45 48 40 3e 3d 2f 25 25 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 17 1c 23 35 3b 3e 3e 38 46 46 42 43 3b 46 43 45 46 41 49 44 43 46 53 50 5d 71 68 60 55 4f 47 47 4c 47 46 4c 4c 49 41 49 44 3d 42 42 3e 49 47 4d 4a 4a 53 4e 4a 4a 41 45 4b 4b 4c 4d 4f 44 42 44 43 40 4c 41 44 3e 3f 42 3e 44 45 44 40 45 3c 43 3f 3f 3f 42 40 3e 41 43 40 3f 3e 38 3b 40 45 41 39 32 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 40 3e 41 41 3f 45 3a 3d 40 3c 46 42 45 3b 46 43 46 41 39 43 3f 3e 3b 3b 45 36 47 3e 45 41 44 44 40 42 41 36 3e 3f 44 48 50 4a 44 52 49 48 4b 45 41 48 4a 4b 4a 4a 41 3f 49 47 54 44 49 4a 49 43 50 44 3d 40 42 4e 3d 3e 3f 2b 1b 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 0f 1a 18 2b 33 3c 40 42 39 49 3d 42 3f 47 45 40 49 42 49 47 46 45 44 51
 64 69 67 60 50 55 49 49 43 42 49 4b 3e 40 46 4e 42 47 45 4c 3f 49 4a 49 4d 49 4b 4f 4b 45 44 44 43 46 44 48 43 41 45 45 41 3f 47 43 3e 3e 3e 44 42 3d 42 41 3d 42 49 40 40 41 44 46 43 47 35 40 3b 42 42 3d 37 40 38 3e 3b 2a 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 37 3d 3c 3e 3d 39 44 37 49 34 3f 41 40 41 3c 40 3c 3c 44 3e 3c 40 41 3a 39 37 39 44 3b 3b 3d 3e 39 42 3a 3c 42 3f 3e 42 47 49 44 45 44 41 3c 39 3b 3a 49 45 48 51 4a 49 4c 41 43 3f 44 47 4e 48 48 48 44 3f 4a 48 3c 3b 2a 24 1d 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 10 19 23 35 38 3e 43 42 45 3e 43 45 47 45 46 41 3e 47 45 43 44 47 55 53 5c 62 59 4e 50 49 45 47 4e 48 3e 3b 48 4b 49 4a 40 45 4f 46 41 4f 45 48 4f 4c 4e 47 46 43 4d 48 47 40 3f 46 45 43 46 47 41 44 40 3d 46 35 44 41 3a 3d 44 44 46 45 3f 39 41 3b 45 42 46 47 43 41 44 3e 41 3d 41 3e 39 34 32 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 16 3e 39 39 3e 38 3c 3f 3c 3c 39 41 39 41 40 3f 47 39 3e 44 42 47 40 4f 37 3c 3c 40 44 43 3d 3c 40 37 3c 41 45 46 46 4b 3d 48 44 46 49 44 40 46 45 49 43 42 41 4d 4c 3f 46 46 41 4b 44 49 4c 4e 47 50 45 42 49 3d 35 3f 36 34 1d 1a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 10 22 21 33 36 41 3c 3b 45 45 40 41 47 47 3f 47 45 44 44 40 40 4e 56 60 56 56 53 50 49 45 45 4a 42 49 49 49 4a 4a 4a 46 47 4a 42 4b 4d 45 4c 49 47 4c 4a 4f 4e 47 45 48 47 3e 41 3f 42 47 45 3c 43 45 41 48 37 42 41 3c 3d 42 34 46 3e 45 3c 43 45 44 49 3f 3b 35 3c 39 3d 3e 3e 41 3a 3f 3c 35 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 11 36 3b 3b 42 3f 37 3a 34 3d 39 3e 43 3f 3e 3c 41 47 3e 3e 45 41 3d 48 3e 40 3c 45 3b 44 38 43 44 3b 41 3f 3e 46 44 49 4b 43 43 3f 46 43 39 41 42 43 44 42 43 3f 49 47 47 45 40 4f 4b 45 4c 4a 40 4a 45 48 41 47 3d 35 36 2a 17 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 12 1d 24 28 36 39 3d 3f 3f 44 37 3e 3d 44 41 3f 41 48 47 43 45 42
 40 51 4e 51 4c 4b 47 46 46 4e 45 44 46 47 44 44 41 40 4c 4d 45 49 4a 45 42 48 3e 46 40 48 41 44 44 41 41 44 40 47 41 48 40 3d 40 42 3c 40 3d 40 3d 39 3e 3a 3f 3f 3a 3b 41 44 49 41 41 45 45 3a 3f 34 45 35 37 3b 3b 34 32 31 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 32 3e 39 3e 3b 36 3d 3c 44 41 3b 44 44 40 3e 3e 3a 3e 40 3c 41 42 35 45 3d 3e 39 41 40 42 46 44 3e 3c 45 3e 44 42 46 45 40 3e 37 4d 3f 3b 41 44 3c 41 41 48 4c 47 44 3e 42 3e 49 47 45 46 42 44 3b 43 42 3e 38 2e 28 27 12 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 0c 1f 22 35 2f 39 3f 42 41 49 3e 40 45 44 43 4a 49 40 40 41 39 44 4b 48 49 48 49 48 3e 48 3f 42 42 41 46 44 40 43 44 4b 47 4a 46 48 44 47 46 4b 45 44 46 4a 40 48 4a 48 49 3a 43 44 45 45 44 49 43 3a 3f 47 40 49 3a 41 43 43 40 40 3a 43 51 4e 4b 4b 42 3e 42 38 34 41 3b 3e 42 3c 3a 2f 33 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 33 35 39 4a 3d 3f 41 43 3e 42 3b 3c 45 3d 3e 3e 3f 3c 3e 35 3c 3a 3b 42 35 41 3e 4a 47 3c 42 3e 49 3b 3b 41 3d 43 3e 47 47 4a 45 40 41 41 3f 3e 3f 3f 4b 45 49 43 3e 48 41 40 48 44 43 4c 4f 47 49 40 43 45 3c 36 33 22 21 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 19 23 29 42 3b 43 44 3c 3c 42 41 4a 40 42 4c 43 4a 4b 3d 42 40 4b 44 52 49 47 44 45 48 4f 3e 44 40 45 4a 4c 48 46 48 42 41 4c 44 45 49 47 4e 44 44 3f 45 50 45 49 52 45 4a 41 3f 41 43 4e 43 4a 3b 3c 42 3c 40 48 3e 44 47 52 4d 4a 4a 46 54 4a 45 47 3e 46 3f 3f 3c 38 38 3e 36 3d 2d 31 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 10 30 37 3f 3b 40 41 43 40 3b 35 44 39 43 3f 47 44 44 3d 41 3b 41 39 45 3f 41 45 46 45 40 45 47 3c 42 40 42 49 3f 3c 44 3e 40 3f 3c 40 43 41 3e 3e 43 3a 42 49 43 40 3d 44 44 47 4e 47 44 44 54 4d 49 46 46 3d 38 30 27 18 0f 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 10 1a 2b 2b 29 33 34 40 39 40 3a 3e 46 40 46 3e 44 3e 3b 41 41
 48 41 4d 49 4b 4d 40 44 40 3d 49 4c 45 43 41 43 52 40 4d 45 48 3e 41 48 45 49 4b 44 41 43 45 45 4a 44 4c 4b 43 41 3f 42 46 4f 50 48 41 3a 3b 3b 3b 39 43 42 45 50 46 45 45 4a 42 54 4b 45 3c 3c 3d 3e 3c 3b 3f 38 34 3b 3c 33 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 36 44 45 3f 44 44 43 39 45 43 37 42 3e 43 45 3a 3c 39 42 43 3f 46 49 42 3d 41 45 42 45 39 34 3f 40 3f 39 43 44 45 37 42 41 3a 42 43 3d 40 48 3a 3f 41 40 3a 47 3f 4b 47 41 49 4b 44 44 3c 44 48 46 44 4b 47 3e 2e 24 0d 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0e 18 24 26 35 43 3f 40 38 41 44 45 3f 44 49 44 4c 48 40 3d 43 3e 49 47 42 42 46 40 41 4f 49 41 49 4c 47 47 47 49 49 44 3f 4e 48 47 49 41 4a 4d 42 49 4f 47 50 4d 50 4b 47 40 4a 4c 44 49 4e 43 46 44 3e 44 3e 44 46 3e 45 4b 41 44 49 4c 49 51 4e 4d 4d 3f 42 3c 38 35 34 3b 42 39 35 2b 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 27 34 46 44 42 46 47 4a 4c 4b 4c 3c 44 43 3f 44 41 43 49 41 45 46 4c 45 41 42 4a 44 3d 37 41 3f 39 44 3f 4b 47 45 48 3c 40 44 3d 41 47 42 43 43 3e 42 48 44 49 41 3b 4e 4b 49 43 40 43 51 47 46 46 4a 48 40 37 24 1d 11 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0c 12 1c 22 2e 38 34 37 37 3d 3d 3d 47 47 40 42 41 44 43 40 44 45 40 47 41 48 3f 45 43 50 50 47 4c 50 45 53 44 42 43 50 3d 3e 50 47 4b 54 40 50 48 46 41 48 53 4a 53 4b 3f 41 3c 44 4b 4b 4a 44 3c 3e 3b 44 3d 3e 43 37 41 43 3e 38 40 42 47 54 48 58 4e 41 3c 37 39 32 35 30 3e 37 37 29 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 3a 44 55 52 59 5a 5a 54 4c 4a 46 49 46 44 43 4b 43 4d 45 47 46 47 47 41 4a 4a 45 48 3f 40 49 44 3e 3a 44 42 41 43 40 3d 4c 49 48 47 41 3d 45 46 35 4b 44 45 49 40 43 49 44 44 46 45 48 46 4a 48 4a 3e 35 28 1c 14 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 10 25 34 2c 3e 39 42 3a 38 41 3c 41 3b 3a 3b 42 45 43
 47 3d 3e 3f 48 46 42 3d 47 4b 4d 4e 4d 51 54 50 4d 49 47 47 3e 52 49 4a 47 49 4d 46 47 45 4f 47 41 49 45 42 49 3e 3d 44 42 46 43 48 3e 38 40 42 40 36 3a 3b 36 39 39 3c 3c 39 3f 46 47 4e 45 40 3d 3a 3d 40 41 39 3e 37 31 30 21 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 32 3f 4a 62 59 5f 67 5b 58 55 4b 4f 48 49 4e 4f 50 41 46 4b 4f 40 4e 47 44 48 45 47 47 44 46 48 4c 4d 49 4c 51 49 51 4e 4c 47 50 54 4e 50 44 43 47 41 42 49 46 48 3f 4a 42 3f 49 46 41 43 44 50 48 3f 39 30 1b 18 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0b 1d 28 38 36 3c 35 3b 3b 3f 3f 42 42 45 44 41 3b 41 45 46 42 38 3d 41 3f 43 44 48 4e 47 51 4f 56 57 50 4e 41 50 45 52 4c 46 47 47 40 45 41 45 3d 48 47 41 45 3e 41 41 41 42 40 36 47 37 43 42 3e 3e 3d 3a 35 3a 3a 31 38 37 3f 3e 3e 43 40 41 44 3c 3f 3f 52 4e 45 3b 3c 36 38 2b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 08 34 3a 48 54 5b 5f 5b 56 5c 4d 4a 41 48 49 4d 44 4d 4d 52 4b 51 4d 52 52 58 59 5c 5a 61 59 59 65 61 62 5c 61 5c 59 5a 58 5c 53 52 57 52 57 4b 48 4a 43 3e 41 44 45 41 49 42 42 47 44 42 4e 4b 47 42 3d 32 2c 14 09 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0d 18 21 28 34 36 37 39 3e 3b 3f 41 47 41 3e 42 49 44 41 3f 48 46 3f 3d 3f 3f 42 46 49 4c 55 51 55 56 59 4d 4b 47 4c 4b 4f 4c 4b 50 45 48 43 41 43 45 49 3e 3d 42 41 39 3a 3d 41 43 3e 3c 43 37 34 3d 3c 3f 36 3a 3b 38 30 34 3d 3a 3d 40 3a 41 3c 39 3f 46 43 44 3c 3e 35 39 3a 32 2a 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 3d 46 49 49 51 57 4c 4f 45 41 4b 4e 56 4c 56 58 53 56 58 66 6a 6c 6a 67 6c 6f 73 75 71 6f 7d 76 6e 75 70 76 77 72 75 6b 65 6d 63 6b 5e 5a 49 48 40 44 49 49 4a 4f 42 44 42 48 45 4b 3e 45 3f 3d 34 33 1e 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 08 10 21 1c 2a 37 33 39 38 38 3c 4a 44 3e 48 3f 3f 47
 49 41 44 46 3d 40 44 3e 46 4a 4b 4c 52 50 52 57 57 4e 47 4c 4b 4e 46 46 56 4c 4c 42 3a 46 41 41 42 41 3a 3c 37 3d 36 3c 43 33 33 34 34 34 35 3c 32 3d 38 34 3f 31 3c 43 39 3b 36 3b 40 3e 39 38 3b 44 44 46 44 36 41 38 31 31 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2d 46 48 51 4b 45 4f 49 4e 45 4a 4e 52 5c 59 67 64 6c 73 71 75 78 80 81 79 83 7d 7f 7f 7a 7b 7a 7e 85 88 7f 84 81 78 7d 7a 7c 7b 77 76 69 68 56 49 42 45 3c 46 41 3e 42 3d 42 41 44 3e 3f 3b 34 2d 26 18 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 0e 1e 2c 2e 30 31 36 3d 42 3f 3a 4a 37 39 46 37 45 42 3d 3e 45 3b 42 44 3e 46 46 51 48 57 55 55 49 4c 4f 44 46 48 4c 49 4c 48 3a 41 3b 3f 3f 41 3f 3a 3c 3d 39 38 39 39 3b 34 40 3b 38 42 35 3a 33 31 30 35 37 39 37 37 3b 34 3c 3d 34 36 39 33 3d 33 3b 35 3a 39 36 34 2b 34 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 24 3c 41 49 48 47 49 52 4d 59 5b 69 66 67 70 72 7b 83 86 7f 82 85 88 83 83 87 8f 87 81 88 83 8d 86 87 81 86 8c 88 87 8c 88 83 78 7a 74 6e 71 65 57 4b 45 3f 4b 3e 43 3e 3f 3f 44 40 3f 40 3e 32 2d 15 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 14 26 2b 31 32 3d 3b 39 41 40 46 44 44 3e 43 41 46 45 44 43 44 44 43 41 47 4d 4e 48 5a 4d 52 4c 43 4e 47 40 48 45 43 4a 3f 42 4a 36 3f 41 3d 41 43 3e 35 39 31 40 3b 3a 3a 3b 35 2d 3e 3c 38 3f 3a 34 3c 2d 38 3b 31 36 3b 42 37 36 3f 3a 39 39 3e 3e 3d 39 31 37 37 32 36 27 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 2c 36 43 49 47 52 52 67 6b 6d 6f 6d 72 80 7a 86 89 84 85 82 84 8a 90 91 89 8b 8a 8a 88 8c 85 87 84 85 88 90 8c 91 85 81 84 81 80 82 7a 72 70 69 50 4d 43 41 43 40 40 41 46 40 47 41 3f 3d 40 35 27 13 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 12 1e 25 2a 2f 34 33 46 37 38 40 3c 34 39 46
 40 47 38 3d 3c 44 39 44 45 3f 47 46 4b 4f 4d 42 42 47 3c 41 45 44 45 40 3f 3c 38 3f 3e 3e 3f 40 35 3f 3e 3c 34 3a 3c 37 3b 31 3b 32 35 39 35 35 38 35 33 3a 36 38 37 32 39 32 39 31 2f 38 37 3a 39 34 30 38 35 2f 36 32 30 2b 26 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 32 3f 4c 52 56 65 69 72 6e 7b 7d 7d 84 87 8d 84 83 85 89 88 8d 95 82 8a 89 92 89 86 8b 82 8b 88 80 84 8f 86 8e 88 84 84 8b 7f 7c 7b 7e 73 70 5e 57 47 3c 3f 3e 47 43 46 3a 3f 45 40 38 40 2f 27 18 13 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 13 20 23 30 2c 33 40 39 37 3c 38 44 3d 38 43 43 43 43 3e 47 3c 41 43 41 3f 42 45 48 41 3e 3c 3b 39 43 42 40 45 33 3d 3c 3d 3c 3b 3a 39 40 3d 39 40 3d 35 39 40 36 3a 3d 41 3a 36 33 39 39 30 32 34 39 38 3b 3a 32 3a 32 37 39 3c 2f 35 35 35 32 32 28 32 27 30 34 35 2c 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2e 4b 5d 6a 6a 6a 77 85 81 87 81 80 89 81 8f 83 88 86 86 8d 8b 8b 8e 80 87 86 81 7e 87 89 87 81 83 88 87 85 82 84 84 7f 82 7c 77 79 71 6e 64 5d 54 43 3e 39 42 43 46 43 40 3a 36 42 39 34 33 1d 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 10 17 17 29 33 2f 36 3d 3b 41 3a 3b 42 3f 4a 47 42 40 3f 47 46 45 3f 44 3e 44 41 4c 42 3d 43 3a 42 40 3c 40 3e 3e 42 49 37 40 40 38 3f 3b 3a 36 37 3f 36 34 38 39 3a 39 32 32 41 36 3a 3e 3f 34 37 35 38 39 38 32 36 2f 43 3c 3c 33 31 34 2d 35 33 2f 2b 30 33 2c 2a 2a 21 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 34 55 6a 77 73 7b 83 81 88 87 89 91 86 88 89 82 88 87 85 8e 85 8d 8a 82 86 8e 8a 8e 8c 89 7f 88 89 86 7f 7f 7e 84 82 7c 7c 79 74 7a 6d 68 5d 57 48 45 3c 3c 44 46 3e 43 3f 3f 43 3e 39 38 2d 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 15 1a 25 32 37 3a 39 3b 39 40 44 39 4a
 45 4b 3b 3c 3b 4c 42 49 43 49 38 41 3b 46 4a 3d 44 43 40 4b 45 3b 3f 41 43 3a 3f 3f 39 42 3b 46 49 3c 42 40 36 47 3d 3e 3e 3b 34 3e 42 3b 2f 32 39 35 39 37 35 36 34 2b 3c 2e 32 35 37 3d 38 32 2a 33 32 34 32 2e 2b 28 30 2d 1f 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 40 67 7c 87 8a 88 84 89 8c 87 87 85 84 89 8b 87 92 84 8e 85 83 7d 89 7c 7c 84 80 85 7f 82 84 87 84 83 7f 7e 83 75 79 7f 57 7e 75 68 6d 5b 50 4a 4b 42 44 42 42 3e 42 43 41 36 3a 36 31 2f 20 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 12 1c 23 2d 2a 36 39 3e 3c 37 3a 3e 45 3c 3a 41 3d 43 3e 3b 42 43 42 48 40 3e 43 3f 47 47 40 43 47 40 42 34 3e 3c 42 43 3a 3d 3d 3a 3d 3b 3b 43 3e 37 35 3a 3a 3d 36 38 3c 35 33 3c 3d 39 2e 37 30 33 35 2a 33 3b 39 3b 35 2f 31 33 31 2d 31 31 32 29 28 27 28 2d 22 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 37 6d 80 8b 7f 83 84 89 8a 85 86 88 8b 8a 85 85 7d 7f 84 83 80 81 82 80 83 75 80 81 84 7a 7c 83 77 7c 85 77 78 7e 75 7a 7c 68 69 65 5d 4d 50 41 42 44 42 3d 45 44 41 45 46 3d 3a 34 28 1b 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0b 21 26 38 39 35 36 3d 37 40 3e 3b 3f 43 3e 3d 4c 40 45 3f 46 44 43 3b 44 3d 43 48 49 41 3f 40 47 43 3f 3b 3d 3f 38 3e 41 45 3a 3c 3c 3c 40 3c 3b 40 3a 39 3b 31 40 3d 34 32 36 3b 33 36 37 38 37 33 37 2f 33 33 32 2d 35 33 34 2d 2b 2b 37 2a 2a 36 35 2f 26 24 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3f 76 7c 8f 81 8c 81 7d 89 84 86 88 83 84 7e 84 83 7e 84 7a 84 79 81 76 79 79 7f 79 80 83 7e 81 79 76 79 7a 72 75 6a 73 6c 62 67 5e 62 57 45 4a 41 40 4a 40 41 3e 37 38 3b 39 30 27 1f 19 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0f 1a 2c 2e 37 38 41 42 3a 41 3b
 3c 42 40 3b 3c 45 3c 40 3f 44 42 47 46 3e 3d 3f 44 41 3e 45 3a 40 44 3f 46 3a 3b 3c 3e 44 48 44 3d 3e 3e 46 39 3a 35 3e 38 34 39 3e 40 41 31 38 38 37 31 3a 3b 33 38 39 34 2f 3e 2f 36 37 35 2e 30 31 29 2d 27 35 2e 30 21 2e 24 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 44 79 80 8e 80 7f 84 80 81 83 85 7c 7e 7d 7d 7f 82 7b 7d 77 7e 79 7a 7c 6d 7a 81 7e 7b 78 7b 7a 71 7b 78 74 6f 6a 6e 68 70 64 64 5c 4d 4f 4a 42 41 3f 42 3f 3c 45 36 36 35 30 31 27 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 16 26 28 3c 35 37 39 37 36 3f 3b 44 3a 41 3e 37 43 48 43 3e 48 3a 3b 3f 40 3b 3f 40 4b 39 3e 43 36 3e 3a 3c 37 3c 36 39 43 46 3a 39 41 39 34 3c 39 3a 31 41 38 37 3d 32 3f 39 38 2e 31 35 36 36 35 3b 33 35 35 34 34 33 3e 32 31 28 31 30 2f 2f 33 2b 27 27 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 71 84 8c 87 79 7f 7c 7d 7e 7d 7a 75 7f 79 76 7b 7e 7c 79 78 76 74 70 77 70 74 76 6d 78 75 71 73 6b 6e 74 72 6e 66 63 62 60 59 55 4b 50 44 42 3a 3c 3a 31 37 3b 3c 42 39 2c 27 11 0a 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0c 0e 24 29 34 40 30 3f 39 3f 3e 41 40 3f 48 3d 41 37 38 4f 46 45 43 42 42 43 40 3e 45 40 44 32 3c 3d 41 39 44 47 43 35 3c 3b 3d 39 3e 43 31 3a 35 31 33 3c 36 3f 35 3d 35 3e 34 33 3e 36 33 3c 3a 37 34 30 39 37 3b 35 30 34 2e 2d 32 33 2c 30 36 2c 2f 32 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 34 6f 84 86 89 7a 7e 80 84 77 81 73 79 7e 74 7c 72 77 71 6e 79 78 7e 6f 76 79 6e 73 77 71 77 6a 75 6e 6c 70 6d 6d 58 62 58 5b 5a 5a 4c 48 4e 43 46 3f 3b 37 3e 3a 39 36 34 21 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 17 1f 22 30 33 2e 36 3b
 3b 39 42 3c 3f 43 39 44 3a 38 41 41 3a 45 43 42 41 41 44 45 3d 43 41 43 39 43 3a 3c 39 33 3f 3a 3d 3b 41 3d 3b 3c 38 3e 44 3f 41 39 3c 42 2f 3b 3a 3a 35 3d 35 38 3a 35 37 35 2c 36 33 32 37 3b 36 2f 32 27 2e 2f 2d 2f 27 29 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 31 6d 86 7e 85 7d 7b 7a 7a 74 79 7d 78 7e 71 76 7b 72 78 75 70 73 77 69 74 75 6d 74 6d 6e 6f 71 74 6f 6b 67 60 5f 57 5a 55 55 5a 4a 49 50 45 48 4a 40 33 41 3e 38 31 32 2b 18 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 07 1c 1f 27 28 30 36 35 35 3a 35 40 41 38 38 35 3d 39 39 35 3b 45 43 3b 41 41 3d 3d 41 32 42 44 47 45 40 44 3c 3e 3e 3b 3c 44 41 3b 37 3b 3a 40 40 35 36 38 3b 3b 3c 39 34 34 32 3a 3a 38 3a 35 2f 3a 27 38 2f 31 32 32 32 30 34 2f 29 2c 34 25 28 24 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 06 05 03 00 06 05 03 00 06 05 03 00 06 24 5c 81 84 78 71 74 79 7a 6d 6b 6c 73 76 74 6e 76 75 75 73 79 6c 6d 6f 6b 6c 64 6d 75 6a 6a 6c 6c 66 69 5c 5f 60 5f 58 53 51 4c 50 4a 4a 4b 4a 45 39 36 3a 3d 37 3a 25 1e 11 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 17 24 22 24 33 31 36 3a 34 3e 3a 41 36 43 3a 44 42 46 3d 3e 3f 3e 3d 42 48 36 3d 3b 30 40 3e 3e 3b 3c 3d 40 41 46 3d 42 3b 3b 3d 43 3b 3e 41 38 3b 42 36 3a 3e 36 39 30 30 36 34 38 34 35 36 37 3b 3c 2b 37 2d 33 35 2c 2c 30 34 29 31 2c 33 2c 2c 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 06 05 03 00 06 05 03 00 06 05 03 00 06 21 6b 7a 7d 73 6a 6b 77 73 70 6d 73 69 6d 6f 6c 6e 6c 74 72 77 73 6c 6f 60 66 6b 71 6b 6b 6e 68 64 62 62 68 63 63 52 53 55 46 46 44 52 46 46 4a 3e 3d 3d 35 33 30 22 1e 12 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 00 0e 1f 21 22 31 35
 33 38 38 39 3a 38 3f 3f 3d 42 39 3f 3e 44 40 3d 46 42 3d 42 47 3a 3b 41 3c 3f 46 3f 3f 40 3b 38 3e 3d 3e 43 3d 3e 3b 37 42 3e 3c 3d 32 41 31 39 41 38 38 3f 3f 35 32 3b 30 39 33 2e 2e 2e 37 35 3d 33 36 30 2d 2e 2c 2b 30 2c 27 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0f 06 05 03 00 06 05 03 00 06 05 03 01 06 26 69 79 7d 71 76 74 76 6f 6c 6e 6d 6f 6b 74 6a 71 69 66 63 69 6b 67 6d 65 67 72 69 67 72 64 69 64 5b 61 56 55 5d 58 52 54 49 47 42 49 47 4b 46 39 39 33 35 37 2c 1f 16 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0f 15 22 2a 32 2b 33 39 37 3f 3c 36 38 3c 3c 3a 3c 38 45 3e 38 40 3e 42 40 37 3f 39 3c 3a 44 39 3e 41 46 40 3c 3b 41 3d 37 3a 39 3e 3c 44 39 3c 38 37 3e 32 35 3b 36 33 3f 2d 34 3f 30 33 35 34 37 2b 36 33 31 34 30 2a 33 2d 2b 31 30 2c 2b 23 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 06 05 03 00 06 05 03 00 06 05 03 00 06 20 59 6e 7d 79 73 6f 6c 50 68 66 67 6e 65 6e 67 65 6e 70 69 74 6a 6b 67 65 6e 69 6b 67 65 61 58 5b 5d 5d 5b 50 50 50 56 4d 44 3f 44 3e 43 40 40 37 35 38 2e 2a 20 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 0f 16 21 25 2d 37 35 33 3a 39 36 35 42 36 3a 44 3e 3d 39 3c 42 3b 41 41 3c 37 41 3f 3e 34 39 3c 3c 3e 3c 38 3b 38 39 40 39 39 38 3a 3d 39 3a 3a 3a 3c 32 39 32 31 32 2f 34 34 35 33 37 2e 36 3b 30 33 36 2b 2c 2a 32 31 2b 34 2e 29 2c 2f 26 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 59 73 74 75 62 61 61 66 63 62 68 66 69 66 61 6a 6d 66 6a 67 5f 63 68 62 61 69 63 58 5f 5e 5d 53 54 58 4a 56 59 54 4a 42 40 40 40 3f 3d 3a 39 31 31 2e 25 25 15 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0c 15 25
 25 2e 34 30 32 38 3b 35 3b 40 43 45 3b 42 39 39 48 40 43 42 3c 41 3a 38 43 40 45 3e 3d 3a 3e 46 48 44 49 3f 42 3c 3b 41 37 39 40 37 3e 36 33 38 3e 3c 3d 3d 37 34 30 39 2d 36 38 37 2f 36 37 35 2e 30 37 2e 2e 2f 32 35 31 2c 28 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 15 4a 66 77 6d 69 69 6c 6c 63 65 66 69 62 69 69 67 65 63 5e 6e 64 5d 5c 58 65 5a 5d 5b 5d 59 51 4e 5a 4f 56 55 4e 42 46 45 3c 40 39 39 42 3a 35 32 2a 21 25 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 0d 15 1d 24 2b 32 33 3c 3d 3e 3d 3e 39 42 3e 42 3d 42 38 38 3c 41 3a 38 48 39 43 3f 3c 39 38 43 40 3f 45 3b 39 42 37 3b 3b 3b 3c 36 40 3b 3b 3a 3d 41 3a 3f 3d 35 3d 3b 3e 34 36 37 35 3c 34 3a 32 31 34 32 34 2d 33 28 39 34 30 29 2e 21 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 14 46 61 69 65 6a 69 61 65 65 5f 61 67 54 60 64 64 65 59 64 65 62 63 63 59 62 5b 59 59 54 51 51 58 51 45 5a 52 53 45 3b 3c 40 32 44 36 3e 3e 30 32 26 20 0d 0a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 0d 16 1f 25 26 34 36 31 2f 3b 36 42 3d 3b 3a 3e 45 3d 3b 35 3d 42 42 40 37 38 36 36 3f 3e 3a 3e 3d 3f 3e 3f 3e 39 34 3e 3e 39 3d 3f 3c 41 3b 36 35 3e 36 35 32 2f 32 38 3a 3a 31 34 32 34 3a 35 3c 35 30 2d 31 2f 29 32 34 2f 36 33 23 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 46 69 66 61 65 62 58 64 60 65 62 62 62 5f 62 5f 5a 5c 5d 61 64 60 52 5b 4e 58 51 4b 57 4c 52 49 50 51 51 4a 46 44 42 3e 2e 37 39 30 36 2e 30 25 17 15 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 0c 19 1b 25 28 34 33 3b 35 3c 3e 3e 3a 3b 37 40 3d 3e 3e 3e 40 42 38 3e 3b 39 40 3c 39 41 3e 42 40 3b 41 44 3b 3d 3f 3a 45 36 43 3e 38 39 35 3d 43 3c 3b 36 36 39 37 3d 37 33 39 37 34 41 35 37 2f 29 35 34 33 34 39 35 40 3b 37 35 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 3d 5c 6c 68 62 5f 62 5d 63 5e 56 5e 5c 67 5f 60 5d 59 62 59 5b 5c 52 54 54 54 50 52 55 54 53 52 52 51 4f 45 48 3f 3f 3a 3b 3c 38 3c 2e 25 25 1d 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0c 1a 1b 1e 2d 34 35 36 41 38 39 3d 35 44 3b 39 41 37 3c 3a 43 40 39 37 40 3e 40 3a 41 3f 3f 46 43 39 42 42 3e 3e 42 3e 3e 40 35 3b 40 3e 3b 39 38 3e 3c 35 3b 36 35 3d 3f 32 34 3a 3a 2f 33 36 34 31 2d 33 34 36 40 3f 46 49 38 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 38 56 6a 64 62 65 5c 61 53 5b 5b 5e 61 60 5f 51 55 58 56 54 51 57 53 4d 4e 45 4d 4b 55 51 57 57 59 56 4f 3e 40 3b 37 3b 33 31 37 33 28 21 17 08 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 0e 13 20 26 2d 2c 38 33 35 3d 38 42 43 36 3a 36 42 3d 40 39 2f 3c 3d 43 3b 35 44 3f 44 43 44 45 40 3b 44 3d 3a 3f 40 44 42 45 43 37 3c 3c 40 38 36 38 33 35 3b 37 2c 32 39 3d 31 3b 3e 31 34 34 32 35 33 37 38 43 4f 55 5c 44 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 3a 60 64 62 52 5b 5c 58 57 57 5a 56 51 59 57 55 53 52 55 55 4e 50 4b 4a 48 51 4d 52 55 56 5b 56 54 46 3a 3a 3a 3c 3c 3f 37 3b 2a 2a 2a 1a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 03 06 09 16 20 1f 25 31 3a 3c 3d 40 42 3c 3a 38 3b 42 3c 3a 3c 39 3d 44 3c 3e 3d 39 4a 4a 4e 51 47 4a 47 47 42 3f 4a 39 3f 42 41 3c 39 38 3b 42 3f 44 3a 3f 3d 3a 40 37 33 3e 38 38 3e 39 3c 37 3a 35 30 39 35 44 53 5c 64 66 4d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 38 5e 64 61 5c 55 5f 56 59 57 55 57 59 59 53 4b 50 4e 47 51 4e 4d 49 4c 4d 53 52 56 5d 51 54 45 43 41 3a 3d 3a 34 3c 31 36 2a 26 1f 1d 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 10 1a 25 22 2e 32 38 39 3b 3a 3b 34 41 36 3b 39 3e 3f 41 40 3b 44 42 4e 50 56 57 58 53 56 54 41 48 44 3f 3d 47 46 47 41 4c 3c 41 3f 3d 46 44 3a 45 3a 3f 40 39 3b 3a 3c 38 35 42 31 3a 39 3e 38 45 54 55 59 68 65 51 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 33 54 62 59 58 5a 52 56 52 55 55 56 53 52 4d 51 50 48 45 47 49 53 4d 4d 4c 50 54 5f 53 4e 48 46 46 3e 3e 38 35 39 32 30 2b 26 20 17 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 12 1c 28 22 31 37 3a 43 35 33 3b 3b 41 3d 48 41 3a 49 44 47 45 4d 56 55 61 5b 62 56 58 57 46 42 45 3f 42 46 44 47 46 42 45 43 3f 41 3f 44 3b 40 3c 3c 37 42 3e 39 3f 38 38 39 37 3b 39 3f 42 4e 57 5c 66 5e 51 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 2c 56 59 58 5c 58 52 51 4c 50 4c 4a 4e 49 49 49 46 4d 47 49 4d 4b 50 47 51 54 49 50 4b 42 3e 3c 3d 37 33 36 37 30 2f 29 1b 13 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 05 06 0e 16 25 22 2c 33 3a 3b 41 3a 38 3c 43 3e 43 3e 43 48 4d 48 46 4c 59 5b 63 5c 5e 63 64 55 54 52 4a 50 44 47 44 3f 46 42 45 49 3e 47 42 3d 3f 41 44 3d 36 41 44 4a 3b 3d 3a 38 3d 36 3b 39 47 47 59 59 53 51 45 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 4e 5a 57 4d 4f 48 4a 48 4e 4d 50 45 4e 44 44 4e 4f 42 4b 44 50 4c 4e 4c 4a 49 48 43 41 3f 3d 3a 3f 32 2f 34 2d 25 1c 12 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 16 1a 22 30 33 31 44 3b 3d 41 42 41 46 4c 49 54 4a 4e 48 4e 58 59 63 67 68 66 60 60 5c 58 4a 4b 46 46 47 48 48 40 40 45 46 3c 42 48 3e 41 3a 41 3d 3c 43 42 45 3a 37 3b 3a 35 39 3d 42 4a 49 4a 46 4e 3b 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 43 4b 4c 4c 43 52 4d 3c 43 4d 44 48 4b 49 50 50 4b 4c 4f 4e 4a 4f 44 48 4d 3b 3a 37 3d 32 3b 3a 35 36 39 2d 24 11 12 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0d 17 1e 2e 29 30 2d 3a 39 43 47 47 51 53 52 56 48 4e 50 4d 52 59 5c 5d 5c 5d 61 5d 53 58 4d 41 3c 47 41 43 46 47 40 3d 38 3d 3d 47 3a 35 41 36 36 35 3c 3d 3a 38 35 33 30 38 3a 31 41 3f 3d 46 3e 35 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1a 40 45 44 45 46 48 46 41 3b 44 48 47 4b 42 4b 4b 4d 48 4b 4c 4d 40 3d 39 42 3a 3a 36 39 31 3b 2f 2a 2a 26 20 13 0d 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 0f 1e 26 2b 2c 32 43 3d 4a 4f 4b 52 5b 57 4e 4b 4a 53 57 55 54 52 55 58 5d 5e 50 4c 4e 4a 48 4d 47 46 36 40 45 42 46 46 38 3f 36 39 3b 3a 31 2f 32 34 37 37 34 31 32 3e 2f 31 40 36 35 34 32 2e 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1d 3c 4b 44 43 3b 3f 3b 44 45 43 42 47 41 3b 40 4d 4e 45 43 3d 47 3e 37 38 3c 3a 39 39 38 3a 34 25 21 24 1f 0e 04 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0f 0f 17 2a 27 2e 3e 3e 4b 47 54 56 52 55 54 5b 5c 57 51 4e 57 51 54 4c 56 52 4f 59 50 53 4d 4a 51 4f 45 4b 40 3d 3e 39 37 3a 35 33 36 38 39 35 35 34 27 32 2e 31 32 35 31 3e 41 33 3c 37 28 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 34 45 47 3b 47 3b 41 41 3d 40 44 3f 42 44 41 3f 3f 46 44 3a 36 35 3d 37 36 38 33 2a 2c 26 19 28 1f 15 0f 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 17 15 2a 2a 31 33 39 44 44 4f 5e 57 5c 54 56 55 58 51 52 4e 45 3a 50 46 50 50 4e 54 55 58 50 54 48 49 45 41 45 38 3a 39 2c 32 2b 29 30 31 2d 22 26 2e 2e 38 2d 34 29 38 3b 2b 33 33 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 42 47 39 3d 39 3b 44 48 41 3f 40 40 3d 3c 41 45 3c 3b 41 35 3a 3d 33 3a 36 2e 2c 29 20 29 16 14 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 15 1b 27 36 3a 3e 3c 3f 47 50 56 56 5c 54 58 55 58 55 51 48 3f 42 4a 50 5b 52 4c 51 4e 55 52 4d 46 48 3e 3c 3b 36 2b 2f 30 35 38 2b 29 2d 28 28 2c 2b 2b 26 2f 31 27 2b 23 22 25 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 30 35 42 37 35 40 37 3c 46 38 3b 40 38 41 44 3c 3c 34 3a 30 3b 33 2f 2f 30 29 25 29 1d 1e 18 0d 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 07 10 1f 20 2d 31 36 3e 45 4c 49 47 50 52 5b 57 53 55 50 49 42 47 44 48 42 4e 4f 50 55 55 4d 4b 46 45 3f 3c 39 32 25 2e 2e 33 30 29 2c 25 29 27 2a 27 28 2b 2e 31 25 27 23 2a 1e 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 33 3b 39 3e 3d 3b 3d 3c 37 42 3d 3e 2b 3b 37 38 3a 3b 35 40 33 23 32 29 31 22 1f 1b 16 0e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 11 0f 1e 19 26 35 34 3c 38 40 3f 48 4b 51 52 53 4d 3d 40 3d 42 47 43 41 4c 48 45 47 48 49 47 3e 3b 37 34 37 2f 2c 28 2f 2a 24 30 26 23 2a 21 21 25 1c 29 23 2a 23 2f 29 1b 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 2d 39 31 37 3b 34 3b 36 36 33 36 37 32 33 32 2a 31 36 2f 2e 29 27 26 21 21 1a 18 0f 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 09 12 19 14 24 23 28 34 38 2f 35 48 42 45 45 47 43 3f 36 39 3d 3c 3a 41 41 49 3a 42 38 3a 34 2c 30 2f 2c 2a 2d 29 25 2a 2a 2d 22 2d 20 20 23 24 29 24 1d 26 1e 23 21 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 28 2f 25 33 33 2a 37 31 28 29 2a 2c 26 2b 37 1f 29 2b 2a 1e 23 17 13 16 0f 10 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0f 10 16 1c 1f 29 37 35 3a 2d 33 35 41 3c 34 32 39 3e 39 38 3c 38 31 3b 36 3d 39 31 2b 2c 2b 2d 2c 25 2f 21 2d 29 21 29 23 29 21 23 22 25 27 1f 25 21 1f 1e 1f 22 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1e 2b 28 26 2d 2c 33 25 2c 1f 24 26 29 2b 25 23 24 20 1e 1f 1e 16 13 0c 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0e 0e 1d 23 1d 29 30 36 2c 2f 30 33 36 34 2e 2e 2b 31 33 32 2f 24 2a 33 2b 22 27 22 2c 27 28 2a 2b 1d 27 21 23 27 1f 20 1f 27 24 1c 24 17 1f 1d 1c 21 1a 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 15 12 19 15 24 1b 1b 20 26 1b 15 1b 20 20 1b 1f 14 1a 15 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 08 16 0f 17 21 2c 1f 24 2a 20 25 26 23 2c 26 25 27 1f 20 16 21 1c 1a 1b 1f 22 24 27 21 22 1a 1e 22 14 1f 22 22 1c 18 19 1e 17 17 1d 17 19 13 17 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0e 0a 0b 0e 0c 0d 10 0f 0d 0a 1c 17 0f 14 0f 0b 06 0a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 0b 19 18 17 24 1d 2c 24 1d 24 23 1f 1c 1d 10 11 0d 16 16 12 13 1c 24 1d 21 21 18 20 1a 1d 19 1f 23 1d 16 15 14 11 15 14 14 17 14 0b 11 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0d 05 10 0a 0b 05 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 07 14 18 1b 1b 1e 19 19 16 10 0c 0d 05 06 05 0f 07 11 0b 17 1b 1c 1a 10 10 14 10 0a 14 0d 0b 15 0f 0f 0e 10 07 0b 0e 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 05 08 06 05 0a 09 06 05 03 00 06 05 03 00 08 06 09 0b 06 07 06 00 06 09 06 0e 06 05 07 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
