 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 04 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 02 06 05 03 00 06 08 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 01 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 01 06 05 03 00 08 05 03 03 06 05 03 05 06 05 03 09 06 05 04 00 06 05 03 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 02 06 05 03 00 06 08 03 02 06 05 08 00 06 05 03 07 0e 05 0b 03 06 09 0a 01 06 05 03 03 08 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 04 0b 0d 0b 0d 0e 0c 0f 0c 12 06 08 03 04 06 05 0a 05 06 06 03 00 06 05 07 06 06 05 04 00 06 0a 03 03 06 05 03 02 06 05 05 00 06 05 03 00 06 05 03 07 06 07 03 00 06 05 03 03 06 05 03 02 06 05 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 06 06 05 12 0a 06 05 03 00 06 05 03 08 06 06 0b 01 10 09 0b 08 08 0b 06 0e 06 05 05 04 06 05 07 04 06 05 05 00 06 05 03 09 06 08 0a 0a 0d 0b 12 14 0c 0e 0a 0f 11 09 08 0e 06 05 09 05 09 08 0a 0f 06 05 05 09 08 05 09 01 06 05 03 01 06 07 03 02 06 06 04 00 06 05 06 04 06 05 03 00 06 05 04 02 06 09 03 02 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 04 04 06 05 03 04 06 05 05 00 0a 08 13 16 0d 05 03 0a 0d 07 0e 0a 0a 05 0b 15 0e 07 0a 05 11 15 08 06 0a 05 07 05 06 08 03 05 06 05 03 08 06 07 04 09 06 06 0d 0e 10 11 1a 18 13 14 10 1a 17 14 0b 11 10 11 0d 14 15 13 1d 16 10 09 0b 09 12 0e 0d 0b 0a 12 10 0a 06 0a 0e 06 06 05 07 06 06 05 03 04 06 05 05 01 06 05 06 0e 06 08 03 00 06 06 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 01 06 0a 0b 05 10 05 09 06 0d 05 0c 0d 0c 11 0b 0e 06 13 04 09 19 12 16 06 09 08 06 10 15 11 13 1a 1c 1c 0d 07 06 05 0a 08 09 0a 08 06 09 05 04 09 0e 14 08 1e 22 22 21 1c 17 1f 27 2d 31 2f 2f 3d 33 30 2a 29 23 2b 2a 30 2d 2c 1a 22 26 23 1f 1b 25 1f 14 1c 16 14 17 13 16 16 1d 19 07 0c 11 06 0a 06 09 0e 07 05 03 07 06 0a 0c 11 06 05 05 0c 06 05 03 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 04 04 08 05 04 02 06 08 03 07 0a 05 0a 07 06 0c 08 0e 13 14 0c 1a 11 15 1a 16 1f 19 16 16 10 1a 20 24 29 2f 37 3e 41 44 22 1a 1c 13 18 0f 11 0f 18 0e 0c 09 05 10 0e 16 1f 2a 4c 4e 42 3f 35 3c 44 52 52 55 59 5e 65 5c 53 46 44 4a 42 47 3f 3f 3e 3e 3e 44 39 3b 35 2d 29 31 31 28 23 29 28 2d 2d 2b 17 0e 0e 19 18 12 17 05 12 11 0d 05 13 06 13 0f 0f 0e 08 0c 06 06 03 09 06 06 0e 00 06 05 03 02 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 07 09 04 09 07 0d 0f 09 0b 04 11 10 0c 12 0d 16 14 10 1c 21 23 26 27 25 29 2f 2f 2d 34 34 45 55 5e 70 60 51 45 46 39 2b 32 2e 2c 2d 38 2f 1e 0c 0f 0f 25 31 21 2b 54 73 86 77 6e 69 5d 72 70 81 80 76 7e 70 6f 52 55 47 44 3b 40 44 36 43 49 42 45 4c 42 3e 47 3c 3a 2f 2e 3c 3d 42 44 3d 40 3e 35 2f 24 20 14 15 20 28 25 1c 1c 1a 13 1b 1d 0a 12 0a 09 10 0a 09 07 06 05 05 09 0e 05 03 00 06 06 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 06 06 05 00 06 12 0b 05 06 07 0e 15 16 16 13 18 17 1e 1e 29 2b 28 27 31 35 38 42 44 44 50 54 5e 68 69 72 85 86 92 89 74 5a 58 4c 46 40 45 40 43 4a 50 4b 3e 1f 1e 23 3d 49 50 55 5b 6f 76 7c 87 89 88 86 8c 85 79 67 64 61 54 46 4b 41 3e 40 44 50 41 44 42 44 44 44 4f 46 45 41 41 47 49 4d 4c 44 49 4e 55 5d 81 71 54 4a 3f 33 3b 39 36 2d 2d 25 26 19 20 1c 1f 17 14 15 15 16 18 08 05 0f 14 0d 0c 0e 00 08 05 07 0e 0a 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 00 06 05 11 00 07 05 05 0d 07 0c 0f 14 0c 18 15 11 18 1e 1c 16 1e 1f 2a 2f 2b 3a 3d 3e 3b 49 3e 4f 60 5f 75 72 81 83 82 8d 96 97 97 ab a8 9f 89 6e 65 58 59 59 51 56 4f 59 5b 5a 5e 56 4b 40 49 54 5a 62 5f 5a 61 61 62 66 70 6a 6b 6f 6a 65 57 53 55 47 4e 47 44 4a 42 44 41 45 43 43 4a 4a 4a 47 3f 48 4a 46 4d 4a 4c 49 4e 51 54 53 61 89 a2 95 7d 66 5a 5c 5d 58 4a 53 40 3e 47 36 3d 33 2a 23 2a 25 2b 2d 1e 1f 1d 11 13 1d 0e 0a 0b 06 0e 0c 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 09 0b 09 03 0a 0d 12 0f 10 10 14 12 16 18 18 27 27 3c 43 44 4c 46 48 4f 49 4c 4a 52 65 72 6f 79 8b 98 9c a3 a7 ab b4 a9 b5 b8 bb b2 a6 8d 6e 66 60 5c 5c 54 61 5d 5d 5f 59 60 59 5a 5c 6b 65 60 5d 5c 61 65 5e 61 5e 59 5b 59 5a 53 55 53 50 4f 55 4e 41 48 40 49 3b 4e 4d 43 43 4a 47 4a 44 4b 4c 52 51 4e 4f 4a 48 4d 4f 5c 59 5f 65 78 a0 b7 b7 9c 8c 85 85 8d 7b 71 6f 60 6a 67 62 5d 4e 4e 46 4d 42 3e 33 33 2b 28 24 2c 1d 1c 13 08 09 15 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 05 00 06 10 05 0b 06 0e 10 09 09 14 16 24 20 18 25 25 2d 3a 3a 49 62 6b 7c 76 7f 81 84 7a 78 80 82 8b 8f a7 a9 b0 bd c9 d4 cf da d8 d5 d7 d0 c0 b1 8c 79 68 5f 67 5e 59 5c 61 61 61 62 62 5a 5f 5f 67 60 65 65 66 69 6b 63 65 6b 65 60 5d 54 5c 5a 58 5e 51 52 4a 4f 51 49 46 43 4a 47 4c 4a 4d 4f 50 52 50 4b 51 54 52 51 54 54 54 51 51 51 56 5a 5f 62 6d 7b 9a c0 c5 c2 bc b8 b4 ad 9e 98 98 90 8c 85 76 61 5d 5f 5f 65 60 4f 54 56 4a 42 35 3b 33 2a 2e 1e 17 1a 12 16 15 0a 09 0a 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 02 0f 09 11 11 11 06 17 11 14 28 2a 29 36 44 46 4a 5e 67 7c 92 aa b7 b8 c3 c3 c0 bd b7 ab b2 b3 ba c3 cd d2 dd f8 f2 f5 f3 f0 e4 d5 c5 af 96 84 68 62 5f 5b 56 60 5f 57 5f 5f 62 65 61 63 62 61 64 6b 6b 69 70 6a 65 68 67 6a 66 60 5e 65 5e 59 59 63 58 49 56 4e 52 45 50 4d 48 4a 50 4d 4d 4f 57 4f 56 5a 54 54 5c 5e 55 54 55 53 5b 4d 5e 59 62 6b 71 75 80 8e a5 bd cc d4 c7 c8 c3 b9 b5 ae a8 93 80 5b 58 55 5d 59 5d 5c 63 67 62 62 68 57 47 3c 31 30 20 28 28 26 21 21 12 0f 0b 06 07 0a 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 07 03 11 09 11 1a 0b 15 14 20 25 2a 35 47 50 60 71 79 7f 81 87 85 99 bc d7 ed fc fe f2 f1 e8 df e1 e4 e4 f5 fd f9 fa f7 e5 db c8 bd a6 9b 94 85 7f 6f 6d 65 63 5c 5d 66 57 59 63 65 64 5d 67 58 6d 67 66 65 6b 66 67 6b 65 65 6b 64 66 60 62 61 52 5b 55 53 5b 51 5a 50 59 4c 4e 49 4f 47 4f 4f 4a 50 53 54 58 53 5a 51 55 57 52 59 59 54 5f 5e 62 62 60 68 6d 6d 75 6d 7e 8b 99 b5 b7 b9 b9 b6 b0 a0 82 7d 66 5c 5d 65 5d 5f 5b 57 5f 60 7c 81 84 77 6d 56 4a 3f 34 2f 38 33 2e 29 1f 10 10 06 13 0c 09 0f 06 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 10 05 0f 01 06 06 18 19 1d 14 22 26 35 3e 4c 4e 47 5b 5c 6d 7c 87 93 8d 88 84 85 8d 9b a6 c5 da f4 f7 f7 fb fd ff ff f1 ed e5 d5 cb be ad aa a7 9f 94 87 8d 85 84 77 6f 70 60 5f 61 64 60 58 5c 60 5e 62 6a 6c 6d 6e 6e 6f 6d 6a 6d 6c 64 6b 6a 62 69 5f 5c 66 61 5f 61 65 57 5a 5b 54 4b 48 4a 4d 51 47 50 55 4c 4a 54 56 5d 60 5a 62 60 60 65 55 5c 5b 5f 64 5f 6a 67 61 72 77 71 75 72 78 7a 7f 84 80 85 8a 75 78 70 67 65 5b 60 65 64 62 5b 64 64 68 7c 8b 98 9c 83 7c 78 5c 52 4e 58 5f 4c 34 27 18 1d 11 17 13 10 14 11 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 02 0a 05 04 0d 11 0b 0c 18 11 19 16 1e 23 2f 43 4a 5c 65 60 5f 64 67 66 73 79 8b 95 8f 8f 8c 85 90 8a 93 a3 a8 b5 b7 c3 c9 cd c8 d4 cd c3 b6 ad a7 a4 a5 9d 96 9a 95 91 8d 88 83 7b 79 75 6a 69 6b 69 5f 5f 5e 64 66 65 73 70 72 72 70 76 73 77 79 75 75 6c 6e 69 6a 62 65 66 68 62 64 66 5c 56 60 57 5a 55 50 4f 58 50 5b 52 56 56 60 5c 60 60 5f 61 65 63 5e 60 65 62 65 60 69 60 69 6e 6f 72 73 77 73 71 78 79 70 6b 66 6c 74 73 67 69 6a 64 65 64 6f 64 64 63 6d 69 68 75 89 90 90 8b 79 5e 5f 6a 78 82 6f 55 3f 2f 28 27 2a 20 27 17 14 0a 06 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 0a 0f 08 07 10 0a 14 17 10 21 1f 25 36 47 49 56 60 70 76 70 62 71 69 76 79 7b 7b 8e 92 95 8b 8a 97 88 9b 97 9f a7 ac a4 a8 a1 aa b0 a7 ac a7 a3 a7 a9 a1 99 96 9e 8f 94 91 90 8d 7c 76 82 6c 71 6a 64 63 60 65 64 64 68 70 6f 75 71 78 74 7e 72 6e 78 7d 70 75 64 6b 68 65 66 69 63 69 67 64 5d 5e 55 5b 5b 57 4c 57 53 52 5b 5a 56 5f 5b 5d 5f 61 60 64 64 5d 59 63 63 61 63 61 61 69 70 74 6e 6e 7d 74 68 6f 73 6f 6e 6e 64 6e 6b 66 67 6d 6a 63 70 69 67 70 67 69 64 66 64 74 74 70 70 6e 60 65 74 92 a7 8f 76 5a 4f 47 36 3b 35 31 2b 1d 13 12 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 11 18 14 0b 14 0e 1b 21 24 2b 38 4c 55 57 68 69 78 7f 78 76 6f 6d 75 74 7d 85 82 89 8f 95 99 96 8d 8b 8e a3 9d a2 b5 b1 a4 a6 a9 a7 9c a7 a9 a3 af aa a5 9e 9b 95 8d 8b 95 92 93 86 82 7d 77 77 71 6b 71 6d 6f 66 6e 72 75 76 77 77 7e 7d 75 7d 81 7b 7d 77 79 71 6f 70 6f 6a 70 6d 6e 6c 67 5b 64 62 64 58 5d 5b 5b 5b 59 57 54 59 55 5c 65 69 64 61 69 63 64 67 65 61 5f 65 64 67 65 69 72 7b 73 77 76 70 6b 70 6f 72 6a 66 6f 71 6a 6c 6f 6e 65 70 6b 70 6e 6b 69 67 67 6d 70 6d 6d 6f 6b 65 67 6c 87 a8 ac 99 80 6f 60 53 64 54 4b 2f 23 1b 23 1a 16 0b 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 06 06 05 0b 0b 06 09 10 0c 13 18 13 1e 20 24 36 3b 4f 5f 61 65 71 75 75 76 84 7c 7b 74 79 7a 80 7e 85 87 8a 8e 97 99 92 92 8d 96 9b 9f a5 b6 b5 af ae af b0 ad ae af ad ad b3 ac a2 a1 a1 a4 9c 98 95 8d 8f 87 85 7d 7f 78 75 70 64 72 75 70 7b 7a 83 86 79 87 7e 80 7e 7c 84 81 7d 7b 7d 70 6d 7f 7d 77 71 67 6e 6a 6a 68 6d 68 60 63 67 5c 5c 5f 5e 5e 63 68 62 6d 63 62 69 6e 72 68 67 68 5f 61 63 6c 6e 72 70 6f 7d 75 76 76 77 78 78 6b 70 6f 71 73 74 76 74 70 69 6e 71 6f 6e 76 77 72 6f 6b 6f 6d 72 6f 70 6c 65 6f 6b 7a 8e a9 b7 ac 9a 99 88 87 6b 60 4f 39 2a 2f 2d 22 1b 0f 0a 0d 05 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05
 0f 09 0f 10 12 10 1e 23 27 31 3c 47 4e 6f 7a 86 76 6f 76 77 7a 80 83 80 8a 7d 79 77 7e 7a 87 89 89 85 8f 92 92 96 8d 98 9e a2 a8 be ae b5 b5 b4 bb b0 b2 b3 ad b4 b0 aa a1 97 9d 9a a0 9f 9d 9c 92 8d 86 88 79 7d 80 7b 78 78 7e 7b 7a 7a 85 84 83 88 86 87 80 8b 7d 84 7d 84 7c 7a 77 7e 7e 7d 7a 80 78 79 74 6e 6b 74 73 66 5e 66 5b 5c 68 5b 5e 69 6d 6d 6a 6c 6d 71 72 67 67 64 60 61 65 64 69 6d 6b 74 6f 78 7c 7e 7c 79 75 75 73 73 77 75 73 74 77 7a 70 76 79 74 79 70 75 72 7a 6f 74 73 78 71 73 70 6d 74 74 72 77 87 a5 be b8 c0 b1 aa 8f 7d 6a 5a 41 4e 47 35 2a 26 16 12 0a 07 11 1e 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 0e 13 1a 1c 21 1a 1f 1f 25 2e 48 5d 66 7e 83 89 95 83 79 74 78 7d 7f 7f 83 7e 86 7e 80 7f 80 8a 88 84 87 89 85 8e 8f 97 95 94 9f a5 a8 ae a3 a4 bf bb b7 be b6 b2 b5 b3 af a0 aa a0 9f a2 9c a7 a0 99 93 96 91 87 8b 7e 8b 84 7d 7a 84 7a 85 88 89 8c 93 95 92 94 89 8e 8c 90 8b 86 83 84 84 85 88 83 80 7e 7b 7e 78 7b 81 7e 79 72 70 6a 65 64 69 60 6b 69 60 67 61 6f 6a 68 72 71 69 6b 6b 66 61 67 66 6d 74 6f 76 72 79 79 7c 7a 74 7e 72 79 78 7e 85 73 7a 7f 73 7d 84 7e 79 79 76 78 77 79 77 7d 76 7b 7d 76 6f 75 65 6e 74 76 84 93 af c1 c9 c2 b9 a4 85 7d 70 79 68 5b 46 2c 13 0e 0e 0b 0e 1d 20 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 01 06 05 03 07 06 0a 05 03 06 06 04 06 1a 27 25 25 29 2b 34 44 4e 5e 6e 84 8b 97 99 99 86 83 75 76 7b 7b 7f 81 81 83 7f 84 81 84 7e 7f 8a 8c 95 8e 93 94 91 93 9c 9b a0 a9 b1 c0 c1 c7 c2 c9 c7 c6 c1 c5 b1 b2 af b0 a3 a0 9d a5 9c a0 a0 90 9f 93 92 96 8c 8b 90 8a 89 89 88 8d 91 95 90 91 a0 8d 97 94 9b 92 8d 95 92 8e 8f 93 8d 8e 85 8f 89 8f 85 84 85 7d 87 7c 83 86 7c 73 75 72 6a 6c 67 6e 65 6e 6a 71 74 6d 75 74 65 72 6d 70 6d 6d 66 6c 70 71 77 82 7a 78 7f 79 7b 83 80 7d 80 81 7b 86 7d 78 86 8c 8a 7a 7d 7f 83 7b 71 78 78 84 76 78 7c 7d 75 75 74 73 73 72 71 79 80 96 b4 c7 cf ca b9 ad 9b 90 88 88 70 45 27 0c 12 0d 07 0b 1e 13 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 09 03 07 06 05 0f 01 06 1b 10 19 1f 20
 32 2e 35 41 59 66 7a 91 a6 b3 a9 98 8c 83 7c 7c 7a 77 85 8b 79 86 84 82 89 85 84 84 81 86 8c 8e 9a 98 9a 96 92 9d 9a 9c a4 a1 b3 c5 c1 c7 cc c4 d0 ca c5 bf c5 be b4 a8 a2 a9 a7 a8 a3 a4 99 a0 94 9a 9d 90 95 8d 93 9b 97 95 9c 95 9a 97 9b 9c a5 a7 9e 9a 9c 9d a2 96 9c 99 93 9a 95 94 96 95 94 93 8b 91 89 8b 87 88 81 86 7f 7d 73 76 6f 76 72 6f 76 7b 71 70 77 73 76 74 6b 6f 6f 6d 6a 6e 67 72 74 7e 7a 7a 84 84 7e 84 7f 84 7e 86 88 8d 90 80 90 8b 8d 8f 93 8d 87 80 7e 84 81 85 7d 8b 86 82 81 7f 73 73 7a 75 73 72 75 75 85 7e 88 95 a7 b3 b5 b2 98 90 8e a2 99 67 3e 26 18 10 15 18 1f 1c 0f 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 06 05 03 01 06 07 07 14 12 14 1c 2b 2a 30 3a 4c 57 6a 7d 83 a3 bf d0 bb 9e 82 80 7e 75 7b 85 7f 7c 89 8b 7f 88 89 86 8b 8a 84 8a 8c 8b 90 9b 9c 96 9e 98 a0 9a 96 a7 9e b6 c1 cc ce cb d6 c7 cc cb c7 be bf ba b1 9d a7 a0 a5 a4 a1 a1 a0 a0 98 9d 9b 9d 9a 9b a3 8e a3 a1 a7 a5 9e a6 a2 a8 ac aa a5 a4 a6 aa a8 a2 aa a2 9c 9b a0 99 9c 97 91 8a 91 8b 8e 8d 8f 90 8c 8d 87 77 79 77 71 73 6e 75 78 72 79 78 74 6f 73 75 66 6e 64 66 64 74 71 77 75 7e 81 7f 82 84 86 83 8a 8e 8f 8a 92 8e 8f 90 94 8e 93 92 8c 8d 85 85 89 88 8b 8c 83 8b 85 7e 7d 78 74 71 77 78 7b 76 75 7d 81 85 7e 7d 8b 8b 84 83 8e 93 b0 9e 70 4f 3f 27 1d 18 11 1b 1a 11 0d 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 07 01 0a 08 0c 09 10 13 19 18 1b 31 2c 36 42 40 5b 72 7e 88 9f c2 d4 da c9 96 85 7d 82 85 82 7c 7d 84 87 84 87 8b 8d 90 8a 88 8a 8e 83 8a 93 97 9d a8 a4 a2 9d 9f 9a 9d a5 a9 b4 bf c3 d1 d9 d5 d7 d1 ce cd c4 c8 bb b1 ac a3 a5 a5 a2 a4 a5 a4 a9 a3 99 9f a5 a0 a0 ac a4 aa ab a7 b1 b3 a5 b0 b1 b2 b4 ad af af a8 ae ad a4 a4 af a5 a8 a3 99 a0 9b 9f 99 8f 95 94 95 93 81 8b 8c 89 8a 88 76 81 74 6e 6d 73 74 77 71 72 79 6e 73 68 70 68 68 66 72 7a 79 81 81 89 8b 87 86 88 91 8f 93 94 91 9d 9c 9a 95 95 98 9d 9e 98 8d 8b 89 92 8e 93 93 88 88 87 84 7d 7e 79 7c 78 7d 7a 7c 79 7e 75 82 7f 8c 82 8b 7a 87 9a aa 9b 72 5d 57 4d 3e 24 20 19 10 0c 06 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 06 0b 0f 0b 0f 12 10 1b 24 2a 3d 3e 47 66 73
 7a 8b 9e b6 d1 df d2 a7 94 8a 7f 86 83 8f 77 83 8a 8a 90 8d 91 95 8e 99 a0 93 91 99 93 94 8e a3 a8 a6 ad ab a8 a6 a9 9e ad af b7 c8 d0 d8 dc d4 d8 d1 d5 c5 d0 c6 c4 b5 ae a8 a7 a7 a4 ac ab a3 a5 9f a5 a3 ac a4 a5 a5 a6 ae b4 b6 b7 b9 b9 b7 b4 bd b7 b8 b1 b5 b5 b6 b7 ae ae aa ad b0 a6 a7 a4 9e 9e 9f 98 99 9d 9b 9a a1 95 91 85 89 82 7e 7c 80 7d 7d 75 72 7d 76 7a 78 73 72 72 69 68 74 74 6b 73 75 81 85 8a 8c 8f 8f 95 92 9b a2 9b a1 a1 9f 9f 9b a3 9f 9c a5 9d 95 9a 9d 9c 99 9a 99 93 90 86 84 83 82 81 84 7d 7d 80 78 80 7c 81 7f 80 7d 85 83 88 84 9c 99 98 71 60 58 5e 5a 4c 2f 25 13 0e 05 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 04 0f 0d 0c 0f 0d 16 17 22 26 39 50 52 6e 81 8d 9e b0 c4 da e8 c6 a9 89 84 88 8a 7b 88 8a 8d 85 8e 8d 85 8c 91 9f 9f 9f 9f 9e 9d 9c 93 94 93 a3 aa a5 b3 ae b5 a8 a4 ac b2 ac ba c6 d0 d7 dc dc e0 e0 d7 d0 cd c8 b9 ab b3 a3 a2 aa a2 a7 a4 a4 ac a3 a3 a4 a7 a5 b0 ae b0 b1 b2 b3 ba b5 b9 bf bd c2 c1 c4 be bc b9 ba bd b6 b8 b1 b5 ad ab ac ac a4 9f a9 a3 a0 a9 9e a5 9f 94 99 8f 91 8b 7e 84 89 85 81 7a 7f 7e 76 79 6e 77 78 73 75 70 75 72 6f 77 7e 8a 85 8b 90 95 98 9c 95 99 98 a3 a8 ab 9f ac a4 a5 9d ac 9e a3 9e 98 a1 95 90 95 95 94 8b 97 86 88 84 83 89 8a 86 85 7c 7d 7a 84 80 84 80 82 88 83 86 94 a2 8c 6d 62 63 66 61 5d 4b 34 2c 15 08 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 07 0d 08 08 0b 15 16 1b 25 2d 35 44 57 7a 8a 8f a5 a7 c1 d0 dc dd b7 9b 8c 8b 89 98 8b 8b 8b 8a 8d 8c 90 8e 96 94 96 9d a9 a5 ab a2 a2 9c a3 9b 9e a7 b8 b3 ba c2 bf b0 ad b5 b7 c2 c8 d3 d5 da e1 e3 e1 df d7 d1 d3 d0 c2 b6 b1 a5 b0 ac af ad a5 a1 ad a3 a2 a4 aa a4 af b1 b1 b4 ad b7 b9 c6 bd c6 c0 c1 bb bf c1 bf c2 bb ba ba b8 b1 b2 ae b0 ba af ac a8 a4 a3 a4 a5 a9 a8 a3 9d a8 9c 94 8a 92 8e 8c 87 84 6d 7d 78 7e 81 73 7b 7e 76 78 6e 6d 79 7c 7c 7b 85 86 8c 92 9f 9e 99 ae a5 a1 ae ac ae a5 af a9 a6 a5 ab a2 a4 a2 a6 a6 a2 9c 97 9a 90 8f 8b 92 8d 90 88 84 89 87 80 89 80 85 82 86 8a 84 88 8e 84 85 97 9f 8a 79 67 78 79 70 65 66 5b 3a 2f 1f 10 09 06 05 03 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 15 14 18 13 17 11 1b 16 24 37 42 52 68 78 94 a1 ab b7 c3
 ca c3 b9 a9 91 8d 8f 8d 8c 8f 86 94 92 8e 97 8d 92 94 97 99 a2 a7 a5 ad b1 ac a9 a9 ac a1 a9 b4 b0 c2 c5 d2 c8 c2 c6 c0 c9 c6 cf d8 db df e5 e4 e4 df d9 d8 db d1 bb b6 b5 a6 a4 a6 a9 a6 a6 a7 ac aa aa aa a4 a5 ae b4 b2 bc bb c0 c0 c0 ca c3 bf ca c8 c5 c7 c0 c9 bd c5 c5 be ba ba b3 bd b3 b3 b0 ae b0 a3 ae a6 ad af a6 9c a0 9b 9e 9c 93 8a 8c 85 85 86 7d 83 7e 7d 7b 82 78 7d 70 70 7c 75 76 7e 82 8e 95 96 96 9b a4 ab ab b3 af b2 b5 bd b1 b3 b9 b0 b2 b6 b5 b6 a1 ab b0 a4 a6 a4 9a 9c 9a 93 94 96 92 8d 95 8a 8f 85 7d 81 8e 85 89 8e 8c 8d 8a 7a 90 96 a2 98 82 79 6f 74 6d 6f 81 79 5d 41 24 1e 0e 06 08 04 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 01 06 05 03 0f 13 12 11 11 1c 21 25 35 54 5b 70 85 96 94 81 91 96 9d aa a1 90 8b 81 85 88 8c 89 90 8e 94 8d 8b 8b 94 9d 93 97 9e a3 a9 a6 aa b2 b6 b5 b2 aa ae ab b5 b6 c4 c6 cc d2 cf ca d2 d0 cd dc d8 df e9 e6 ea e4 df d9 d9 cb cb c9 bc b5 ad ab b2 a5 ab a4 aa aa 9e a2 a2 a7 a9 b6 b5 b7 bd be c3 c4 c2 c9 c6 ce c9 c4 c5 bf cb cb c3 c1 be bf c0 bc be b3 bd af b3 b6 b1 b0 b0 ae b1 a7 a4 a3 a4 9c 9a 98 95 95 94 92 90 8d 86 86 83 83 74 83 82 74 7a 76 78 74 7d 85 88 95 93 9a a3 a1 af af ad b2 b6 b4 b2 b9 b7 b9 c0 b6 ba bd b9 bb a7 ab 9f a0 a5 a6 a3 9e 9a 9e 95 8c 9a 92 95 8a 8a 8c 8b 85 87 95 90 86 8a 80 84 88 84 94 9e 9b 8b 82 73 72 70 7a 87 92 71 45 30 1b 12 15 0b 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 05 08 04 0d 0c 07 07 11 12 17 21 2a 2e 44 5b 6b 82 86 a0 90 7e 73 72 7d 85 8e 8c 8a 88 84 7d 8a 87 89 90 93 90 95 95 93 98 9b 99 a0 a2 a8 ae b0 b0 bc b4 be b9 bc b0 b8 b9 b8 c5 cb da d2 d5 dc db dd df e0 e7 e8 e7 f1 e7 eb e1 e6 da da d2 cd b8 b6 b4 b5 b8 ad a5 b0 af a1 9f ac a6 aa ae ac b1 b3 b5 b9 c2 c0 c7 c6 c6 c4 ca d2 bd c4 c3 c0 c4 be c5 b9 c4 b6 bd c0 b2 bf b5 b6 b9 af ae bb a8 ac aa a4 a5 a5 a1 9b a0 9c 94 98 97 91 8f 8a 8a 83 82 82 81 80 82 7d 78 76 78 80 82 8b 94 9b a3 a4 ad b5 bd ba b6 b9 c1 c2 bd bd c7 b1 bf bd bb bc b7 a9 a9 ab ac a5 a8 a3 9b 9f 9d 94 9b 9c 96 90 8e 8f 93 89 8e 8a 88 91 87 8a 82 8b 8e 95 a4 99 94 86 7d 73 78 77 92 a9 8e 60 43 22 20 16 12 08 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 05 07 09 0c 09 18 10 25 20 2c 3e 49 5f 79 87 a1 aa a1 71 7d 7c 72 7e 81
 76 84 92 8d 8b 83 85 78 85 9a 97 97 9d 97 98 99 a2 a8 a0 ab a4 ac c2 c0 b7 b8 bb c0 c2 bb c2 bd cc ca cb d4 dd df e6 db eb e6 e0 eb e4 f2 ed ec e7 e9 e4 de db d3 ce c5 be ba b6 b6 b2 b6 a3 a6 a6 ad aa ad af ad b5 b2 b6 bc bf c1 c8 c1 c4 c9 cb cf c9 c6 c7 cb c8 cb c4 c9 c5 bc ba bb b7 be b7 b9 bf be af b0 b7 b2 ac b0 a9 a9 a1 9f 9c 9c 98 a2 92 9a 9d 91 8b 87 8f 86 87 82 77 7e 7c 86 7c 87 89 85 95 98 a1 a9 b2 af b3 bb c1 c1 bf be c6 c3 ba c3 c6 c1 be be b9 b7 b5 ad b3 af b0 af a3 a4 aa a5 9f a0 a0 94 9c 92 92 8c 90 91 92 91 8f 8a 85 89 88 89 96 a0 97 96 8f 87 79 7f 80 90 ae 9e 69 47 37 22 21 0e 0e 0d 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 09 0b 0b 0f 12 1a 23 25 3c 48 5a 77 7f 96 a1 b4 a2 84 69 67 63 70 79 72 7d 80 83 8a 8b 89 82 84 87 82 88 95 9b 9d 9f 9d 9e 9d a6 a5 ad bc b5 bc c5 bd c0 c2 c6 be c3 c1 c3 cc ce d4 db e7 e6 f4 ec e4 ec eb eb ef e3 ed e9 e9 e0 df d8 d3 cb be bb bc b0 b7 b4 b1 b6 ac a6 ae a2 a9 ad a3 b1 af b7 b3 bc bc c0 cc cb cc c6 c7 cb c9 c9 c7 c6 c3 c0 c7 be c0 c1 c3 be b4 bc bd c2 ba b4 b9 b5 b2 b8 ae ab a4 a3 a4 a6 a3 a4 a0 9e 9b 9f 99 9e 98 8e 88 87 8a 7c 82 7e 85 81 8e 8c 8e 99 99 a1 aa b7 b9 bc c5 c8 c2 c4 ba ce c5 c2 c5 c0 c2 c7 bd bf b4 b6 b1 ad b2 b7 b0 ae ac ad ab a0 a0 9e a1 9c 96 9e 94 92 8f 91 93 8f 8c 8a 84 8b 89 97 9a 9f 95 91 85 84 84 82 90 b2 a9 82 5b 3d 26 1d 21 18 11 0c 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 07 09 0b 11 1a 14 1a 2d 31 43 57 6e 84 94 a3 a2 ad a0 85 6e 63 6f 6a 71 7a 77 7e 7c 86 83 89 91 8a 82 7c 95 88 8e 96 95 97 a5 a8 a0 ab a6 ab b6 be bc c0 bd ba c1 c8 c6 c6 ce c8 cf db d6 e6 e1 e4 e9 ee f0 f3 f5 ed eb eb e5 e6 eb de e4 d7 d1 ca bb ab b9 b6 bc b8 b1 b3 a8 ae a7 a9 aa a8 a6 b4 b0 b9 ba ba c5 c1 c6 c6 ca ce d1 c8 c4 c7 c9 c1 c9 c8 c1 c8 be c1 bd bf c8 ba ba b4 c3 ba b9 b7 b6 b9 af a7 af a6 aa a9 a2 9a a6 a2 a4 9e 9c 95 9c 95 90 8c 87 86 8b 82 84 86 89 8e 88 93 a4 a6 ad b0 b8 c0 bd c5 cb c9 d1 d0 cc c9 c5 c3 c7 c9 bf ba ba b2 bc ad af b4 b4 b6 ae b8 b3 9f a7 9d a8 a4 97 9a 9e 95 8f 95 94 92 90 8a 87 8a 86 82 8f 90 94 9c 93 85 86 87 8a b7 b5 93 6c 46 3a 2d 28 1e 12 0d 09 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 07 14 14 1c 1e 28 2c 48 50 5f 68 89 95 97 95 8a 86 79 6b 71 72 6e 6f 71 6d 73
 80 7a 80 89 87 90 8e 84 8c 87 8b 8d 8e 9e a3 a5 b1 a2 a3 af af b0 b9 c1 bd c8 c6 d2 d3 cd cf d0 d2 db e0 e0 c6 e1 e8 e9 f8 f2 f1 f5 f8 ee f5 f4 f1 e8 e2 d9 d5 d2 cb c3 ba b7 c4 bd b9 be b6 b6 aa aa a9 a7 a4 aa ad b9 b6 b6 bd bc c2 ca c9 c5 cc c9 c6 c7 c7 c4 cd ca c1 c6 c6 bd c1 bb c1 c5 c1 c2 bf ba b7 c1 b7 bd b0 b2 b1 b0 b0 ad ae a8 a8 aa a8 a3 a1 a0 a4 94 92 94 9b 97 8c 90 7e 84 90 90 90 96 a3 a3 a4 b0 b4 c2 c3 c9 c9 ca d3 ca cc cf c7 c6 cd c4 c6 c4 c9 c1 b7 c1 b6 bd be c5 bc b6 b1 b5 b1 b0 ad a7 a5 9f a7 a5 a3 a9 95 99 92 93 8a 90 8e 86 8a 8d 91 89 97 8c 8f 91 83 8a aa c5 a6 81 60 42 30 30 2c 1f 17 09 07 07 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 06 05 05 12 10 1a 21 20 2d 3f 50 5d 5f 5f 68 6d 72 6c 6d 6b 67 6e 6e 6b 6a 70 72 76 75 7d 7f 7d 7d 84 8f 87 8c 91 93 95 90 90 90 93 95 a3 ab aa aa b4 ac b5 b0 b4 bd c4 cf cc ca d5 d4 cd d5 d5 d6 e2 e2 ec ec e7 f1 ef f6 f6 f9 f6 f0 f2 e8 e5 eb dd df cb c3 c5 c0 bc c3 c0 bb be bb b4 b9 b7 ae a6 a5 a7 b9 b5 ba bc c2 c0 bf c5 c3 c0 ca c9 c0 cc c8 c5 c8 c6 c8 c9 bf cd c3 c1 c4 bf c2 c0 be ba b9 bf b9 b8 bd b7 ac b5 ab a7 ae ae aa b2 a8 ae a2 a4 ac 9e ac 96 9c 97 90 8f 89 91 94 9b 9d 9b 9e a3 ab b8 be c5 cd d5 ca d3 d0 c8 d0 cc cb c8 cb c6 c9 c7 c8 c6 c7 bb c0 c0 c0 bf b9 ba bc b6 b1 ad ae ab aa a7 a6 a5 9d 9e 8d 9c 8d 94 8d 95 90 87 85 8c 83 82 90 8b 8d 85 88 8b a1 cc b8 9a 6e 56 3f 40 38 25 1f 08 03 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 1a 1e 1e 1f 33 47 54 5a 64 64 65 6a 68 6c 64 62 64 67 68 6e 6c 6b 6b 69 74 77 79 7f 7c 7b 80 84 88 91 94 91 8b 89 92 93 97 9a a0 a5 ac b0 ab ab b1 b4 b7 c0 c5 cb c7 ce d4 d7 d1 db d9 d7 e7 e1 e0 ee f2 f7 ee fc f5 fa f2 f0 ee ef e4 ea de d5 d2 cd c5 c2 c3 b8 c5 c3 c1 bc be b9 b1 b5 ae af a3 af b2 bc b6 bb b7 c6 c6 c0 c4 c0 c2 c3 c3 cc d0 c7 cc cf ca c9 c4 c4 ca c8 bc bd bd be c3 ba c1 b9 ba b9 b7 bb b6 b8 b8 aa b3 a7 b0 af b1 ac af a6 a5 a9 9d 9d 9c 97 97 94 94 94 95 93 9d a3 b2 b5 ba ba c9 c7 d3 dc cd d5 d0 cc ca d0 cc c9 ca cb cb c0 c7 c9 c1 c1 c6 c3 c6 c4 ba bb b6 b9 b4 b5 af a6 af ab a0 9c 98 98 9c 93 99 8c 87 96 87 8f 88 8e 83 83 84 86 87 89 84 95 b7 bf a7 7a 62 5a 46 3e 30 2e 18 16 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0e 0c 0f 1e 1a 25 28 3e 50 5e 5d 68 66 6b 68 6f 6d 6b 64 6a 66 6c 68 65 6e 71 6d 72 73 7c 73
 79 80 83 82 8b 91 8e 96 96 99 93 98 9a a0 a0 9d a4 a0 ab b2 a9 ad ac b4 b9 be c7 d1 d2 d7 db d7 e0 e0 db e0 db e0 f3 f5 f3 f6 f6 f8 f9 f9 fa f4 f2 e4 ea de d6 d1 d3 c2 c0 c8 c2 cc c9 c1 c1 b5 ba b5 b4 b2 ae b1 b5 be bd ba bc c1 c5 c4 bf c9 c2 c5 d1 c6 cc cb c8 ce cb d0 d0 cb c7 c5 ce ca ca c7 c7 bd bb bd b9 bc be be b4 bf b8 b8 b7 b4 b7 b6 b3 b8 b3 b2 af a9 aa a9 a3 aa a6 a6 9d a0 98 a3 a1 a6 af b2 ba bd c5 cd ce cb db d9 db d6 d4 d2 d4 d1 ce ce cd cf cf cb cc c9 c4 c2 c4 c3 c3 bc bf c5 b5 b9 b2 b5 a8 ac ac a0 9e 9b 9b 95 90 93 84 8d 8e 8f 88 90 89 81 8b 84 8b 86 85 80 8f b1 d2 c0 a3 86 6c 5c 4a 38 25 23 14 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 09 1d 16 25 2b 2c 3a 56 6d 6c 67 69 6c 6c 70 67 6a 6a 74 68 6e 6b 72 73 70 74 75 79 7a 7d 7e 7d 87 84 8b 8f 90 94 96 95 9c 95 90 9d a0 a3 9e 9b a7 b0 b4 b8 b2 b4 b6 c6 c1 cc d3 d1 d6 d3 df e8 e1 e5 e4 e7 ef ee ea f3 f0 f4 fe fa fd f1 f5 ec eb e5 e1 e0 cf d0 c6 c4 c6 cb ca c7 c7 c6 c5 c0 b8 b8 b1 b0 b0 b4 b2 c2 c0 bd bf c0 c8 c7 ce c6 cf ca cb d1 cd cc c7 c5 cd cd d0 cd ce d1 cc c5 c7 c9 c4 c1 c1 bb be c3 c0 b2 c1 bf b7 c0 b6 bc be bb b6 b5 b4 b6 b7 b1 ac a8 aa a1 a4 a9 9c a5 a5 a3 b1 b5 af b3 bf ca cd da d4 d6 d0 d8 de db d6 cf d5 da d4 d8 d3 da d7 d0 d2 cd c9 c9 cb c8 c7 c6 be b5 b9 b1 b3 b3 ac a9 9c 9d 9f a5 9e 96 90 8b 98 90 8b 90 8b 8e 8b 90 88 8b 86 86 84 8b a4 c7 c2 af 97 80 74 61 4f 3e 2d 1d 1c 11 08 06 00 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0d 17 16 18 27 2b 3b 49 6f 83 7b 74 68 6a 6f 70 6d 78 73 68 75 72 71 73 6e 7a 77 7d 7f 74 7e 7e 8a 80 90 8e 93 90 90 91 9d 9b 97 9e 9b a0 a3 a8 a8 a9 b2 b0 b8 ba b9 b7 bb c0 cb d0 d2 da d8 de dc da e4 e6 f0 ee f2 f0 f4 f3 fe fd fc f6 fd f2 ec e4 e4 d6 de d2 c8 cb cd ca c7 c6 c3 c6 cc c0 c0 c4 be ba b6 af b4 b6 b7 c2 c3 c2 c4 c0 d0 cd cc db d5 d3 d6 d8 d4 ce d1 d3 cd d1 c4 d6 d0 c7 ce c9 c0 c5 ba c4 c8 c2 c7 c0 be c2 bc c7 c3 bc bc b9 b7 bf ba bb b6 b9 ba b5 af b2 ae ac a1 a6 aa a8 a8 af b4 bc bc c5 cb d4 d7 dc d7 d8 d9 da db d9 d5 d5 ce db d8 d4 d6 d1 d3 d2 c9 cd c8 cb c8 c6 c2 c4 be b6 b9 bc ac ae a9 9d 97 98 a0 94 89 92 90 90 89 8c 85 8b 8f 90 8e 89 7f 7f 86 81 84 93 b1 ce b4 ae 97 84 71 5e 4d 36 2b 1f 17 19 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0e 17 1f 23 34 3c 47 64 8a a6 89 75 76 6e 72 74 75 6f 77 6a 6b 71 77 7b 78 7e 78 7d 77 80 80 81
 8b 8f 89 92 98 98 93 9a 9e a2 a2 a0 a9 a0 ae a7 b0 a7 b5 be bd bc c1 c2 bd c2 cb d3 c6 d0 d2 d8 de e2 eb ea ea e6 ee ed f3 f1 ec f9 f6 f2 f6 ec f1 ec ed dc d0 cf ce cc c6 cc c9 c5 ce ca cf c4 c9 c6 c2 bd c2 c1 bd c2 bb c1 c8 c9 cb d3 db e0 db d9 e3 e4 e2 e3 de dc dc de db d7 d9 d4 d7 d1 cd d0 c6 cf c2 cc ca d1 be c5 b5 c4 c0 c0 c8 c5 c4 c3 c1 c1 ba c1 c1 c3 be b5 b1 b8 b4 b3 aa b3 b6 b3 b9 b5 bf bf bc c7 c9 d7 d7 dc dd db db e2 e4 d9 db d7 d6 db e3 db de d0 d5 cf d2 cf ce d2 d1 c9 c0 c4 b5 b0 b5 b5 b6 b3 a7 9c 96 9e 96 8e 99 93 92 94 8e 8d 8b 84 91 95 86 84 88 78 7d 81 7e 86 aa c5 cb bc a9 90 7e 6a 5e 53 32 2d 29 1d 09 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0a 0f 15 16 27 39 4c 55 6a 84 a9 ad 85 7a 73 75 78 75 74 74 71 72 73 74 81 7d 80 81 82 83 87 8b 87 8a 8b 91 8a 8c 94 9a 9a 9e 9e a5 ab a7 a9 b0 a3 b4 b2 ae b9 c1 be c7 c3 c7 c3 c7 d0 d0 d3 d0 d9 d8 d8 d9 e2 e6 ea eb f4 f0 f4 f1 f6 fb fb f1 f3 f1 f1 e8 e7 df da d5 cc c2 ca ca d2 d8 ce cb d4 ca cc c5 c8 c8 be c6 c2 c2 c9 cd cb d4 d7 dc ed fa ff ff ff ff ff f9 fd ed f0 f2 ee eb e0 de dd dd d4 d9 d1 d4 d4 d0 d2 c9 d0 d1 cb c5 cb c2 c8 cd c7 cb d0 c5 cf cc c4 c9 c9 c1 c2 c4 bd b4 b9 b5 b8 b6 be bd c5 c9 c5 c9 d3 db e4 da de dd e9 de e2 d2 d9 dd db dd dc db dd d8 ce d5 d9 cf d6 d3 cc cc bd c0 b6 bb b5 ae ac a7 a9 a6 9c 9a 9f 91 91 99 8e 97 8c 8e 96 8d 93 89 8a 8c 7f 81 7b 79 7b 7b 91 bf cb c8 ae a2 91 77 6b 59 4d 40 28 10 05 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 09 06 12 1a 1b 30 41 57 6c 85 a7 b1 96 7b 77 76 7b 7c 75 75 74 73 7a 7d 82 81 84 85 85 85 8e 92 86 82 8f 91 92 92 91 94 9e 97 a4 a5 9e a9 a5 a8 ae ac ad b6 b0 bf bc c1 c3 c4 c2 c7 d0 d2 d4 d1 d2 da d6 df e1 e5 e4 e6 f2 ed f3 f9 f0 f2 f4 f6 f7 f5 f4 f2 ed eb e3 dd d9 d0 c9 ce ca cf d2 cf d9 d6 ce d3 c9 c6 c5 c7 c7 c7 c6 c7 c8 cb dd ea fd ff ff ff ff bc ff ff ff ff ff ff ff ff ff ef ee e0 e7 e2 d4 da d3 d1 ce d2 cd cf cd ca d4 c6 d0 ca d1 ce d1 ca d7 cf cd c7 c6 cf cc c7 c8 c6 c4 c4 b8 bc b9 be bb c7 c9 cb cd d4 d4 db e2 db e0 db dd e8 d9 df da df df dd e3 da da d6 d7 d2 d6 ca d4 c6 c9 bc b6 b7 b3 b3 aa aa aa a5 a2 9d 98 94 94 93 9a 90 94 8d 91 89 95 8f 91 85 8a 83 7a 73 74 78 74 7c a7 be be bd af 9a 8f 7c 64 54 48 35 21 12 01 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 10 12 14 20 29 3e 4d 5c 82 9a b9 b5 87 85 82 73 7b 6e 7b 81 74 84 7c 72 80 87 88 8a 89 8e 8d 90 8e 8e 93
 94 95 92 91 a4 99 9e a4 a0 ab ac aa b5 b7 b5 c0 b7 b9 bc b9 c2 cc c7 c1 d0 ca cc d4 cf d0 d9 dc dd e2 e5 e6 e9 e7 ea eb f1 f1 f6 f8 f7 f0 f2 f0 e3 e3 e6 e5 db d0 cd cd c9 cd d7 cf d3 d0 d1 d9 e0 cd d4 d3 d2 cf cd d2 d6 e1 e9 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ea e8 da d9 d7 d4 d5 d7 db d6 df d4 d1 cf d5 d9 d2 d4 d9 dc d1 ce cf d4 d4 d4 d8 d4 c9 ca ce c7 c5 cb c7 c2 c8 c6 cb cd d9 d6 e2 dd e1 e0 e3 e7 eb d9 e6 e2 dd df ea e8 e1 e0 e1 de d6 d1 d8 d9 c5 c9 c3 bf b6 b7 b4 a5 a8 a6 a5 9e 9c a0 95 9b 91 94 8a 91 91 8f 8d 8b 8b 87 87 85 78 74 7e 72 79 75 7b 8d ac ce cc b9 ae 9a 88 6e 5c 4b 32 1c 11 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 10 20 2c 33 4a 5d 76 91 b4 b9 9b 86 79 81 7e 8b 7d 87 7b 80 85 79 7e 82 87 85 88 8a 8d 92 8c 91 84 9b 99 96 93 94 9e 99 a2 97 a7 a4 ac a8 b9 b9 ba bf be b8 bf ba c4 c9 cb c5 cb cf cd d8 d6 d2 cf dc dc dd de ea e7 ee e9 f1 f4 ed f4 ef ed f7 eb ea ef e6 e8 e0 d6 da d6 cf d0 cf d2 d1 d2 db dc d9 d6 d4 d3 d7 d5 d0 d6 d8 e5 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed ea df db db d2 e2 dd dd d6 da d6 df d6 db dc d9 da d5 d5 df de dd db df de e2 d7 cb d0 cd c9 cd cd c5 c4 c2 cb cf cd d8 dd e1 e5 e6 e0 df ed df e2 e8 df e1 e6 e4 e7 e8 d6 d8 db d0 d2 c9 d0 c5 bd be b8 af ab b0 a8 9b a0 9e 9b 9d 94 8e 93 98 97 99 93 98 90 8d 8b 88 7f 81 7b 75 71 76 74 7d 76 7e 95 ab c3 c7 b0 a1 94 7d 65 48 32 1a 12 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 07 15 18 18 2c 44 4d 66 86 a4 b6 a5 92 8e 83 84 81 89 80 7f 86 7a 81 7c 81 8e 82 8c 89 87 8d 8a 97 8f 8e 96 97 91 9a a0 a1 9c a2 a5 a5 a1 aa b2 b1 b9 b7 c5 c0 b6 b5 b8 c1 c6 c1 c0 c2 ce d4 c8 d0 d0 d0 d5 de dd e1 e2 e3 e0 e1 e4 eb eb ed f3 ee eb eb e4 eb e9 e8 dc d7 d2 d3 cf d2 d1 d5 d6 d5 e2 d0 db d6 df d7 de d9 d4 df e6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 e3 e2 e5 df e1 e6 e0 d9 d5 e1 dd dd e4 e7 e0 e3 e6 e4 e9 e4 de e3 e5 e5 dd db d0 cc d2 cc c9 c5 c1 c7 c6 cb cd d4 d9 db e4 e0 dc e6 e4 df df e0 e8 d9 e8 e4 e0 df e0 e1 da d8 d8 d1 ce c8 c1 c5 ba ad a8 aa a5 ad 9d 99 9d 92 99 96 97 95 99 95 90 96 96 93 8b 8d 7d 7d 7f 78 79 72 80 79 78 74 77 7b 98 b4 ba b7 a8 95 82 64 54 2f 2a 0e 00 0d 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 04 06 05 10 1b 1a 21 3b 4e 5f 79 88 9f aa 9c 9b 88 8e 88 81 88 88 80 80 84 8a 88 84 86 7f 8b 8b 89 86 82 92 8f 96 9b
 a0 9e 9b 9e a5 a5 a9 a3 ab ae aa be ba b2 be c4 bf be bf bf c4 c3 be c4 cd cb d0 d0 cd d1 d5 db dc de d5 de e1 e5 ea ee ef ec ed e9 f2 ed e9 e2 e8 e0 df dd da d8 d6 ce cf d1 d6 d4 db da e0 de db e7 dd e2 df e4 e8 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e3 ed ea ec e1 eb dc e2 e5 e5 e8 e6 eb ee ea ee e3 ef f5 ec e9 e8 ea e0 db d6 cb d2 c9 c6 c6 cc cc c7 d3 ce da db d9 d9 e6 dc ea de e3 df e3 e7 df e5 e6 e1 da df d7 df d4 d4 d0 d0 cf c6 bf bf b3 af a6 a1 a5 95 9f 8e 8c 99 96 99 8e 9d 95 a1 99 93 8d 92 83 7b 80 77 6e 72 7a 76 7b 6d 75 6d 7c 89 9d c0 ba a5 93 7a 66 5c 40 34 21 0b 15 05 05 00 06 07 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 07 0a 15 15 21 21 28 40 54 6d 84 81 8a 90 8f 95 8e 87 8c 84 86 87 86 82 88 88 89 8d 8d 87 8f 8c 87 90 93 93 92 9a 8e 97 9f 97 96 a8 a1 a7 b1 b4 a6 b6 b5 b9 b1 bb b6 bc c3 ba ca c8 c4 c8 c8 c7 d1 ce c8 d5 d4 d8 d3 d3 d9 e1 e1 e3 e8 e4 e4 f0 e9 f2 e9 ef ed e1 e6 e6 de e2 e0 d7 d4 d2 cd d4 d2 d2 da d8 de e2 dc e8 e0 ea e2 e5 ea f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef f2 ee ed e6 ee e3 e9 e9 e6 e6 ed f5 ff fe fc ef ef ed e7 ea e6 dc db de d0 ca d0 d2 d4 cc cc ca cf cf d0 db df e4 e1 df e0 e1 df e0 d9 e5 e0 de e8 e3 e6 e8 db df d4 d4 d0 d5 d2 c0 c5 b9 b6 b0 a3 aa ac a4 a1 9b 9a 8e 97 92 9c a4 91 9b 9b 91 8f 88 88 84 82 7e 86 70 75 7c 76 71 7d 72 7c 6f 74 8e a2 af a4 86 7a 76 70 5d 48 2c 15 0f 09 10 05 06 05 03 0a 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 06 17 1b 1b 28 3c 50 5e 71 6e 72 6c 7a 82 91 8e 8a 87 89 79 80 80 8a 90 87 7f 88 8e 8b 8b 89 87 89 90 8d 9a 9a 95 9c 98 9a 9b a7 aa a9 b2 b0 ab ae b5 b7 bb b8 bb b7 c5 c0 c2 c7 c6 c0 c6 c9 c5 cb d4 d8 d5 ce da d7 d8 db dc da e2 e1 e0 e4 ea f2 ed ee eb e3 e4 e6 e4 e6 db d8 dc d0 d3 c9 cd d4 d4 d8 db d7 de d8 db e5 e8 f0 e6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 f3 f0 f3 ec f0 ed ef f0 fb f4 f5 fe f6 ff fd f0 f6 e8 e4 e7 dd d7 dc d2 cd d0 d6 ca ce d2 c9 cb cc d5 ca d7 df d9 dc d9 e2 da e5 e5 df eb e3 dd e6 e5 e7 e1 dd de d6 d5 d4 d1 c5 c4 c6 bd b2 a8 a6 a3 9c 9d 9e 98 9f 97 98 92 98 92 9a 96 8d 86 81 7f 82 7c 81 76 75 73 75 80 81 75 72 74 77 6d 6f 85 84 98 8a 7f 77 72 78 65 4e 3a 28 17 11 0b 0b 0a 05 03 00 06 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0b 17 1a 25 2a 2c 3b 51 61 71 69 6a 6f 70 7a 7d 8a 88 84 80 87 7b 81 8c 8d 8d 87 80 89 87 8f 8c 91 90 93 93 93 9e 94
 9f 9a 9f a6 a3 a7 a6 ac a7 b1 b3 ba bc bb c2 ba c6 c2 ba c9 c6 c4 d1 c7 d0 d1 d0 cd d6 d3 da e3 d9 da e0 e0 e4 e1 e1 e4 e5 e3 eb e6 e5 e1 e3 df e5 e4 d8 df d3 d4 d5 cd cf d8 d8 cd db da db e1 e3 e7 e7 e7 f2 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f4 f0 f4 f3 f3 fa f9 fc fd ff ff ff ff fe ff f3 ef e6 e5 df e1 d4 e4 d8 d0 cf ca d1 cf c7 c6 c8 ca db d0 d2 d8 dc e0 e3 e7 e0 e9 de e2 e6 e5 e3 e4 ea e8 df dc e2 da d4 d4 cd c2 c0 c2 b5 b5 ac a6 a2 a6 a1 9e 9c 9b 90 96 95 92 97 90 88 8e 8a 81 80 81 78 7d 7c 7d 7d 7d 7a 78 75 6a 70 73 76 75 75 84 7e 83 77 7d 8c 84 76 62 44 2c 1d 12 0c 00 0b 05 09 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 20 22 2a 32 3b 41 51 57 5a 63 68 63 65 66 74 84 86 84 88 81 85 82 84 84 90 8c 84 83 8e 8c 8e 8a 8f 8a 8a 8e 96 9f 9f 9c 9c 9f aa af a6 ab b2 b4 b2 ad b5 ba bd c3 bb c3 c5 cb c7 c6 c6 cc ca ce d5 ce d2 d3 d8 de da de e0 e1 e2 df e0 e9 ea ec e6 e0 e8 ea e2 ec e0 dd de dc d7 d8 d5 d4 d0 d6 d1 d7 d7 d1 d7 d5 e2 e7 ed ed ee ef fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff ff ff ff ff ff ff ff ff ff f7 f6 f6 e8 ec de dc de cf d8 d3 ce cc ce cc d1 d6 ca d2 cb d5 d4 d7 dc dd e6 e5 dc e9 e5 eb e3 de e4 e3 e7 e9 ef de e1 e2 d4 ce d0 c4 c5 ba b2 ad ab af a5 a8 9e 9e 9b 99 94 98 94 91 94 95 95 88 8e 86 86 80 81 7c 7c 7e 7a 77 80 80 7c 72 76 6f 79 73 7c 73 80 85 70 78 72 89 95 85 73 58 39 22 1a 15 13 06 10 04 03 06 06 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0d 16 1f 29 31 3e 4d 5b 60 61 5b 5e 63 62 66 66 71 76 81 83 7d 82 80 84 7f 81 8e 8a 8e 8c 86 86 90 86 8e 92 94 94 91 90 94 a5 9a a3 a4 b0 a1 b1 b1 b3 bd be bb bd b9 ba c7 c4 c7 c8 c3 ca c9 cd d0 da d8 d0 db d5 d8 dc e0 e0 e1 e3 e8 e5 e8 e9 de e5 e6 f0 e4 df e7 e3 df e3 db dd d0 d1 cf d0 c8 d2 d2 d6 d4 dc df e2 e3 e9 e2 e7 ed f2 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 ec eb e0 d7 d6 d3 da d4 d4 cf d1 ca d4 cb d4 cb d1 d2 d4 d6 d7 d6 d9 da df e0 e6 e5 e4 ea e4 e5 e5 e0 e6 e4 e4 dd da da d7 ce d0 bf c8 b7 b1 b6 b1 a8 a5 a4 a0 9c 9e 9b 9e 9c 95 92 8f 8e 90 8e 8b 84 86 82 80 80 79 7e 7f 7d 7a 6c 71 78 75 73 76 6d 72 70 80 73 73 71 70 86 94 88 7a 60 47 31 25 18 12 0e 08 10 01 07 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 07 1d 2c 2c 2e 35 36 4c 63 64 55 5c 5f 5f 69 6e 72 75 72 79 83 86 88 80 81 80 7e 82 83 86 90 8d 97 94 95 8f 99 93 8f 99 99 94
 97 9c a1 a5 a1 b3 a7 b3 b8 b9 b7 bd ba be c2 c1 be bf c6 ca d1 cf cd cf d4 d6 cf d7 d8 d3 d6 e2 e2 e1 dd e0 e5 e6 e6 e4 e9 e7 e7 eb e2 e9 e6 d8 df dd e0 d3 ce cb be c8 d5 cd d6 cf d4 d6 e2 db df e0 e9 f2 f0 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ed f0 e3 dc db da d3 d8 d8 c6 ce d3 cc ce d1 cd d6 cf d3 cd d1 d5 de da df db e0 e6 e2 e5 e1 e9 e8 e3 e8 e6 e0 e2 e0 df d9 d6 cc cb c2 c2 bb b5 b4 b7 b0 a7 a0 aa 9b a0 94 91 94 8e 96 8d 8f 8c 91 8d 89 79 7e 80 81 85 82 85 80 7c 7c 7c 74 79 74 74 6d 75 72 79 78 73 68 6d 64 73 85 91 84 6a 50 37 30 1f 16 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 03 0f 0d 1f 2e 32 3f 37 42 4a 5a 63 5d 61 5f 59 5f 68 73 76 77 74 77 7f 8b 86 7f 7c 7d 85 86 8c 85 8e 8f 99 98 93 96 95 94 98 9a 97 98 9a a6 9c ae a6 ad b2 bc b6 bc bd c2 bb b8 c5 c4 ca c5 cb c5 cf d1 d9 ce d2 d4 dc de e0 de e4 e4 df e9 eb ef ee e0 ef f0 ef ee f0 e7 e5 d6 de dd dd d7 d7 d2 cb cb d0 ca d2 d7 da d9 d9 e6 e3 e5 e6 ea f1 f0 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 ff f7 f7 f1 f1 e4 e5 dc d9 d5 ce d5 d4 d0 d5 d0 cc d4 d2 d1 dc d0 d7 d7 dd db dc e2 de da e4 dc e4 e7 dc ef e1 e1 e8 e7 e3 e3 e4 da da d8 c6 cc be b9 b9 b7 b1 b4 a3 a8 a1 a7 9b 9f 9a 9c 97 98 97 96 89 8a 8f 82 8a 84 88 81 75 87 82 88 83 7b 7a 75 75 7c 6f 6e 76 76 70 7f 7d 73 6e 65 65 6b 84 8e 87 75 5b 4a 2d 1d 1e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 0b 14 0f 20 2e 38 36 45 4d 45 45 50 5a 58 64 67 63 68 65 6d 6d 73 7b 75 77 81 87 82 7b 76 73 7a 87 87 8b 96 92 95 8f 93 96 8c 8f 9a 9c 9e 9a a2 a9 ae a6 b6 b2 b5 c2 b5 bc c0 c3 c4 c5 ca cf cb d0 c9 ce cd d4 d7 d9 d9 e0 e6 e1 e6 e9 f2 e8 e8 eb ef f2 e9 e9 ea ee f0 f1 e1 e1 e2 df e2 da d5 d9 d2 d2 d1 cf cc d0 d7 d3 da df dd db e8 e7 ea e7 f1 f3 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff f5 f9 f1 f6 f4 e6 e5 e0 db db d3 d3 d0 ce d3 d2 d2 cf ce dc d3 d5 d4 db d2 d3 d5 db d4 da d9 df e4 e3 e3 db db e2 ee db e3 e4 e0 e2 e4 de d9 da cc ca c7 be ba b7 bb ae b3 a8 a1 9e 99 97 9d 96 95 97 8d 96 8a 8b 90 8d 8b 8d 7d 8c 8f 84 87 80 7e 7b 7a 7e 76 7b 6d 7e 74 72 76 79 75 71 73 6d 6d 65 73 7f 95 96 75 6c 52 3c 2b 18 0c 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 17 22 23 2d 3c 4b 4d 59 50 54 52 56 5f 5c 65 5f 64 6c 6d 71 73 72 78 7d 7c 79 84 84 75 7a 7f 7a 89 81 92 90 8d 91 8d 95 97 94 90 9a
 98 99 a1 a1 aa ac aa b3 b7 b3 ba bd be c6 c5 c4 c9 c4 d1 cc cf d7 d4 d6 da e2 da d5 e2 e5 de e3 e8 e3 ee e8 ec ee ef eb f0 ed f0 f0 e9 e2 e2 e4 d8 d9 d6 d3 da d3 cd c1 cf cd d7 d5 df e0 e2 e7 e9 ec ed ee e5 ef fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff fe fa fa fc f4 f1 f1 ea e4 db df db d8 d3 d4 cc cd d2 cb d0 c7 cc ce cf d9 d1 d2 d8 d5 d1 d1 d9 d2 db d6 dd dc e1 e3 e3 e5 d9 e6 dd df e5 d8 e3 df d6 d6 cf c6 c8 bf be b8 b3 b5 a6 a6 a7 a4 9d 9e 9e 9d 95 91 91 8e 93 98 8c 93 90 8a 86 8d 86 85 80 7f 79 76 79 78 6f 72 79 73 71 74 72 75 71 6f 6f 6b 6e 66 66 6b 7f 85 8f 87 6e 52 39 23 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 1c 2b 2b 34 49 4a 59 66 5a 54 56 5e 60 63 69 6a 62 66 6c 71 70 78 74 72 7d 80 7e 81 80 7d 80 84 88 8a 92 87 91 91 95 94 96 90 96 95 9b a0 9a a6 ac a7 ad b1 b3 b6 bd bf c2 c1 c3 cf cd cb d6 d5 d0 dc dd d8 e1 d6 e1 da e4 e4 e6 e8 f0 eb ef f4 ea f1 f5 ef fb f0 f1 ef ea ea df e2 e2 d8 d2 d1 d0 d6 cc d0 d5 ca d6 dc dc df eb ec ee e7 f2 f5 f4 f3 f8 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fc f9 f4 f5 ec f1 e7 e2 e7 db d6 d8 d6 d3 d0 d3 cd ca cb d6 ce cc d0 d6 db cf ce dd d6 d9 d7 d9 e0 db d7 dd e1 e2 dc e0 e1 df dd e6 e4 e5 e2 e1 d7 d4 db d1 c7 c9 bf b9 b1 ae b3 a9 ab a7 a4 9e a3 95 9e 98 9b 9c 96 9d 90 8e 8a 92 8e 90 90 8c 87 83 7d 7d 76 78 77 70 72 78 78 74 6f 70 6f 6f 75 7b 6b 70 70 6d 6b 77 85 90 83 6d 5e 42 28 1d 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 00 0a 19 21 2c 2e 42 4e 58 67 6b 62 5f 56 6a 61 61 70 69 66 6b 6e 69 77 75 6f 77 75 7a 7a 7c 7e 7a 81 7b 83 89 85 8a 92 93 95 9e 92 94 93 95 9e 9f 9d a3 a4 aa ab a5 af b7 b7 bd c1 cb c7 d1 cc c5 d5 d5 d0 d1 d9 d6 e2 e2 dd e4 e4 e4 ec eb eb f4 f1 f7 e9 f1 f7 ed f5 f8 f9 f7 f2 ed f1 ea e6 df e0 d9 d5 d1 d7 d3 d7 dd dd e2 e3 ea ea f2 f4 ff fe f8 fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb fa fa f6 ea e6 e8 e3 db e4 d1 d3 d6 cc d3 d0 d4 d7 d3 ce cb d1 d3 cd ce cb d4 d0 d6 d6 d3 d8 d6 de df dd e0 e0 e3 e3 e0 e1 e2 ea e4 e2 e5 e1 df e0 d2 d5 c7 c4 c4 ba b6 b5 b1 b1 a7 aa b0 9f 9c 9f a1 a1 99 97 9b 9a 9b 9d 97 94 90 8e 8e 8a 88 89 88 77 7e 7f 7b 7d 7e 6e 75 79 76 70 73 6f 6f 6d 6a 6f 6a 6a 64 6e 6b 76 8c 82 71 5e 4b 32 22 0d 06 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 0a 18 1a 2d 31 4b 4d 60 69 78 72 5e 61 5b 67 65 60 63 68 70 67 6b 6d 6e 72 6e 79 76 81 7d 76 7f 84 7d 86 82 83 8f 94 8d 93 99 98 99 97 98
 a5 9a a1 9b 9d a8 a5 ae b4 b7 bc c0 c7 c3 c9 d0 cc d0 d4 d2 d1 db d9 dd da e0 e6 e4 e1 ec ed ec ee f1 f5 f2 f3 f1 f8 f3 fc f1 ee f6 ee f0 ea ed e1 e6 e3 e1 de d9 dc ca dc e0 d9 e5 e1 ee f8 f6 f7 f2 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fe fb f7 ef ea e3 dd db d8 dd dc d5 d0 d2 c8 d1 cd cb ce d4 ce cb d4 d0 cf d0 d4 d9 d6 d9 d6 da da db da db d9 e1 e3 e1 de e7 e5 e2 de e2 de d4 d9 d8 cd d7 cb bd c0 b9 b5 ad b1 b3 a5 a6 a4 9e a0 9a 9d a6 a2 a0 9e 92 94 9a 91 98 8f 91 92 84 8b 7a 81 7f 7e 7d 6e 7a 7a 75 6d 78 71 6c 65 67 69 6f 74 74 6b 6c 65 59 5f 74 84 87 70 62 47 2d 23 0c 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 15 14 27 35 37 4b 58 62 80 84 72 63 63 60 6b 6b 68 6d 71 70 6b 6d 70 70 78 72 78 79 76 7e 78 7a 7d 78 7d 80 7f 86 90 8e 94 9f 95 9f a3 9e a0 9f a3 a2 a4 a5 ae af b3 b1 bb c1 bd c4 c4 ce d8 cd d5 d2 d2 dc e2 df e0 e0 e3 ea f1 ef ee eb f4 f9 f3 fa f4 f0 f4 ef f5 f3 ee f9 f1 f4 f0 e7 ea ee e9 e5 d8 d8 d7 d9 d6 df e6 e8 f2 f4 ec f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f1 e6 e0 dc d7 e4 da da d9 d8 d6 db d5 da d8 d4 da d4 d2 d1 cf d9 d1 d5 d4 d9 d2 df e3 de de e0 d8 de e4 de e7 db d6 e6 e9 de e8 db db d3 da d8 ca ca c2 b6 b8 b4 b2 ae af 9e a3 a8 9e a5 a4 9d a2 9a 9f 9c 97 99 94 93 92 8e 89 8c 84 7f 85 7a 81 78 73 7e 74 75 72 78 7a 6b 71 6c 68 6e 72 6c 75 68 64 5d 5a 60 6f 7f 85 78 5e 4b 30 24 0d 0c 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 0e 24 2c 31 46 4e 60 6d 85 84 73 64 61 69 66 6c 6f 69 6e 6d 6e 6c 74 75 75 6d 76 79 78 78 7c 80 81 86 83 86 7a 7f 80 88 8f 96 9a 9b 9b 9e a7 a0 a5 a2 a6 a4 aa af b3 b5 b6 bf c0 cb c9 c8 cc cb d2 d5 d4 d9 dd de d9 e0 ea dd e9 f0 e5 fa f9 f4 f6 fc f8 f8 f7 f6 fb f8 fd f9 f1 f1 ed f5 ec e0 e6 dd e2 e1 dc d2 df e0 e8 e7 f2 f4 f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f4 eb e5 e4 e0 db e2 d6 da e4 de db d9 dc df d5 d7 d3 d5 dc d9 dd df e3 d3 e0 d6 cf d9 dd dd e5 e1 e3 e4 e6 e1 e2 e6 e2 e8 df df dd dc d7 d7 d0 cb c9 c2 bf b9 b0 b4 aa b1 b3 b0 b5 a6 a0 a0 a7 9c a7 a0 9b 98 9d 93 98 8c 8e 89 8b 83 81 82 73 78 7d 74 78 80 75 75 75 72 6c 69 6a 68 6e 6d 6b 63 64 65 58 58 60 6f 7f 85 7d 6a 4e 3c 24 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0f 07 16 22 46 41 53 67 71 82 83 70 68 5f 64 68 66 6e 65 69 67 67 70 73 72 71 74 6e 72 7b 79 7f 88 7e 83 84 84 82 7f 7f 89 8d 8f 8f 8d 99 8f
 a3 a0 9a a2 a6 a6 ae ad ac b4 b2 b2 b9 bf c2 c4 d1 cf cc ce db d4 df dc e8 e9 e0 e6 e7 e7 ea eb ea ec f2 ff fb f9 fc f6 f5 f8 f6 ff f5 ed f2 f1 eb ed ef e1 dc de da d8 dd e1 e5 ef eb f7 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f2 e7 e9 e2 e1 e0 e2 e6 e2 e2 de da e0 d7 e5 d7 d6 e0 dc d7 db dc da de dd df df d9 dc e0 df e4 e4 e4 de e2 e0 e0 ed e2 e7 dc db dd d9 d6 d9 ca ca c6 c2 c1 ba b3 b3 b2 ad af a4 a4 a2 a0 a5 92 9a 96 9d 9a 93 94 8e 86 87 8c 8c 87 84 7c 7e 7b 7a 7c 7e 76 70 6f 74 6e 6f 6b 69 65 60 5f 68 5c 60 5e 5a 58 58 5f 66 83 85 7d 6a 54 39 29 13 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0d 14 26 3f 48 5e 66 7f 81 7d 69 6a 67 6e 69 63 67 6c 6b 6e 6d 6b 6c 72 73 75 71 7b 79 7c 77 84 80 84 7b 80 7f 80 83 84 88 8b 8d 93 a3 9d a0 9c 9e 9c a5 a3 a3 a8 ae ac ad be bb bb c3 c9 cd d2 c7 d3 ca d7 df dd e6 e4 de e3 ec ec f0 ec f6 f1 f8 f7 fd f4 fb fa f6 f6 fa f3 f9 f9 ef f3 e9 e0 e9 e2 de e0 e3 de df e3 e5 eb f0 fb ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 f4 f6 eb ee ea e6 f5 ea ef ec ee e8 e3 e6 de e4 e5 e3 e4 df dc e2 de db da ea e4 e4 dd df e0 df e8 e9 e4 ea e3 e0 dd dc e6 dc d9 d7 d8 d2 ce c7 cd c5 c0 c2 bd c4 b4 bb b3 aa a9 a5 a2 a1 a1 a0 a4 90 94 92 8d 8f 86 8c 8c 89 84 86 8b 81 79 7e 76 79 7a 77 6d 76 71 78 6c 6b 63 67 5d 63 62 60 62 63 57 54 5b 56 6d 84 89 7b 67 55 39 28 16 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 13 18 1b 3d 4c 60 70 72 86 70 63 6b 6c 6a 62 69 68 64 69 6f 67 6f 6f 70 72 6a 6d 72 73 81 86 84 8a 8a 87 84 8c 85 80 84 8d 8e 8b 99 96 94 97 9b a3 a2 a7 a6 ac b3 af af b7 b7 b9 ba bf c3 c6 d0 d1 d5 d6 d8 e1 db e1 de e4 e8 ee eb ec f6 ee f7 f6 f5 fe f1 f5 f8 ff fb fc ff fb f7 f2 ee f2 e8 e5 e7 e6 e3 df df e7 e2 e7 eb eb f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 f1 fa f4 ee f2 f2 f8 f4 f4 f6 f5 ea ee ed e7 e6 e6 ea e7 e9 e3 e0 e1 e3 e9 e6 e8 de e7 e1 e7 ea e4 ec e4 e4 eb e1 db e7 ea dd d8 de d6 d1 c7 c5 c2 c5 c3 bb bd ba b9 b3 ad af af aa 9c a6 9b 9c 9a 9e 9a 93 97 89 87 8a 8b 85 87 81 7b 7e 81 78 77 74 7e 77 76 73 76 72 6e 6f 6b 6a 64 5f 65 64 6a 59 56 55 59 61 66 80 8b 7e 6f 53 3e 27 17 06 05 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 14 1f 2e 44 62 75 7e 76 68 62 6d 63 69 6e 6b 65 63 6b 64 68 62 68 6e 70 6a 73 71 76 82 83 80 8a 8a 7e 80 89 82 85 88 88 91 92 90 9a 9a
 a2 9d 9e a5 a6 a6 a5 ac ad b4 b6 c0 b8 c1 bf c5 cb c5 c9 d0 d7 d4 db e1 e0 d9 e4 e9 e8 ea f3 e7 f1 ef ee fb f7 f2 f2 f6 f6 f5 fb f5 f1 f1 f1 ef e9 ea e4 e4 e3 e5 e3 e2 e3 df ec f5 f5 f8 f9 fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 ec f4 f6 f9 fa f8 ff ff ff f8 f6 f1 f6 f4 f3 ef ec ec e5 e8 f2 e9 e9 e7 e0 ef f0 f2 e3 e8 f0 e5 ed dc e3 e6 e7 e3 e7 e3 e4 e5 dc db d6 d8 d5 ca c9 c8 c4 c2 bc b9 b9 b5 b3 ac a6 a6 a0 9a 9a 9f 9f 92 95 94 90 92 83 8c 83 86 7e 85 87 7b 80 76 7a 7b 80 77 79 73 71 6f 6d 6e 6c 64 6b 62 62 64 61 5d 55 66 57 53 61 69 82 8c 7a 6f 54 3e 2c 0e 0f 07 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 0b 19 1c 34 41 58 72 71 7b 6b 5d 66 5f 64 6b 60 65 67 67 6d 6b 6a 71 6b 6b 72 70 72 79 7c 85 88 88 8a 8e 87 89 84 86 85 8a 9b 8b 93 99 94 9e 9c 9f a3 a9 a7 b2 b4 b6 af b9 b4 bf b8 c0 c8 c4 c6 c9 d0 d7 d3 d6 d0 e0 e1 d9 e3 e0 e4 e5 ee f1 ef f1 f4 f3 ee ed fa f9 f4 f7 f9 f0 f2 f1 ec e8 e8 e2 eb e3 df e6 e1 e5 df ef f1 f3 f1 fb f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ed f5 f9 f7 fb ff ff ff ff ff ff fc f8 f1 fa f7 f2 f5 ee f5 ec f2 ea ea e9 f0 ef ea e8 ec eb ed eb f1 ec e3 ec e5 de e0 e6 e6 e5 d8 df cc cf d2 c7 c7 bf c5 be be bb bb b6 ad ad 9f a5 a4 a4 a1 a3 9c 91 a0 8b 94 86 8c 8c 87 8f 82 81 81 81 7f 7c 75 78 6f 76 79 72 6f 74 75 64 63 62 5f 5e 64 5f 5e 5d 5d 59 54 5e 5f 6d 83 81 7b 73 56 48 2f 19 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 06 15 1c 28 47 59 6c 80 7b 66 64 60 60 68 6c 63 68 64 64 67 6a 62 6d 6f 70 70 70 74 78 7d 7c 82 88 8b 8a 80 85 82 86 84 86 93 8c 8b 94 99 9a 9c a9 ac a4 aa a7 b5 be b0 b5 b5 b7 b4 c2 c7 ce c8 c9 cf d2 ce d5 da d8 dd df de e3 e4 e7 e8 f0 ed ee f2 f7 ef f7 f2 f6 f5 fa ec f1 ea eb eb e8 e6 e4 e3 e1 e7 e9 e4 e5 e0 e8 eb ec f1 f2 f5 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 fc f9 fe fb ff ff ff ff ff fb fd f8 ff f6 f5 f7 ed ef f0 f5 f3 f3 f1 ef ed ea ec ea f4 ee e4 e7 e7 e6 df df e4 d7 da dd d6 e4 d4 cf d4 d2 cb c4 c7 c4 bc be bb b3 ba b5 b3 ae a4 ac a2 9f 9d 92 95 97 90 97 99 88 96 85 85 88 8b 8a 84 76 7f 7c 7e 7d 74 78 79 77 71 73 72 73 66 66 67 5b 6a 62 60 63 58 63 5d 57 64 6e 82 86 7f 6d 5a 42 30 15 0c 08 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 09 17 1e 32 3e 49 6d 7e 7e 7d 69 62 62 61 63 63 68 64 64 6a 69 6d 70 6f 6d 70 72 7a 7a 7e 84 80 82 86 84 8b 88 84 85 8e 87 90 8a 91 90 9b
 99 97 9e a4 a3 ad b1 a9 b2 b1 b7 b5 bb b9 b9 c0 bd be cf d0 ce cd cd cf d7 d8 e0 d9 e1 e2 d5 e4 ec e9 e3 f0 e6 ed eb ef fa ee f4 eb ed df ee ee e9 e9 e8 e3 e3 df e1 e6 e2 e4 e1 e3 e6 e9 ef eb f1 ee f0 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 f4 f9 ff fe fe ff ff ff fa ff fa f9 ff f8 f2 f2 f2 e9 ed ee ec ec e9 f0 f0 ec e7 ea e9 e8 e4 e7 e4 e0 dd e0 dc de df dc d8 d9 db ce c3 ca c4 c5 c5 be b5 c0 ae b3 ad b3 b8 a9 a1 9d 9b 9e 94 8f 94 91 92 90 8f 87 89 86 83 81 87 7a 80 7a 7a 78 7f 77 75 7e 73 6f 6f 67 69 67 68 66 60 65 64 5e 54 5c 5a 53 52 5a 65 8b 82 7e 70 54 3f 29 17 06 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0e 1b 1e 2f 3e 57 69 7c 85 80 67 5f 65 65 64 69 66 65 66 66 65 65 70 71 68 72 73 70 77 7d 7f 7f 89 85 7f 87 87 87 86 81 81 87 90 83 8e 95 97 95 a0 a0 a2 a5 b0 a4 ab a7 b4 b5 b1 ba be bd bf c0 c7 cb cc c8 cd cf d6 c7 d3 d8 dc d6 dc e5 dc e3 e0 ed eb ec e8 ef ed e1 e7 e2 ef e4 e6 e1 ec e5 e2 e1 da de dd de dd df e1 e6 e0 ec e7 e6 e3 e8 f1 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fb fc fd ff fc ff ff ff ff ff fa f6 f3 ea f6 eb ec ef eb ec f2 e3 e8 e4 e3 e6 e7 e8 e4 e1 e1 dc dd e1 d8 de d9 d9 d6 da db cf ce d1 c7 c4 c4 c1 b7 b5 bd b5 b8 ae ad b1 ad a1 a7 a4 9a 95 94 90 90 8c 8b 85 8a 8d 83 82 7f 83 7d 82 7e 79 71 76 78 71 77 71 64 6a 68 74 68 58 65 5f 62 64 57 59 5c 4e 5d 59 58 60 6b 84 88 77 6e 58 33 30 14 0b 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0f 10 19 2e 36 42 56 60 7a 8e 82 74 65 63 68 60 65 63 69 69 6a 66 6b 64 73 73 75 78 7a 7a 7c 80 80 83 88 8d 86 86 86 8c 87 84 84 8b 8d 97 9e 9b 9b 99 a3 a7 a5 9d a8 a7 ae b1 b5 b3 b4 b9 bd c5 c4 b9 c2 c4 ca cb cb d3 d2 ce d5 d5 cf db e1 e0 e2 e5 eb e7 e2 e9 e6 f0 e6 e6 db e9 ed e2 e6 e9 df e3 e1 e0 da d9 e4 d5 dd da d5 d9 e1 e2 e4 ec eb f1 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 fa fc fd fc ff fa ff f4 f3 fb f2 e7 e9 e9 ea e8 e6 e2 ee dd df e6 e5 e3 de e6 d8 db df de de da dc d4 d7 d7 cb d1 ce cc ce cd c8 cb bc bb c0 c1 bc b9 ba b3 b0 aa ab b1 a5 a5 9a 9e 99 9e 9c 8c 90 88 8e 87 8b 87 88 85 85 6d 7e 76 76 7b 77 73 75 74 71 71 67 68 6a 65 60 65 69 66 66 5a 58 5f 5f 59 56 52 59 67 7d 7c 7c 6d 5b 4b 2d 12 08 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 11 13 1b 30 3a 49 56 66 73 85 91 81 76 66 67 64 68 69 64 62 6b 64 6f 74 71 74 77 75 7a 77 80 84 7e 86 81 88 85 7f 89 8c 82 88 94 8d 92 92 99
 9a 9d a2 a0 a6 a1 a1 a4 ad b0 b1 af b2 b3 b4 b8 b7 bc be c4 c3 c4 c9 c7 c9 d0 cb ca d3 d0 d5 d7 dd e0 e1 e4 db e0 e3 db ea e1 e5 e5 e0 e1 e4 d9 e6 d8 e1 e7 dc de de d7 dc df d7 da db d9 dc dd e0 e9 f9 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f5 f3 f1 f1 f8 f3 f8 f2 f1 f3 ea ee ee e6 f0 e4 e4 e0 e1 e3 dd de db e2 d3 dc d7 d9 da dd d9 db d9 da d1 c8 ce c1 cc d1 ce c3 c9 c5 c6 bb c6 b9 b9 b4 b7 ae b5 b3 a8 b3 a9 a3 a6 9e 95 98 90 8d 8d 94 8b 84 85 8b 88 86 84 87 7f 82 76 7b 76 77 79 6e 75 75 71 72 6c 68 6b 62 62 67 63 60 5e 67 5c 54 57 54 5c 5d 68 82 7e 74 6f 5e 41 34 14 0a 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 13 1c 28 31 46 59 6b 79 93 93 89 6b 67 61 5c 6b 6a 66 6a 60 64 65 72 6f 76 81 74 74 79 76 7f 79 78 84 7e 80 8a 85 87 81 7b 86 86 8d 92 94 91 92 95 9c 9e 9f a1 a0 96 9f 9f ad a2 ad b7 b1 b5 b6 b5 be be be c2 c4 c8 c2 ce ce d0 d3 d6 d2 e1 d3 d6 d5 d6 d7 dd e2 de e5 e0 df e0 e8 db e4 e4 e4 d9 e0 db e0 d4 de d8 d2 d3 d9 d3 e7 da e1 e6 e3 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ee e9 ed f2 f4 ea ed ec e9 ec eb eb e3 e5 df df de dc e0 df d4 d6 d8 d6 d8 d8 cf d4 d5 d5 d9 c9 d1 cb d3 cd c5 be c4 c2 c4 c4 bf c8 b6 b6 b4 bc ba b2 af a5 ab af ac ae a6 a3 a7 94 94 8b 92 90 8c 90 87 8d 85 7b 84 7a 7e 82 83 7f 7e 7b 77 78 70 69 74 6b 72 66 71 69 6c 5f 63 5e 5f 69 5e 62 57 56 57 54 4f 4c 72 7c 89 7f 6d 57 3d 2a 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 18 15 23 36 44 57 5b 6f 7d 86 91 8d 7e 69 6f 63 6c 6d 69 63 66 6a 6e 6e 7b 71 76 75 7e 7c 82 7b 80 80 80 80 7c 80 7e 8b 85 81 8b 85 90 8f 8e 9b 99 92 9a 9b 9d 9e a0 9e a6 a0 a5 a7 a8 af ae b8 b6 ae ba b9 b5 be c0 c7 c5 c1 cc ce d0 d0 d2 d6 cd d4 d5 da d2 db da db e5 d6 dc de da e9 e6 e2 e9 e2 e3 dc dd d7 d7 d2 d4 d9 cc d2 d7 d6 d5 de e0 e7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f4 ef e4 ea e8 eb ea e9 e9 de e3 de df dc e3 e0 dc df d6 d0 e0 d0 d4 d4 d6 da ca d0 d2 cb cb cc cf cd c7 ca c2 c2 c0 c2 cf c2 bc c0 b3 b6 ba bc b3 b7 b5 b0 ae ac ac a5 a1 9b 9e 9b 95 92 91 91 88 86 86 86 8a 85 87 7d 7d 7c 7d 80 7c 78 74 74 73 70 6e 75 73 6e 74 6d 65 60 64 64 63 5f 5c 5e 58 5b 5c 54 5a 5b 68 7a 83 7b 68 59 3a 29 0f 05 04 08 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 19 1b 2d 31 40 56 61 6b 7c 8c 9b 94 8b 67 65 6e 65 65 66 63 70 68 6d 6e 70 7c 71 73 7e 85 82 89 80 7f 84 7c 7d 7f 82 87 80 89 89 80 8c 93 8d
 99 9a 98 97 9d 99 9a 99 97 a6 98 9e a6 ae ab b0 ab b3 ad b5 b4 bb be be c5 bd c1 c5 c2 c1 cd d2 c8 d1 ce d4 d5 d4 d2 d6 e2 d6 e2 e1 e0 e4 e1 e3 e8 e9 de dc df da d2 d8 d2 ce d3 ca d2 d6 d4 d9 d6 e0 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed e4 dd df e3 e7 e6 e4 da e4 dd e3 e3 e0 db e4 d8 e0 da d7 d5 d9 d0 d3 d3 ce ca c5 d1 ca c7 c2 c5 c4 c3 c4 bb c1 be c2 c3 b4 bc ba ab b2 b2 b3 b5 b5 ae b3 b0 aa aa a7 a7 a1 9d 98 91 8e 94 87 85 85 87 93 84 7e 7e 82 83 81 79 7d 7a 71 6f 78 74 6f 73 6e 6d 6f 6c 6b 6d 6a 66 62 65 61 63 57 60 4c 5c 4f 54 58 69 78 7f 74 6f 5c 3e 2c 13 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 05 0d 0d 17 22 32 44 57 69 71 7f 8e 9c 9f 85 72 64 6b 5f 67 6b 62 6b 68 6a 73 6e 78 72 74 75 7b 86 88 84 85 7e 7c 7d 77 7b 77 7f 83 7e 84 7e 8d 88 93 96 9b 94 90 92 99 95 9d a0 96 9f a5 9f a6 a7 a3 ab ab ab a7 b3 b6 bd ba b9 bd bc ba bc c7 c5 ce c7 c7 d1 d0 d1 d6 d7 d8 e0 db de dc e0 e3 e5 e5 e1 dc dd d4 d4 d7 d3 d3 c1 d2 d1 cd cf c7 cb cf dd ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e9 d1 db d3 e0 e1 e2 da db d6 d7 db d9 d2 d0 dc d3 d4 d4 cb cc ce c5 c7 cb c4 c9 cd c6 c2 c1 bc b9 bb ba bd b8 bb bd b2 b8 ae b0 b3 b0 a6 ad a6 aa ac ac a0 9e 97 a9 9c 9c 9e 8f 8e 8c 89 8d 8b 8b 87 87 78 79 7e 76 83 7b 7a 84 73 75 79 71 70 72 6d 72 77 6c 7b 6a 6e 6b 68 6e 5c 5f 64 5b 53 51 5d 51 5d 5d 63 7c 89 70 6c 63 44 23 10 0e 05 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 1b 23 3d 4f 5c 63 70 81 8f 97 9e 97 76 69 61 61 61 64 6a 65 6b 66 72 6e 71 73 73 70 78 78 84 82 82 86 77 7c 7b 7e 85 82 88 86 81 88 8a 8e 8f 8d 8e 94 91 9a 95 95 8f 8f 96 93 9a 9d 9e 9c a0 a2 ac b3 aa ad b4 ac c0 b6 ba be bb bc b9 c2 bf c2 ce ca d2 d4 d1 d9 d8 d5 db d7 d9 d5 da dd dd d4 d9 d6 d1 cf c9 c3 c6 cf ca cc c6 c8 cc c9 c4 d5 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e2 d2 d6 d5 d6 d3 d1 db d8 d1 ce ce d4 d1 d8 d0 cc c3 ce d3 c5 c8 c7 c2 be b7 bf b8 c3 bd be ba b5 b6 ba b9 a9 ae b7 b1 aa b0 a5 9e a5 b0 a1 ab af a5 a0 9a 9f a5 96 98 90 8e 8d 8c 8e 8d 89 7f 82 87 88 85 7a 87 75 7f 7b 80 7a 76 7a 77 7f 75 74 6a 6c 6f 75 74 6c 6a 64 6c 65 60 65 59 5e 5b 56 59 51 5c 60 6a 7c 7c 71 71 5b 40 2c 12 05 14 0a 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 05 0f 15 16 27 36 50 5e 71 74 7d 8f a4 a2 9a 7b 6c 5c 67 66 67 68 69 73 6a 69 72 6e 71 6f 71 77 7b 7f 7c 85 84 7c 7c 7c 80 7e 84 8d 88 91 84 8e 94
 92 94 97 99 9f 8e 96 8c 92 90 93 94 92 9d 92 9c 9c a0 ae a5 a8 b4 b5 ac b3 b3 b3 b3 ba c3 b9 c2 bf bf c4 cd cc d0 d6 d3 d2 cb d0 ca cd cd d2 d0 d8 ca d1 cb c8 cd c5 cd c9 c6 ca ca bc c0 c7 c9 c7 d6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e2 cf d5 d7 d2 d4 d3 d4 d4 cb c6 d2 d4 d0 cd c8 cb c8 ca cb c7 c3 c1 c4 ba c0 ba b9 b8 bc b6 b5 b6 b4 b0 ad ad ae b0 b0 b3 ab ad a3 9f a7 a0 a6 a0 95 98 95 a1 9c 9c 99 91 92 8e 8c 84 88 8c 7a 8f 81 82 83 82 78 81 7b 83 7b 7e 78 79 70 6b 6b 71 70 72 6f 6b 76 67 68 64 62 63 63 5e 63 62 60 55 4d 5b 5b 5d 67 7b 83 72 6a 54 40 31 1b 10 0e 0c 0c 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 12 0c 28 38 50 58 66 76 80 8e 9e a0 99 7f 62 5d 64 5d 63 62 61 67 6a 69 66 68 66 60 64 71 77 7e 78 78 7b 7d 7e 7c 7b 7f 7a 8a 88 84 92 8e 94 99 9b a3 9b 93 97 90 92 9c 90 94 91 90 8e 8e 9c 96 9f 9e a2 a1 ac b0 a9 ae ab b3 b2 bd b6 b1 ba bd bc c0 bf c8 bd be c9 c2 c1 c5 c4 c4 bd c8 c8 c1 c3 c1 c3 b5 c1 b7 b1 bb ba be bb c5 c5 c6 c4 cc da ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ef f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 d5 d2 d1 cf ce cd c8 cf cb c7 ca c4 ca ca cb c5 c1 c6 c1 c0 c0 c0 c0 bd bd b0 b1 b9 b7 b1 a7 ae aa a4 a1 a7 9f a7 a6 a0 9d a4 98 9b 9e 96 9b 9a 99 95 92 8f 99 8e 91 90 8a 88 86 87 84 7c 83 80 87 84 76 82 73 7f 81 7b 84 77 72 72 73 74 71 6e 75 78 71 6d 68 6e 6a 67 63 64 60 5d 5e 59 5a 52 5e 55 50 58 5b 76 85 77 69 56 41 30 26 18 0a 0c 06 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 08 12 0e 1e 35 4e 64 6b 7d 87 98 a2 a8 9f 84 6e 61 66 60 64 66 65 6c 69 69 6d 64 72 65 69 6d 6e 6f 6d 79 79 7b 81 89 8c 8a 84 8a 8b 8c 91 94 90 99 9b 9b 96 9f 99 90 90 92 92 93 91 8c 91 8d 96 96 9a 9f a0 a3 a5 ad ae a8 a8 ae b3 aa ad b3 bc bc b9 ba bb b8 be ba c5 ba b8 b2 b7 b3 ba bb ba bf b3 b6 bc b5 b1 ad b5 b3 b6 b9 be bd bb bd ba c4 d0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed e9 e4 f3 f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e5 d1 d4 cb d6 d0 ca c8 c6 c7 ce c4 c5 bf c3 c1 c0 bf c0 c0 bc be bd b4 b6 b1 aa af aa ab af a5 a2 a9 a3 a3 a0 a2 a5 a8 97 98 a1 95 8f 96 93 98 94 8b 8e 83 8f 86 8e 8c 88 8c 87 81 82 83 81 80 7b 7a 7c 7d 7d 7f 7e 86 80 80 78 74 70 6c 6e 70 75 70 74 6b 66 6e 6d 6b 60 6c 5d 55 5f 57 60 59 58 59 60 5d 59 68 7a 83 72 65 5d 46 3a 2d 1c 17 0b 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 1b 1c 31 50 65 75 7d 8c 8d 99 b0 a3 7c 6f 65 5b 68 61 62 66 6c 67 6b 6b 65 66 6c 6c 71 73 71 6a 76 73 72 6f 84 88 89 8b 8e 91 8c 89 8f 92
 90 94 92 92 98 90 92 9a 90 97 95 91 94 97 9b 9a 98 95 9f a1 a2 9f 9f a6 a4 a5 ae aa a3 b0 aa b2 b2 a9 b0 b1 af b5 b6 b7 b2 b0 ae b4 b7 b1 ab ad b2 b1 b3 af ad a8 aa a6 ae b0 b2 b6 b6 ba b6 be c4 d0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb d5 de dd e7 e1 f6 eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e1 ce d8 ca d7 d5 c5 cf c6 ca c1 c7 c2 bf c3 bb b5 b9 be b4 b6 b2 b2 aa af af a8 a2 a9 a7 ae a3 a1 9a 9e 9a 9a a0 9a a1 91 8e 8e 88 95 89 8a 8a 8d 8c 86 83 8d 87 8a 87 89 85 8b 7d 83 83 84 7e 82 7b 81 77 7f 84 7f 79 79 7e 84 78 72 72 71 77 73 70 70 77 6c 73 64 63 61 64 6b 5d 5f 57 64 61 5c 5e 5d 5f 59 6f 75 7f 7c 6b 57 4c 3e 2b 26 0d 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0d 03 09 12 2e 43 69 6c 7b 89 95 9d aa a1 79 6b 61 67 66 64 60 66 65 66 6a 67 62 67 68 68 6e 75 72 67 70 71 70 75 7d 83 7a 7f 90 89 8d 8c 85 80 88 81 90 84 8e 8e 95 8f 8a 90 8b 8f 97 93 91 98 92 91 a1 9e a0 9a a1 9a a0 a4 aa a3 a8 a7 ab b7 b0 b0 a5 b5 b3 b2 ad af ad ae a6 ae a7 b0 af b6 b0 ad b0 af a8 a0 a9 a9 a7 ab aa b0 b0 b6 b1 b0 c1 d0 ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 e1 cc c1 c4 d0 d1 d3 d8 c0 e2 e9 ea eb f4 f2 fc fd ff ff ff ff ff ff ff ea d3 da d5 cb cf d2 cc d1 c5 c6 bf c1 c6 bd b8 b7 b2 b9 af b6 af af aa a8 a5 a6 a7 a1 99 99 a2 97 99 9b 92 93 9a 8f 8e 8d 8c 90 87 8b 90 88 87 87 86 82 88 83 81 87 85 89 87 81 81 7d 7f 76 78 7a 79 81 79 7b 74 7e 74 79 81 76 70 74 6e 70 6e 6f 6e 74 6e 67 6b 6b 66 60 65 64 61 5e 5d 5e 5a 58 5a 52 5b 5a 66 7b 7c 75 6a 5c 4b 3f 34 27 1e 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 0a 0f 17 26 3e 58 6f 78 93 9e a6 a8 98 78 64 60 5d 5b 66 5c 62 6a 66 6b 6f 65 69 5f 65 67 69 6d 6d 6a 6b 6b 69 73 72 7a 84 80 8c 89 86 83 81 7b 7e 81 7f 87 93 8c 90 8e 92 90 8c 95 94 94 97 8d 9b 92 9e 91 9c a1 a1 a9 a5 9c a3 a3 a8 a5 a1 a9 ae a7 a7 aa ac b1 a6 b2 b0 aa a8 ac ad ac af b4 b1 ab a2 a7 a8 a7 a8 a7 a6 a8 ae b0 ad b7 b6 b6 d0 ff ff ff ff ff ff ff ff ff ff ff ff d5 d6 c9 be b6 ac b5 b7 b9 bc c1 c9 ca c7 cb d4 d9 e2 e0 e6 f6 fa ff ff ff ff ff ea d8 d6 d3 d4 d0 d1 ca cd d0 cd b7 bd bf ba bb b3 b0 aa b0 a3 a6 aa a7 a4 a1 a3 a3 9f 9d 99 99 9e 94 92 8f 92 93 91 90 8c 87 82 7f 87 80 80 7f 79 82 84 7f 81 82 84 7e 7e 7b 84 7a 7e 85 81 76 72 70 7b 7c 82 7b 7b 78 7d 7b 76 73 69 73 72 72 6b 73 6f 6a 6d 66 6c 5e 64 64 61 60 5d 63 5a 61 4f 5c 56 53 5c 57 6f 75 74 6e 62 49 42 39 2a 19 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 09 15 10 15 23 3b 5b 6d 7a 85 97 a5 a6 9d 82 70 62 5a 66 63 64 6a 62 72 66 6b 69 69 6c 6c 6d 68 6c 71 6f 70 66 68 64 70 73 7d 85 90 8f 89 81 7c
 81 80 7c 84 7b 84 8e 8a 8e 8c 8e 93 92 92 8e 95 9a 93 99 98 98 9a a3 9e a1 9a 9c a0 aa a1 a3 a5 ab a8 ad bb bc b1 b0 ab b6 ad b3 ad ae b4 ac b0 bb ae b4 ad b1 a4 b1 b5 a5 a5 a8 af b4 b8 ad af b3 d5 ff ff ff ff ff ff ff ff ff ff ff d9 c0 b8 a4 9b a0 9c a4 ac a6 b0 b2 b2 b6 b6 bc c7 c5 d2 da df ec f5 ff ff ff ff ff f9 e1 de d8 df db d5 d4 c4 c4 c4 cc bc c4 bb bc b5 ac b1 b1 aa a6 b0 a2 a7 a8 a2 9c 9b 9c 90 94 8e 90 89 92 8e 8d 8b 89 8c 8d 89 88 7c 7e 77 80 7a 72 80 7a 7d 74 7c 7d 81 82 80 78 80 7e 76 76 79 7d 82 75 7b 7f 7b 89 79 7e 78 71 76 75 6d 75 6e 6d 71 74 71 70 61 60 66 69 60 5d 60 5b 55 60 5d 5a 5e 58 5f 64 6d 7e 7a 70 64 53 50 3f 2b 1b 0f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 10 05 0a 11 0c 10 1a 3a 52 64 7d 8b 90 a8 9b 9d 7d 64 5f 64 67 61 6a 64 63 6c 6c 63 69 6b 5f 6a 6b 6f 6b 6f 6d 71 6d 71 69 72 6b 69 7b 86 89 86 7d 7c 81 7f 80 80 7c 83 85 8d 8c 91 96 90 8c 96 8e 94 99 95 97 90 96 90 96 90 9c 9a 9b a4 99 9f a5 ac ad af af b4 b9 b0 b7 b5 b8 b7 b2 b2 b7 b3 b5 ba ba b3 b3 b0 ac b0 ad b2 aa a9 ad b1 a7 a7 a6 ae ba de ff ff ff f9 f8 f5 ff ff ff ff d5 b2 9e 96 96 95 93 97 99 95 9b a4 a8 a0 ae ac b7 bc c7 ca c4 d1 e1 f6 fa ff ff ff ff ff ea e8 e1 e2 db d2 d4 d1 ce cb c8 c4 c3 bd b8 ad ae ac a4 a4 98 a9 9f a0 a0 98 a0 9f 99 99 8f 93 8f 8c 86 86 88 89 8a 81 87 84 81 7a 7d 76 6d 70 72 7a 6b 71 6e 72 72 74 7a 77 76 78 77 78 7a 78 73 76 77 72 7b 79 81 74 71 7d 6b 70 72 71 6d 6e 6b 6f 65 64 67 65 65 5f 64 59 58 5f 5d 58 60 58 5e 52 56 59 58 66 70 76 67 64 53 54 47 30 25 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 0c 13 1d 22 30 44 62 7c 8b 94 97 99 99 71 62 68 61 68 62 5b 67 69 6b 6f 6a 71 61 67 6c 6b 6c 6b 6d 69 67 64 68 69 70 6c 74 80 84 7e 87 82 81 7d 77 7f 7b 7b 7d 79 8a 8f 8c 85 93 8e 90 91 90 94 90 8f 91 8e 8f 8e 99 9c 9e 93 a1 9f a1 ab b0 b1 b7 b7 c0 b7 b2 a6 a9 b1 a5 b0 aa a7 b1 ae b5 a9 ac ac b0 b0 ac a6 b0 a4 a5 a1 aa ab aa af a4 ba d8 ff ff ff e2 d7 dc d9 f4 e7 cc a8 9a 90 8a 84 89 81 86 8e 89 93 9d 9a a2 a7 a8 af bb c0 c2 c6 d2 dd e9 ff ff ff ff ff ff f8 f5 eb ef de da d4 dc d0 cd c4 c5 c5 c2 bc af ae ac ac a8 a3 a2 9b 99 9b 96 96 91 90 90 90 8c 82 90 89 82 85 77 86 7e 81 7b 7e 7e 7c 6e 67 78 71 6e 66 6e 72 70 76 6b 79 76 73 74 71 74 71 72 72 6d 6f 7a 78 76 7e 78 81 75 76 73 75 6c 73 6b 6e 6a 63 67 5e 5e 5d 5b 60 63 61 5d 58 5a 5b 60 59 54 52 53 57 62 79 7d 71 68 52 4f 3f 2c 20 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0f 0d 1a 18 1e 30 41 5f 6e 7e 96 9f 9c 95 72 5f 5d 5a 6d 64 61 67 60 69 69 73 72 6c 6a 66 60 67 65 6a 6d 65 72 68 67 65 72 6d 7a 84 83 86 7a 7e
 79 76 78 7e 7f 82 8b 85 85 90 92 92 92 8f 8f 91 89 81 87 8f 85 8b 94 84 92 90 97 9a a2 9f aa ba c0 c2 bf b3 a8 a4 a0 a6 a6 a0 a8 ac a5 b5 a9 ae af a3 a6 aa a0 a6 a0 a0 98 a4 a4 a0 a3 a0 9e a3 a8 d4 ff ff f8 da c3 bf c1 b8 ae 9d 8c 88 81 7a 7d 84 80 84 8c 95 96 96 94 94 a5 b4 b3 bc c0 c0 c5 cb de e6 fc ff ff ff ff ff ff ff ff f7 f2 e8 e0 df d5 d4 c5 c5 be c1 b8 b3 b8 a3 ac aa a1 a5 99 99 91 95 99 99 96 8d 88 8b 8b 84 84 82 85 87 8b 76 82 84 79 7a 75 7a 71 71 71 70 67 6e 6b 6d 73 6c 73 6c 69 6e 78 78 71 71 6b 74 73 75 78 7b 7f 7a 79 7f 72 6e 6e 69 72 6a 66 62 62 58 6b 61 65 5e 65 5e 5a 5f 60 57 5d 5a 56 58 54 5a 5d 5f 71 75 80 6c 63 55 3d 38 22 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 18 12 23 1d 2f 3e 53 6d 72 8e a3 91 92 77 64 5d 5c 5f 66 63 64 66 60 66 6b 69 63 66 66 63 6d 61 60 6c 67 62 69 66 69 78 78 82 86 86 7e 7d 84 80 82 7f 76 80 85 87 80 97 8a 82 8a 93 8e 90 90 83 86 86 89 86 87 8b 8a 90 8a 8c 95 9b a1 ac b6 b8 b8 b0 b3 a6 a2 9b 9b a4 ab a2 a9 ac a9 a3 aa aa a1 a5 9f a1 a3 97 9e 9e 99 9e 9c a1 a0 a2 a6 b4 d2 ff ff e7 c4 b3 ad 9e 9b 8d 87 79 7e 70 7b 7a 79 83 85 8c 8a 8a 8d 97 9d a9 b5 bd ba c5 c7 cb ce d4 ef ff ff ff ff ff ff ff ff ff ff fc fb ee ed dc c9 c7 c3 b6 bc b5 b5 b1 b2 a4 9f aa a0 a2 9e 95 97 95 8d 8d 84 89 7f 7e 84 81 85 84 7b 7d 78 80 7a 6c 6f 78 75 71 6d 64 6e 6f 60 66 70 6d 6e 6a 6a 6a 6f 70 74 75 6a 72 73 72 79 7d 7b 7c 7e 81 7a 76 78 78 67 6b 70 65 6f 6b 60 6a 6b 5f 60 56 63 59 5f 5e 5d 61 5d 58 53 4c 53 53 5b 69 78 77 6f 65 5b 40 39 20 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0d 11 1a 1a 19 20 2d 37 43 56 79 8e 96 a0 90 72 64 58 55 57 61 5e 69 5d 64 65 5c 6d 6c 68 69 5d 6c 62 64 62 68 69 65 6b 6a 67 75 7c 84 7d 7c 7e 75 7a 7c 72 7a 81 79 78 7d 80 84 80 84 87 89 88 83 7e 89 7e 84 84 87 8a 89 8d 8a 8a 91 92 9a a5 a5 b1 b0 b1 b2 99 9d 9b 99 9e a0 98 a5 a3 a9 a5 a9 a7 a6 a1 a2 94 95 9a 9d a5 9b 9b 97 9e 9b 9d 98 aa cd ff ff ea c7 aa 96 8c 80 7d 6c 6c 67 6b 72 77 77 7f 89 8e 8f 92 93 9e af ae c4 c0 c2 cd ce d9 df eb f5 ff ff ff ff ff ff ff ff ff ff ff ff f7 f3 e2 da cc c5 c7 b9 ae af b1 ab a4 a7 a4 a4 9f a1 9c 9b 92 93 8c 88 8b 82 7e 83 80 7a 7c 77 84 72 7b 79 6f 6c 72 6f 6d 6f 65 68 68 66 6b 70 62 60 68 6d 6c 6d 71 6a 6a 6d 6d 6e 6a 75 79 78 7f 6f 7a 80 7a 73 6f 68 72 61 6c 70 65 64 64 64 57 61 59 54 5f 58 5a 57 55 5f 55 5c 4e 51 52 59 73 75 76 73 5f 5b 48 2e 25 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 0a 11 11 14 20 23 2a 31 32 40 56 64 7d 8c 8f 88 6b 60 5d 64 5f 5d 56 66 62 6c 60 62 68 61 69 63 64 65 63 63 66 66 5f 62 6d 68 70 7a 7c 79 80 75 80 78
 76 78 73 73 7c 80 76 81 7a 79 82 84 86 86 85 83 79 7e 83 75 7f 87 85 82 80 86 8a 90 98 99 9b a1 a5 b0 ae a5 9b 9a 96 97 99 9e 9b a2 a7 a4 9c a6 a8 a0 9f 9e 92 98 9a 93 97 8f 9a 99 9b 98 9b 9d aa c6 ff ff f7 bd a3 89 7d 76 70 6b 64 69 6a 6c 75 78 81 85 92 93 98 9b af c2 c5 cf cc de e1 df e6 ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e5 db cb ce be b9 b2 ac aa aa a3 a3 9f a1 a2 a1 9c 98 95 8f 95 87 8e 81 7a 7e 7d 7c 80 77 80 74 71 7c 77 6f 6b 6b 70 66 74 71 62 64 65 71 64 6a 6a 65 69 6f 70 69 6e 75 77 72 72 71 7c 82 7a 88 7e 83 7c 71 75 69 73 6e 70 67 64 64 6b 5d 62 5e 65 5d 55 60 5d 54 56 57 52 59 53 53 58 54 5f 76 78 6e 5f 60 4d 38 1e 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0a 11 17 1d 1a 1e 32 30 35 41 47 56 6f 89 88 77 60 5d 54 59 69 60 62 5f 59 63 64 5f 65 58 5d 6b 62 67 62 5f 66 62 65 6a 64 66 75 6d 7b 78 6f 72 78 75 72 78 74 76 79 6f 71 77 81 7c 7c 82 83 7e 83 82 78 7f 76 84 7a 79 7e 78 81 7d 87 88 87 98 96 9f a5 a2 a7 a9 9d 9f 99 9a a0 98 93 a1 9a a4 a5 9f 9c 99 97 a3 95 98 98 93 91 92 94 95 99 98 96 a4 a5 bd ff ff ff bf 93 88 76 66 6a 61 61 66 6e 72 71 7b 85 8f 90 9a 9d ae c2 d3 e1 dd e8 e7 f2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e5 d2 c9 c7 b8 b2 ac a7 ab 9e a4 a6 a3 99 a0 97 90 97 8d 90 87 81 83 84 83 85 7d 80 76 7c 76 76 76 6d 6c 72 72 69 6a 6c 6a 6b 6a 6d 69 66 63 6c 6f 6a 68 65 70 6e 77 71 77 73 84 79 84 81 7d 82 82 7c 74 73 70 6e 70 65 6a 68 64 6b 59 5c 5c 59 5b 5d 57 5b 5d 59 56 4f 55 59 56 4e 61 6d 7d 7e 78 65 60 4b 37 20 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1f 25 28 26 37 36 36 47 56 6e 70 6a 65 5d 5f 5e 5d 5a 62 5a 5e 61 55 68 62 5a 5f 5b 67 6a 6a 67 62 68 63 60 60 6b 76 66 72 71 74 67 6e 7a 75 72 77 77 70 72 72 76 6c 79 78 74 78 7b 81 81 7b 7a 73 79 75 75 7b 6f 7b 7c 82 82 86 7f 7e 8e 94 9c 9f 9f a6 9b 95 9e 98 97 9a 95 95 a0 92 9f a4 a2 9f 9e 9c 95 95 91 8e 8c 93 93 95 99 96 94 93 a0 b6 ff ff ff c5 8c 78 67 5d 54 57 60 5d 6d 75 77 7a 82 8c 95 9b ad c2 d1 df ee f2 fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee d2 ca b9 b5 b1 a3 a5 a2 9d 9f 9e a3 99 9b 93 91 8a 92 83 83 85 7f 7a 74 78 74 74 7d 6f 74 73 77 6c 70 73 66 67 6a 64 6b 64 66 69 67 65 65 6b 63 62 6b 6a 73 7a 72 77 7d 7b 83 7a 81 81 87 80 7f 74 73 73 72 71 73 6d 64 65 68 63 64 63 60 5b 5c 57 5b 5e 59 56 52 5a 52 52 57 52 57 62 7d 7d 75 68 61 47 35 18 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 02 06 05 1b 1f 2c 31 2e 39 35 37 48 51 5a 5c 5b 5d 5b 60 63 5b 5e 5b 4d 58 58 5d 62 5d 5d 61 61 61 63 67 67 64 69 61 5f 64 67 6a 64 68 63 75 71 71 7d 6b
 6e 73 70 6a 7a 6b 77 76 74 82 6d 74 82 7f 82 77 76 76 74 74 72 6e 76 6e 77 7a 81 8a 86 8e 8c 8b 9a 9a 9f a2 9c 99 99 91 a0 9d 9d 9e 9f 9d 98 97 9d a1 9c 98 95 8c 88 90 91 8c 9b 8e 93 90 92 97 aa b1 f6 ff ff ce 92 71 67 50 55 54 5a 68 6a 71 76 7b 90 9e a4 b1 c2 da f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 e1 c6 ba b7 ab af a4 a1 a5 98 95 9c 9d 92 96 93 8c 87 84 84 89 82 7f 7b 80 7a 72 79 72 72 7b 75 74 6b 6f 75 6c 66 69 67 68 68 6e 61 6e 65 63 65 61 69 6a 75 74 78 75 77 77 79 83 7d 83 7e 81 8b 7b 79 75 69 74 6c 72 6c 6a 6d 66 66 5f 57 5e 5a 58 56 5b 57 58 55 52 55 50 52 5a 57 6c 81 83 72 63 62 47 29 1a 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 01 06 05 17 24 2d 34 2f 2f 36 46 4b 54 5b 56 59 58 5e 5a 5e 5d 5d 59 5a 5d 5a 52 5c 59 65 65 5d 63 63 62 66 5f 5b 64 67 60 6d 6b 70 67 67 70 6b 69 71 6e 70 74 71 70 6b 72 6b 6f 77 71 78 76 78 7b 7d 7a 7b 79 79 6d 6d 6f 6a 74 74 74 7f 82 85 81 86 89 91 96 9a 9d 95 97 9a 9a 9d 97 a0 9c 95 9d 9a 98 9f 8b 9b 92 9e 94 90 8b 93 8f 8d 8c 92 93 95 9c a2 b2 e6 ff ff d6 86 60 57 50 4e 51 5b 5f 6a 71 7e 85 96 a5 bd c1 e5 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff de ce c2 ae b1 ad 9f a2 9a a0 98 9c 99 96 9c 94 8c 8a 85 84 7e 7c 81 7b 83 7a 74 77 7a 72 75 79 6a 65 72 6b 67 6e 68 68 6d 6b 68 73 6e 69 6a 6a 6b 63 70 74 70 7c 7a 75 81 8b 7c 84 7e 85 78 7b 75 79 78 72 70 70 79 73 68 65 65 63 64 5b 5a 50 54 5a 56 59 5c 63 54 5b 57 54 58 5d 6f 78 87 78 68 60 48 31 1b 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0d 05 17 1f 27 35 39 30 3f 38 4c 60 59 57 5f 53 53 52 56 5b 55 4e 5b 58 59 5d 5a 59 57 64 5b 54 64 61 5e 67 63 60 5f 62 62 65 65 69 6a 6f 6e 63 6b 73 6d 6a 6d 6f 6a 71 6b 75 6d 70 76 73 74 77 81 7c 78 6f 67 6e 6c 75 6f 66 71 70 72 79 77 81 85 8b 8c 86 8f 91 97 94 91 94 9e 8f 96 9a 92 9a 98 9c a0 98 92 96 8f 8e 8e 8b 8a 8a 8e 89 8f 8a 8b 8e 95 a4 d3 ff ff dc 84 65 5b 48 4a 48 59 55 6c 73 7e 88 9f b8 d0 da fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc e4 d0 bd b9 aa a0 9b 96 9b 9b 96 9b 94 90 8e 8d 89 81 82 81 79 71 7d 7d 77 79 7b 6f 76 70 6a 77 6d 72 72 6e 6b 67 69 6c 61 72 66 66 69 64 6a 64 5f 6a 68 74 70 76 7c 80 7d 81 7b 7a 7e 7c 7e 77 73 78 6d 6a 69 6f 6f 71 64 68 61 62 58 5b 59 51 52 55 55 54 53 5b 4f 52 50 4c 5e 61 71 7f 85 7c 64 56 46 2a 17 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 09 1f 34 37 3c 41 3a 42 48 53 54 56 5b 51 4d 55 5b 56 64 5a 59 5e 56 57 63 57 5b 59 58 55 5f 5a 6b 65 5e 62 62 66 62 6a 62 65 61 66 64 70 72 6a
 6a 71 70 6d 74 67 71 68 6b 73 6b 6e 75 70 74 7d 74 6d 72 6a 77 71 6c 6b 71 75 76 80 79 82 88 8c 87 8a 8c 93 96 93 94 9a 99 9a 94 97 98 93 93 91 97 a0 97 90 8c 93 88 87 87 8a 93 8b 88 8f 86 84 8c 9e b9 ff ff d3 86 5d 4f 42 4b 56 54 5e 72 7d 8c 9b af c9 d9 ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea ce c0 ac ad a9 9f a0 9d 97 92 97 99 8f 95 93 84 86 85 75 7d 7a 7d 72 77 6f 73 6f 74 6e 74 74 71 6c 6c 6e 68 6b 62 6d 6e 6d 69 6e 69 6f 68 63 63 6b 6b 67 72 77 76 7c 75 80 79 7d 7d 7a 75 78 74 71 6e 70 70 6a 72 6f 6a 67 63 5b 5c 54 56 51 53 58 53 56 56 52 52 52 52 52 54 64 6d 7c 7e 73 63 53 3f 21 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 01 06 09 12 20 2f 3f 47 4a 41 4c 49 5b 5c 60 51 59 51 58 5d 5f 59 56 51 58 55 58 60 58 5b 60 5e 54 56 61 61 60 5b 61 5a 60 6f 65 62 6e 69 70 69 6f 72 72 67 6a 6f 67 70 6e 68 6b 69 6d 72 6b 72 6f 7a 7a 79 6c 6b 6b 63 6f 71 6f 73 75 74 7d 7c 75 7c 84 80 7c 8b 90 8f 8e 93 95 9b 9d 95 99 97 9f 90 96 9a 99 9c 93 90 91 88 8c 93 85 8e 8a 8d 8a 87 8d 9d 9d a4 f6 ff cb 79 5b 43 45 4d 4d 5d 61 71 87 8f a1 bc dc f2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 d4 c4 bd ad a7 9d 98 9a 9c a0 94 96 96 90 92 7e 85 7d 7d 7e 77 7c 75 72 70 75 77 74 70 75 76 6e 72 71 75 69 68 76 68 6d 65 6b 66 6e 6e 68 6a 6b 6d 77 71 71 78 7e 78 79 7a 75 77 7d 77 75 75 72 75 70 72 74 6f 72 74 6a 67 62 5b 58 59 58 5b 4e 54 56 4e 51 4f 4c 4a 55 53 4d 63 72 74 7c 70 5f 52 37 1b 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 0f 1d 26 42 4f 49 55 41 4b 5e 57 5a 5c 58 5a 55 5b 5d 54 5c 54 61 5a 5f 5f 5c 5d 60 59 54 5d 5b 5e 61 5f 5b 5b 5f 63 69 63 67 69 6b 63 69 6e 68 64 74 6a 65 6c 71 66 6b 71 70 65 63 6a 6f 71 72 72 66 62 6a 69 6d 6d 76 74 70 74 78 79 7c 7d 79 7c 86 83 8b 8d 8c 8e 94 93 8f 8d 94 99 8f 99 95 9c 95 91 84 8a 8f 87 88 8c 84 88 87 7d 87 8f 94 8a 95 a3 c0 fa bb 72 55 43 47 49 49 5e 62 77 87 98 b3 ca ea fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e0 ca ba ba ae a0 9c 95 99 98 95 97 97 8e 88 8d 83 82 7d 73 7b 6e 73 71 6d 73 6e 6d 66 6d 76 6e 6f 73 63 67 68 6b 6f 60 63 65 68 60 71 5f 67 62 64 71 70 71 72 7a 7b 75 78 6a 74 6f 76 70 70 71 6f 72 6f 6b 67 6a 6c 65 64 59 5c 58 59 55 59 4a 4b 50 4e 53 4c 52 4d 4e 50 52 69 76 85 7e 6f 5b 49 2b 1a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 1a 2f 3d 4e 60 59 55 61 67 64 61 4f 54 55 5b 57 5b 5c 5a 5a 5a 5a 5e 5f 5d 5a 54 5a 60 61 5b 5e 5a 5c 5b 64 60 64 64 64 67 6a 65 68 68 60 6b
 66 64 6a 66 65 69 66 67 68 68 67 60 69 70 74 75 6f 60 62 6f 66 71 72 66 77 67 76 6d 76 77 74 74 7f 7e 80 85 7d 86 94 8e 8e 9b 96 a0 95 99 91 89 97 92 91 92 93 91 8e 87 83 85 83 84 8b 82 8d 8f 92 96 9b a7 c8 ac 76 51 41 41 45 4d 5d 6a 7e 95 af b2 d9 ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 d4 cd bf b0 a3 a4 a7 9b 9d 8a 98 8d 90 8b 87 8f 79 7b 7a 7a 79 75 76 6f 6e 69 75 6c 6e 70 6d 6e 64 6a 6a 6a 70 62 6c 67 6c 66 6c 69 60 6a 66 63 68 70 6d 75 70 6f 77 6f 76 72 72 70 6e 72 66 74 5f 65 6f 68 5f 6a 62 54 60 63 52 55 56 53 51 49 59 53 4f 4d 50 4b 4d 52 52 52 64 78 86 7e 74 5a 45 21 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 08 16 29 42 4e 62 65 5f 6e 6f 7b 6c 5d 51 50 5b 54 5f 52 57 5b 54 5f 5b 57 5a 5a 5c 53 59 61 5a 5a 5b 5b 5f 5d 61 64 62 63 62 66 64 60 65 68 65 67 6a 69 64 6d 6d 73 65 69 67 69 6a 67 6e 68 6a 68 71 6f 6b 68 6c 6a 78 6d 71 78 6f 70 78 73 7a 74 7e 84 85 87 8c 8e 8e 93 93 9d 97 9b 9b 8e 8f 95 8c 8d 8a 8d 91 85 85 87 8a 85 85 86 81 85 89 88 8f 93 91 a3 9e 79 50 47 45 44 52 5c 72 84 9b ae c5 d7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 d9 c4 ba b3 a5 a1 9d 99 99 93 9a 91 8d 8d 82 85 83 80 75 72 72 6c 72 6e 70 6e 72 73 6f 70 6c 69 6d 6e 63 6d 63 73 67 66 6d 67 69 62 67 6b 6a 6a 63 6f 6e 76 7c 78 77 68 74 6e 6d 66 6b 65 67 65 64 67 69 67 66 63 64 61 62 66 5a 5a 50 58 52 50 4f 4a 51 5a 52 58 55 4c 53 53 65 7a 7d 76 67 56 3e 18 07 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0b 25 42 55 60 76 75 76 7a 7f 75 62 5f 55 57 50 5e 5a 61 52 5d 57 5c 60 5e 5a 57 56 57 5d 5c 5d 5a 5d 61 61 5d 64 61 62 6a 62 66 65 5c 63 61 60 5f 67 64 62 6b 61 65 69 6e 69 64 65 6a 71 6a 69 62 68 67 63 6a 6d 72 68 61 6c 6a 6a 64 71 76 7c 7d 79 84 85 91 81 95 94 8f 90 94 93 95 94 94 97 90 92 86 86 84 85 86 82 7e 86 81 82 8a 83 81 84 8d 8f 89 90 96 6d 50 40 4b 4f 47 61 6c 85 a1 b1 cb e2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e7 cf c0 b8 af a6 a2 a3 9f 9c 8e 98 8a 93 8d 79 83 79 79 7b 77 70 6e 72 6d 6d 6e 63 71 6b 72 69 6b 6a 69 69 70 64 65 5b 5f 67 66 66 61 65 66 63 62 62 65 6e 6d 6c 73 6f 70 67 70 68 69 66 66 6d 62 69 6a 62 62 61 62 5e 61 5d 5c 55 56 51 52 54 55 52 52 54 57 53 57 4b 50 51 56 64 74 7c 78 60 48 2a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 13 1a 3b 55 65 7b 75 7c 80 85 83 69 64 52 55 58 57 61 5b 5e 63 50 54 59 59 54 5e 5e 5b 52 59 56 50 64 58 5e 5a 60 64 63 67 62 64 68 60 5c 60
 5d 6b 66 64 5a 65 60 5d 64 60 5f 66 69 60 70 6b 61 68 67 72 67 6b 6e 68 6a 71 66 63 6c 6c 6b 73 77 73 83 84 83 8a 89 85 91 8e 94 9b 8d 96 8e 91 89 84 8d 8e 83 87 8a 7f 84 85 87 84 7e 81 7f 7e 84 84 85 84 7d 8a 76 54 43 43 45 4d 5f 6c 89 a1 b3 ce f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb e2 d8 bf b9 aa ac 9b a2 92 9e 90 90 87 8c 89 7e 85 7a 75 7a 68 71 72 6c 73 65 72 6c 6c 6c 73 69 69 67 6b 6a 68 68 5e 64 61 63 64 6f 61 59 5e 63 64 68 64 66 70 6f 72 6d 66 69 67 62 6a 6b 61 62 5d 61 62 63 5f 64 5c 59 5d 59 55 58 54 54 49 52 4b 55 4f 52 55 52 4e 4f 4e 57 55 6b 7b 7a 70 56 3b 26 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 09 0c 19 30 4b 67 79 7e 83 81 86 91 7c 71 5a 59 5e 68 64 66 68 5d 5a 5c 59 59 62 56 62 56 54 53 54 5b 5d 5a 60 60 57 6b 63 5e 68 63 5f 5f 65 67 5e 6a 63 60 63 64 68 64 5c 5e 5f 61 63 74 69 69 5e 63 66 64 66 64 69 64 6d 6b 64 6e 68 67 70 74 75 7f 76 7b 7c 85 87 8f 95 91 96 a0 8c 90 90 84 8d 8d 8c 84 83 7e 81 84 89 7d 86 7a 89 7b 82 7f 81 88 85 84 82 82 70 4d 3c 41 46 5a 61 76 8a a4 b1 cd f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 d9 c9 b5 b3 ae a6 9f a6 96 a2 95 90 90 8b 85 80 74 78 71 71 65 6d 71 6b 69 70 66 73 77 6b 6a 6f 69 69 6e 64 64 6c 65 64 69 65 61 60 60 66 60 68 61 62 67 71 72 6f 72 69 66 65 69 64 64 6e 5b 69 61 5f 66 5f 65 5f 59 63 5c 60 5a 5f 5d 56 52 53 53 51 52 59 55 53 54 58 4e 54 63 6a 79 76 69 43 22 1d 06 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 05 07 0b 17 28 41 5f 67 77 8e 8a 8d 90 82 79 60 61 60 6a 74 7e 76 6c 62 5d 61 6b 72 62 5f 5a 52 60 5d 5a 59 56 5b 5e 5f 67 6a 5a 5c 5c 63 5f 65 5f 5f 61 62 65 5e 5d 60 65 60 64 5e 5e 69 66 6a 65 60 67 64 64 64 62 6d 5d 67 67 63 6a 68 62 70 73 72 79 7f 7e 7b 83 88 89 8d 8c 97 9d a1 9a 95 92 87 84 85 8f 89 8a 87 8c 84 7a 89 7a 79 80 85 82 7e 7c 7e 75 75 7d 6e 4f 40 49 4b 54 61 71 8f a8 b3 cf e6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb dc cb c0 b7 a6 a4 9d 9c 9d 91 90 8e 8b 8a 81 75 76 6d 69 67 74 6b 6f 6c 6a 65 6a 61 6d 68 66 72 5b 69 66 63 68 62 62 62 5e 5b 61 62 60 62 68 61 61 66 70 6b 69 6a 6d 63 60 6c 62 60 61 67 63 5d 5c 60 66 58 61 5f 5a 61 5a 5b 59 5a 5e 53 58 53 4a 5a 53 61 54 55 52 58 50 56 65 72 7a 6d 58 36 19 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 05 15 17 23 3c 59 67 7e 7c 81 8a 88 79 73 66 60 59 5d 70 70 6c 6e 5b 59 57 6c 76 73 71 60 5b 5d 56 5c 53 55 59 52 61 62 66 65 5e 5d 63 60 61 5f
 64 5f 5b 5c 5a 5e 5f 63 5a 60 58 67 64 64 64 65 5d 5c 62 62 62 60 67 69 6f 67 5d 64 66 6a 6b 6f 6f 6c 6a 82 82 7e 80 87 99 86 a0 95 8f 94 87 8d 81 7e 85 84 7d 85 82 7e 86 7c 80 7c 77 76 6e 76 7a 7c 72 72 6d 74 64 4e 47 44 45 4e 58 69 86 9f b3 c7 e2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 cd c9 b7 b1 ac ac 9a 9e 9d 98 89 85 89 84 7c 76 71 72 75 6e 66 62 68 65 62 67 65 68 64 60 65 66 61 62 66 64 5f 62 62 5e 58 5f 5f 5b 61 5c 5e 69 5b 5c 67 6b 6f 64 5a 64 5c 62 5c 63 5d 64 59 67 52 5f 5b 5b 5d 63 59 61 57 5a 5a 59 54 4f 57 5b 4c 51 52 57 58 57 52 56 57 5c 5f 6e 75 61 48 29 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0d 0b 11 1f 29 52 6a 7b 7c 86 88 85 76 71 5d 5e 61 68 61 66 62 66 58 61 5e 65 73 7e 72 6c 64 64 62 5a 56 53 5b 5f 65 6c 65 60 5a 5c 5d 61 62 63 5d 64 53 5f 61 57 64 5d 62 5a 5a 64 62 64 6b 64 59 60 5e 5e 5e 5f 60 65 63 64 6e 66 67 65 60 68 6e 71 7a 7c 7c 7c 82 81 8e 91 90 91 8b 91 8d 88 88 87 7e 8a 88 7c 84 84 7b 7b 79 78 6d 75 73 7b 73 70 71 6c 6b 72 69 52 3f 49 44 55 61 66 7e 9b ae bd dc f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e3 ce bd b3 ac a7 9c 99 9a 9a 9a 90 91 80 82 76 7c 71 6b 65 69 69 65 65 5a 60 6b 63 63 68 63 68 66 5a 5d 5e 64 64 60 59 5d 60 5f 5d 61 5f 5f 60 63 6a 64 6e 67 67 62 67 69 62 5e 65 62 5b 5b 68 5f 54 5b 5a 60 62 5b 5e 5f 53 54 58 51 52 51 58 54 5c 5b 59 53 58 56 5c 5a 51 54 5c 6b 70 52 34 20 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 0f 0a 08 21 2c 43 63 75 72 7f 89 82 6e 66 57 60 5e 64 67 62 61 5d 59 56 60 58 5f 65 68 69 5d 5f 5f 5f 63 64 5f 69 6e 74 74 6b 60 5d 5e 57 5d 5b 62 60 65 59 57 5c 5b 56 56 5f 5c 5f 66 6a 62 5c 61 61 63 62 61 60 66 63 61 65 67 61 5d 61 6b 69 73 6d 76 74 78 7d 83 86 8c 8b 8d 8c 89 8a 82 83 88 82 83 7f 7d 83 84 84 7b 7b 7b 73 6e 77 72 6f 6c 6e 6b 63 62 67 62 4e 3c 45 44 50 57 6b 7d 92 9c b9 d0 ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed d9 bd b2 b2 ac 9e a4 9c 9d 97 96 90 8c 7e 7f 73 76 73 6c 61 68 6a 66 66 64 5f 5b 63 61 65 60 67 5b 6a 61 5e 62 5d 5f 5d 55 5e 61 61 61 5e 5e 60 64 62 6a 6c 5e 5c 63 64 70 60 64 5b 5a 56 61 63 65 60 55 58 54 5a 59 57 62 5b 5e 5c 57 5d 50 55 5d 58 56 56 58 56 50 53 56 56 54 5d 65 5b 3c 2d 15 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 16 11 1d 19 39 4d 6f 72 81 8b 82 76 60 5f 52 63 66 5c 55 4f 54 59 5c 5f 5b 62 54 60 57 5a 55 59 62 5f 66 66 66 6e 74 73 73 78 6f 64 5f 65 5d
 5d 5c 58 56 5a 53 59 5e 5a 5a 5d 5b 5b 64 5d 64 65 5f 58 64 5e 60 66 65 6a 62 62 5a 5e 65 65 63 66 66 68 72 75 7b 74 81 85 83 83 85 81 86 7d 84 85 82 81 82 7a 82 7d 7d 75 70 7b 72 78 6a 6f 6e 65 67 6f 65 5b 67 65 5d 41 3e 41 4b 5e 67 6d 89 94 a5 bc df ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 d1 c3 a9 a7 a1 a4 a6 a1 9f 9d 90 8f 8e 7b 85 77 76 70 6b 6b 6d 65 64 65 66 5b 60 5b 5e 62 5d 65 61 62 5d 62 61 5d 5d 58 5b 61 5e 59 62 62 60 6b 64 62 61 5f 5b 61 61 59 5c 5b 58 51 5a 60 5a 5a 58 54 59 61 52 58 57 5f 51 60 60 55 59 55 54 5b 56 53 4f 57 59 58 52 48 55 4f 5a 5b 62 52 32 26 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 09 06 05 0e 0f 0e 0f 22 31 49 62 72 7a 84 80 73 68 5c 5d 59 5a 5b 52 57 54 57 5a 57 5f 55 57 56 5b 65 58 5d 5e 5c 63 61 61 6f 6b 71 7c 80 7b 71 65 5b 5f 61 5f 64 5c 5f 59 5d 64 56 5f 5a 5d 64 63 57 5f 63 5e 6a 64 5c 5e 60 60 65 6b 5c 66 60 62 67 68 6d 74 73 72 68 6f 75 7c 7e 82 83 85 80 80 83 85 88 82 83 84 7e 7f 79 70 7a 72 68 73 6c 66 67 63 64 5c 65 6a 5e 5e 65 4d 40 3e 4b 4c 52 5d 71 80 8c a1 bc d1 ed ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e0 d0 b4 ae a9 9f a4 96 98 97 95 96 8b 8b 7f 7b 75 71 66 66 5c 5f 5d 5d 69 66 66 69 63 68 62 66 6c 5c 5b 5c 5a 57 62 5b 5d 5c 61 60 5f 60 62 60 66 5b 5a 5f 5f 5a 63 5e 5e 5f 55 5b 5a 5c 63 5e 58 59 58 53 5b 57 5d 5d 5a 53 58 56 59 61 57 5b 5d 60 56 59 56 54 55 54 52 54 4c 5a 5d 54 49 38 20 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 13 12 19 23 24 3d 49 65 6f 83 81 7c 6d 56 50 58 52 51 53 56 5d 5e 5d 62 5c 5a 4e 5d 53 5f 51 57 5f 63 57 5b 60 5b 64 69 70 79 7a 6e 64 59 5f 59 5f 60 59 5c 56 5c 56 63 5d 54 5e 61 61 59 64 61 64 62 68 63 69 63 62 59 5e 65 64 66 61 66 6c 65 66 72 6d 73 79 72 77 85 7e 85 81 82 80 84 87 7e 80 78 7f 83 83 80 7b 7c 79 7f 6f 6a 6b 62 61 62 5b 59 5b 57 50 59 4c 3c 41 47 54 55 5e 69 77 81 9b ad c6 da f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 db ba ae a3 a3 a0 94 9c 9a 99 90 95 8a 89 7e 7b 72 72 66 65 6b 62 5f 63 62 5a 63 61 62 64 65 64 61 6e 68 5c 63 63 5d 5f 67 56 5e 64 66 69 67 69 61 59 58 5c 61 5b 59 5e 5b 52 57 59 5a 55 54 5f 5b 62 59 60 59 5d 5d 5a 56 58 56 59 5c 5d 5b 5a 54 5c 61 5a 5c 55 59 4f 5a 52 57 54 56 50 32 26 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 0b 06 05 0a 06 11 0d 19 1d 34 42 54 6c 71 88 7a 6a 60 57 56 56 58 50 52 5a 5b 5b 5a 52 5b 4c 48 50 52 59 5b 4f 5b 59 58 58 5b 61 63 65 6b 77 61 5b 58 5b
 56 5f 59 5b 5d 60 5b 60 5e 5f 57 66 62 56 63 62 61 64 65 67 69 5d 66 62 66 5b 5e 5f 5c 62 6b 66 68 68 66 6f 69 6f 71 73 83 73 7c 81 85 84 81 84 83 7b 7e 7c 7c 82 80 79 7b 6b 6d 6a 62 62 64 5d 5d 5a 5c 56 57 4f 59 4a 3d 43 40 48 58 54 58 6f 7a 84 95 b3 c7 dc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee c4 b9 ac 9d 99 91 9b 98 94 97 95 89 85 82 72 7d 6d 6e 68 62 62 63 5f 65 5c 5f 60 64 5f 65 5e 68 68 64 62 5f 65 67 60 61 5c 5f 52 60 5f 5d 5f 5c 5b 66 57 57 60 53 5b 59 5a 54 5c 55 61 57 55 5f 59 57 59 52 53 57 5f 57 5a 51 5a 5b 57 5c 5a 51 5e 59 60 59 56 50 52 51 55 51 51 56 4f 3e 35 12 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 10 12 18 14 24 25 39 41 5b 6e 77 82 6f 66 5d 56 51 4e 51 5c 53 5e 57 58 50 55 56 55 57 53 5a 60 5a 54 58 65 5c 5a 65 5b 65 66 68 65 61 64 5f 5e 58 5b 5d 53 5d 56 5a 62 60 63 68 65 69 56 63 68 5f 69 65 63 6a 5e 66 62 69 64 65 61 65 66 64 62 68 65 6d 66 69 73 77 74 7f 87 80 7b 7d 79 7f 81 7a 7e 81 7e 79 78 75 78 78 76 6b 62 61 57 62 5f 5f 5a 48 50 4e 4f 4d 36 3e 49 48 51 4e 59 69 71 83 91 a2 ad c6 e8 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e2 c4 b2 9d 99 99 96 9a 93 8d 8e 87 8e 7d 7e 7d 79 6b 6f 61 65 5e 5b 57 62 5b 62 63 69 66 6a 6a 61 66 61 5b 5c 60 5e 64 62 5f 5b 61 61 60 64 5c 57 5e 58 57 5a 58 56 5c 5a 54 4e 58 50 53 5f 54 5a 5a 54 61 57 53 52 57 58 53 54 51 54 5e 5a 5e 50 57 5f 59 57 58 54 4f 4e 4d 51 5f 57 4d 39 1e 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 02 06 05 07 15 0e 16 1c 24 27 30 3b 47 5f 76 7f 78 70 60 52 5f 54 55 57 5b 54 5d 57 5a 53 5a 59 59 56 54 54 60 61 55 5c 51 59 62 62 64 67 68 5d 5f 5f 63 61 68 64 5e 5c 5a 61 60 5e 6f 6f 6b 68 6a 66 62 66 6f 6a 70 65 6a 6f 6b 72 61 65 65 6c 62 66 69 62 6d 64 72 70 6f 6e 79 74 81 7f 83 82 7b 80 83 76 84 83 79 77 79 7a 77 71 70 74 6e 63 64 5f 5c 59 55 55 54 51 51 4e 44 37 3d 45 48 4f 50 5b 6d 73 81 82 9e a7 b5 d6 e8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 dd c3 ad 9e 9c a0 97 96 9b 90 8c 8e 86 7c 7e 77 6b 76 6d 62 63 65 64 5b 5f 61 61 60 64 65 6b 69 6b 6a 6f 66 5e 6a 63 65 62 5d 58 53 5e 5c 5e 60 5a 56 5c 52 58 5a 5a 5b 59 5a 58 5c 5d 67 64 57 59 4f 60 5d 5a 5c 60 50 5b 5c 59 61 53 5c 57 54 56 54 5a 5a 53 5e 54 55 5d 55 5b 5c 57 40 32 16 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0c 0e 15 11 16 1c 15 30 31 3c 55 63 71 82 75 5c 55 4f 56 53 53 5b 53 51 58 55 4c 5b 54 58 55 58 5a 58 56 59 58 57 5a 55 5a 5f 65 6d 5e 5f 5f 69
 70 70 63 61 64 59 5f 62 61 69 64 73 73 6d 70 71 67 73 6a 71 64 6e 6e 6d 6c 64 6a 6c 5d 60 65 68 62 63 5f 5f 6c 70 63 76 74 7e 80 7c 80 7e 77 6d 80 76 7b 83 79 78 7a 78 74 72 60 5d 5b 59 58 5a 5c 52 4f 44 49 4e 47 45 36 34 3b 43 51 49 52 5e 64 75 7b 8e 9d ac bd d6 e6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee cd b4 a6 9b 90 92 86 91 90 90 8d 88 80 77 7c 6b 70 69 67 66 5f 5c 59 5b 58 5e 60 68 6b 66 64 67 60 68 64 61 60 63 63 5d 5b 55 54 58 50 5b 5a 58 53 54 57 53 4e 4a 51 5c 59 5e 54 57 52 55 5c 5a 59 5a 59 54 54 5e 4e 54 56 5a 5b 5d 52 57 5a 5e 53 58 55 56 51 52 52 54 50 5a 52 52 48 26 25 0b 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 12 15 1e 1d 1d 1e 27 22 36 43 56 6b 76 77 68 60 58 54 56 50 5b 57 55 54 4b 57 51 55 59 55 5e 5a 5b 5a 64 56 5b 5c 5a 57 66 61 67 67 6b 7a 79 75 78 66 6d 67 64 61 63 67 6c 67 66 6a 69 71 74 72 6c 6e 6a 69 60 65 63 6a 64 68 66 68 66 65 62 68 6c 67 72 6d 6a 6b 78 77 7c 80 70 77 79 74 7d 78 72 74 7e 7a 7d 74 74 6d 72 6b 61 5c 5c 5f 53 51 51 55 45 45 3e 48 40 2a 2f 3b 3d 45 4f 57 57 62 72 73 88 8f 9b ae c0 d7 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dd be aa 9c 9c 90 8e 8f 8f 8d 8d 87 89 7b 7a 75 6a 68 71 63 5f 61 5d 5f 5c 5b 68 62 62 64 67 67 63 5f 6a 5d 5d 60 64 5c 5e 57 5a 5c 57 5b 57 56 54 50 57 4c 50 55 5a 4c 4d 4f 57 51 52 5c 57 54 57 56 56 5e 55 5a 55 54 5a 4c 56 54 58 58 54 55 4e 58 51 54 4c 51 53 57 54 51 58 4d 3e 39 28 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 06 0d 0e 12 0f 18 1d 20 1e 25 2d 42 54 69 79 84 71 63 58 4c 56 51 57 4e 58 51 5a 4c 55 50 52 5b 54 55 5c 5a 56 57 5a 5d 60 6a 68 67 6b 5e 68 75 70 81 85 80 74 65 60 5e 65 5d 6d 65 67 6f 69 72 65 67 6b 6f 6a 64 64 62 69 65 65 71 68 70 70 64 6e 6d 67 6c 6f 6a 71 76 75 78 71 76 7b 7d 71 77 7b 7b 7b 7a 70 78 7f 7e 71 76 74 6a 68 65 61 58 5b 4a 50 4f 43 41 4e 41 3b 2f 25 2f 39 4d 4c 51 4f 65 61 7f 7c 83 8d a3 ac c1 d5 e5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee d4 be a0 94 93 96 92 8f 92 8e 85 89 7b 7b 72 78 72 6a 5f 64 5f 59 65 57 59 5a 5a 5a 61 67 67 5e 5f 5d 63 5c 5d 64 58 64 5f 5f 59 54 4e 55 56 57 5b 50 4f 4f 4d 4f 56 50 53 5e 5b 5e 52 58 57 56 5c 63 5e 5f 51 57 50 59 55 59 57 56 57 50 5c 56 57 4e 5d 59 49 54 55 56 5d 51 4c 47 3c 32 20 08 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 09 0e 19 19 1c 15 1a 24 34 37 47 5c 6f 85 7a 69 5e 53 52 52 57 4d 57 51 59 55 4d 50 5b 52 5c 5a 5f 60 5c 5a 5d 5f 60 62 5b 5f 61 62 64 66 6c
 70 7c 74 6c 6b 66 65 64 69 5b 63 5d 65 69 62 62 6d 64 64 61 65 64 61 69 6a 64 60 62 6e 69 6b 76 77 75 6c 70 60 6e 75 72 7d 74 7e 7a 7e 71 72 73 7b 7b 77 7f 76 75 77 69 73 6f 63 5c 5b 65 59 54 53 56 4a 4a 3e 41 41 3b 26 27 2d 39 3e 46 4c 54 5c 63 71 79 7f 89 95 a5 b2 b6 d5 e6 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd d1 cb af aa 99 8f 8e 84 87 82 7b 7f 78 75 72 6f 6f 62 65 5d 64 5f 5c 5a 52 55 5b 5a 63 60 62 61 62 62 5f 5b 5c 56 53 5a 5c 56 57 50 51 56 54 58 52 52 4f 4e 58 50 57 57 5d 54 5b 58 50 50 55 59 53 56 5f 56 56 4f 55 50 53 53 55 53 52 4f 5a 53 58 52 54 56 56 4a 50 5a 58 54 4b 4b 34 2b 27 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 09 15 11 1a 1c 20 20 2a 2b 34 47 51 65 79 7f 6a 62 53 55 49 4c 54 57 53 5b 58 53 59 5a 59 56 56 5b 5b 5f 59 62 5c 58 5e 58 5e 64 66 6a 6a 5c 66 6f 67 5c 61 5d 5c 55 5b 5e 62 55 5b 5d 59 64 63 61 61 5f 63 5f 6b 5b 66 62 65 64 68 69 6b 7a 79 76 7b 72 7b 7a 7b 76 7e 74 7c 7c 6d 71 72 78 76 78 6d 69 73 6e 71 6e 6c 6c 65 62 53 5d 5b 59 51 4a 44 3f 3e 3d 3a 37 22 1f 26 28 32 42 47 59 5a 69 6e 76 7d 7e 86 87 98 a3 b1 c6 d5 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb de cb b0 a7 94 90 8a 8b 85 7f 85 89 80 81 79 7c 6e 6c 63 5e 60 5a 54 59 5e 5d 5b 5e 5b 5b 57 65 5d 65 5c 59 5e 61 57 52 57 57 50 4b 4a 4d 52 55 50 56 4e 51 4b 54 54 5c 52 50 59 59 56 5c 59 5f 64 61 63 59 5a 53 55 57 57 52 55 56 51 56 56 50 55 4e 4c 4b 51 53 53 50 5a 4b 4a 44 3f 3b 25 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 07 0e 0c 12 18 1d 1c 17 22 24 38 3f 53 5b 6e 83 7c 69 56 53 55 4d 48 50 56 55 52 51 4e 54 59 58 58 5e 5c 5d 54 51 5e 5b 5d 5c 56 5b 63 6b 66 67 6d 6a 65 63 5e 60 58 64 5b 5e 59 5d 60 60 5c 5c 66 60 66 60 60 67 62 69 65 65 65 5e 5e 6e 65 6d 70 69 6f 7e 7f 82 85 72 7b 7e 7e 7c 75 7a 6d 75 73 6c 74 7b 70 70 76 69 6b 61 6c 64 57 59 51 4e 4b 50 4b 4c 44 3b 3e 3a 23 17 27 1b 32 33 41 4e 5b 5f 67 74 71 7c 86 87 91 99 9f b5 c3 d4 e8 ff ff ff ff ff ff ff ff ff ff ff ff ff f9 e3 d0 bf a3 a1 92 8b 88 7e 7e 81 7e 81 76 6e 78 6e 69 6d 60 5f 56 64 52 60 60 5a 60 5f 5f 61 58 5f 5e 63 5b 5f 5a 54 52 58 59 54 4d 54 51 57 57 52 4f 51 51 50 53 5c 54 60 5a 5d 5e 61 5b 60 61 5f 62 5b 62 5f 53 5a 54 56 54 54 58 50 54 55 4a 59 4a 53 54 4c 53 52 44 53 57 50 49 41 39 25 1c 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 05 01 0c 14 1c 1e 1d 25 2a 23 35 3a 47 61 70 75 78 6f 5f 5d 54 4f 56 4f 56 5f 52 52 57 54 54 5a 5b 5b 59 53 5b 56 5d 64 62 5b 60 5e 5e 5f 62 64
 66 67 67 61 5e 5b 5e 60 5a 5e 5d 64 65 61 61 59 67 62 5e 65 5e 60 59 61 60 62 61 6a 60 63 63 65 6b 6a 68 75 79 79 79 7c 86 7b 7c 82 7b 6d 78 76 74 76 74 7a 6f 72 7a 6f 66 6b 68 65 5d 5d 54 54 52 57 50 3e 45 3b 42 3d 25 16 1b 21 28 2d 3d 4c 4e 58 63 64 6a 78 77 7b 8a 8c 8d a2 ac c1 d4 e7 f3 ff ff ff ff ff ff ff ff ff fe f3 da d0 bf b1 a2 96 87 84 80 76 80 7c 7d 7e 7c 79 70 6b 6a 6a 57 5e 66 58 5c 53 52 5e 53 58 62 59 65 66 65 64 63 5f 5e 5d 56 4b 5b 55 4f 53 4c 58 57 54 4c 5e 5c 5a 64 5c 5a 59 56 57 5c 62 5b 5f 5f 65 62 64 61 60 58 53 5e 53 4d 4e 56 5a 55 57 4a 4f 51 51 59 55 4f 53 4d 58 4c 45 49 40 3a 25 14 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 0c 0e 13 11 27 24 2a 2b 2e 37 39 4f 66 76 82 7d 69 57 4d 51 49 52 4d 52 4b 57 4e 56 5f 5b 5a 5b 55 52 57 53 5e 5e 59 4b 51 5b 5e 5b 5a 64 61 64 5d 58 5a 60 57 57 5c 5e 60 56 64 5f 6f 63 5e 5d 6b 60 64 61 60 67 68 6a 5d 67 5a 61 65 64 62 66 6a 6e 73 78 7b 75 7b 78 7e 76 72 78 7a 70 6f 79 7b 70 73 74 77 72 69 65 64 64 57 5b 54 53 51 49 4b 45 45 39 3b 35 25 11 1e 1e 24 27 30 38 45 52 55 5f 6c 77 73 71 77 87 8d 94 9c ac bc c4 d5 dd e9 ed ed f2 f0 ff f6 fd e4 d9 ca be b5 a6 9b 91 85 82 83 76 81 7c 72 79 7a 74 6f 6b 67 66 66 5a 5c 53 58 55 5b 5c 5c 5f 65 59 5f 61 5f 60 59 5b 56 55 58 57 51 54 4c 4d 54 57 58 50 51 5d 5c 61 61 55 56 5a 55 5b 5d 5d 52 54 55 5f 5f 62 5a 5d 5c 58 56 4f 4a 50 54 4e 4e 4f 4a 52 55 4b 4e 4e 48 51 45 4a 49 46 49 38 33 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0e 14 10 1f 23 29 2b 29 30 33 40 51 5e 67 88 7f 6d 5d 50 4e 4d 54 51 4e 53 50 52 50 55 55 55 55 59 5c 52 54 57 5b 5d 57 5d 5f 51 5c 58 5e 66 5b 59 58 58 5e 5d 5b 62 64 5d 64 55 6b 63 61 65 5f 5d 66 5f 5a 67 5f 62 60 69 63 60 63 62 64 64 67 6a 6b 68 67 6f 74 78 76 73 73 73 75 78 6d 76 6c 75 71 75 6c 6e 66 5f 6d 66 5f 5c 5e 59 53 4f 50 4b 3e 3a 3a 38 34 23 14 16 18 1a 20 29 41 44 49 54 56 64 6f 6b 72 79 7e 7e 87 92 9d a8 ab c0 c1 d2 d4 d1 df e4 ea ed e1 de c9 bd b5 a2 9a 98 8c 87 82 83 7a 7c 75 7d 71 6d 70 73 6c 68 64 60 62 5b 61 63 58 5c 56 59 5c 5a 5b 63 5e 5e 60 63 5f 60 56 5d 61 57 54 52 51 52 5e 5c 51 60 5e 5e 58 57 5b 52 56 58 5d 5b 58 5c 52 53 57 56 58 5d 6d 57 56 52 5a 55 4f 53 52 54 4d 4d 4c 52 49 57 49 46 52 4c 4f 4d 4c 45 34 22 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 12 0d 0e 1b 1f 26 23 2c 2b 39 44 46 58 67 75 81 70 64 52 52 4d 4f 57 54 55 54 46 4f 53 64 53 5f 5c 5a 54 50 5b 59 55 55 59 58 5c 58 4e 5a
 5b 4f 55 55 56 5b 52 55 5e 5d 63 69 61 5e 65 5c 62 60 5d 68 61 5f 66 58 66 60 5d 62 5e 68 6e 66 69 68 6f 6e 69 6f 70 72 71 6e 6d 70 72 6a 75 71 73 75 76 70 75 76 6a 6f 68 6f 6a 67 57 5d 54 53 57 53 4a 3a 3c 3b 37 38 19 0d 09 0b 19 19 26 2e 33 43 44 5a 58 63 61 6c 72 76 76 7f 7f 86 97 99 ab ac b4 b4 c2 c2 ca d0 d1 da c1 ba a0 9b 98 8d 8a 86 87 82 7b 7a 79 75 73 77 77 6d 6e 68 66 68 5f 57 52 55 5a 58 5f 5e 59 5f 69 64 65 5b 5e 5a 5f 59 5b 5b 50 5e 56 63 55 58 5d 57 61 56 5e 61 5e 58 56 51 55 5b 5c 5b 58 59 50 58 55 58 50 54 61 60 62 5d 58 5a 4e 50 4b 49 4b 56 4e 4d 53 4c 4d 4a 43 53 4d 4c 41 46 3e 29 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 07 03 0a 08 0d 12 20 26 24 25 2a 35 38 39 44 4d 5e 6b 71 6a 5e 53 51 54 51 53 57 57 58 56 53 51 53 4d 59 57 54 54 4f 4e 5d 50 50 55 53 52 51 55 56 53 5a 53 52 4e 52 54 59 55 59 52 64 5f 5a 5a 60 5a 5f 5e 64 59 5e 65 6b 67 61 66 61 5d 59 65 64 63 6b 61 64 6a 64 64 67 6b 69 6c 6b 6b 78 79 75 73 70 74 76 75 6d 73 66 69 67 6b 68 60 60 54 59 52 51 4c 3f 3f 32 3f 37 20 10 0a 0f 16 10 18 17 2a 32 40 44 4c 5b 67 65 6c 67 72 74 7a 81 7f 91 90 96 a7 a8 a6 af ad b4 bb b7 b3 ab 9f 92 94 84 89 85 81 7c 77 77 75 73 79 70 74 6c 69 6f 63 66 60 56 55 5f 54 60 5b 5a 63 60 64 60 5e 60 61 60 5d 52 52 61 59 5e 59 5f 5b 55 63 61 56 5f 59 5a 5b 58 52 4b 55 5a 5b 58 55 4a 49 54 4d 54 57 57 58 5a 50 5a 54 5a 58 52 58 50 54 58 50 53 51 46 49 49 4c 53 4c 44 3e 42 32 21 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0b 1e 20 21 2a 2a 2c 31 3f 3b 49 44 49 65 65 60 5c 52 50 54 59 57 53 49 52 50 50 54 53 55 50 5e 50 56 58 57 50 4e 5a 56 54 5b 4c 58 55 55 53 55 52 52 56 52 54 5b 56 60 56 57 5b 61 59 57 5f 63 62 5c 60 64 64 5f 5c 5f 5a 61 60 65 65 67 69 60 65 62 67 6d 69 70 66 6a 68 68 6e 73 72 6a 6d 74 74 6c 7c 71 6d 71 65 65 5c 66 59 60 5a 51 4c 47 47 3b 3f 37 37 27 10 07 09 0c 12 14 1d 1d 25 2d 34 43 4d 54 60 58 64 73 66 73 72 76 83 85 84 8f 92 95 88 9e a1 ab a2 a0 9b 86 8d 8a 84 76 76 79 7c 77 72 75 6c 71 75 6f 6e 67 74 69 65 62 5e 58 5d 5f 60 61 5c 61 64 6b 64 54 68 62 5e 62 5f 58 69 5f 5d 60 5f 55 56 5d 55 56 5e 54 5d 5f 56 51 4e 57 50 55 50 4e 50 4c 44 56 59 55 55 59 5e 5b 5b 58 55 54 51 57 4d 58 4c 52 4e 52 4c 4e 4d 51 51 4a 41 44 3a 2e 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 0b 12 1b 1a 2a 23 2d 2d 38 34 38 40 4d 4d 64 5c 52 59 58 51 4e 54 50 53 51 4b 4f 4d 4a 5a 57 57 56 4a 4f 57 54 5a 54 56 55 4f 56 59 58
 5a 56 53 56 5b 57 55 59 5a 5c 56 56 5c 5f 5e 6b 60 5f 5d 61 64 5e 5b 5d 62 60 57 5b 5d 5f 64 5c 60 5d 5a 69 5d 69 5f 65 69 67 69 6b 6c 6d 72 6c 76 71 71 72 74 72 69 6d 6e 66 6d 69 55 62 5b 5c 60 53 4f 43 3c 39 3b 3d 20 0c 0d 08 10 12 13 19 16 23 2f 31 30 3a 47 4d 61 5c 5d 58 60 66 6b 72 73 73 7e 77 7b 83 84 92 98 9c 93 8f 7d 80 7f 7c 7c 78 72 77 79 6d 6e 6e 69 6a 66 68 6b 72 5f 75 61 6c 64 6a 64 68 69 69 67 5c 64 66 63 61 64 64 65 64 61 5f 5f 60 67 57 5e 58 53 5b 58 5b 4c 54 64 56 55 49 54 54 4f 48 4f 4c 53 50 48 50 55 4d 59 62 52 5b 5d 52 58 46 50 52 56 4b 4f 4c 52 53 4d 4d 55 47 49 4a 42 3c 23 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 07 06 05 09 19 1d 2a 24 26 31 2c 3c 3b 3f 47 4e 52 4d 4f 54 52 4f 4f 56 51 4e 49 53 52 4e 48 4b 52 56 56 52 50 57 58 51 51 55 48 4c 4b 4a 52 52 59 53 54 4f 4f 50 5a 5f 50 5f 57 57 62 5d 61 63 5f 66 60 56 66 62 61 57 59 5e 59 56 56 59 57 60 5f 62 64 5d 65 63 5d 6a 64 66 70 73 6d 70 6f 71 6b 79 70 6e 72 78 70 71 68 6b 63 67 59 62 65 62 4e 3f 46 44 40 3e 33 19 04 06 09 03 05 0d 0d 13 1d 1b 27 34 35 44 4a 49 5b 57 55 52 5f 5d 61 5d 65 69 6c 72 6a 70 80 8e 87 89 8a 78 7e 7b 7b 70 77 75 78 6c 69 6a 65 6b 6e 6c 70 60 65 61 6a 68 65 66 62 62 62 66 66 5b 65 63 64 69 66 66 6a 73 61 60 64 59 5d 5a 51 50 53 5b 60 57 51 53 58 61 5f 4f 52 4a 4e 4c 4b 4e 49 51 4e 49 4f 56 5a 5c 52 5e 59 4e 5b 55 4e 53 4f 52 4d 4c 4e 4f 46 59 4c 4f 50 48 49 39 32 18 06 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 0d 14 1f 22 2a 21 29 33 30 3e 47 4b 4e 4b 57 50 50 4b 54 52 57 56 4d 50 4a 54 4d 4b 4e 5a 53 55 55 55 5a 55 4e 50 52 51 4d 4f 50 54 4f 58 52 4b 4f 53 5b 56 4e 5a 49 58 58 59 67 61 62 5e 61 5c 54 5a 5d 58 58 5c 5b 59 54 59 5c 64 66 65 5e 5f 5d 5d 67 65 63 66 67 6c 6e 6b 63 72 74 67 74 71 73 6c 6b 6f 72 6f 70 6f 64 69 5a 65 5b 56 49 43 41 42 48 3a 23 10 11 0a 06 07 06 0f 0f 19 19 23 23 2b 3d 41 46 4d 45 4b 4b 54 55 5a 56 5e 5d 60 5b 67 68 73 81 80 7d 75 72 7e 7c 72 6e 67 72 6e 66 6c 61 65 64 69 69 68 62 60 60 6d 5b 5f 5b 65 5d 5f 5c 6e 69 67 71 62 6a 69 68 6c 66 61 58 5d 5d 59 5a 5a 50 56 50 57 54 58 5d 62 68 58 52 52 48 4f 48 48 4d 43 4c 44 4c 4d 5b 54 59 5c 5f 54 5d 5b 53 51 44 4d 47 4a 4e 4c 4f 50 51 4b 56 4e 47 3c 34 25 18 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 04 06 05 03 00 06 0a 09 1d 0d 1f 26 26 38 31 32 3b 43 44 4d 4f 56 4e 53 51 50 53 54 52 49 4e 57 50 50 54 4d 4a 52 53 55 51 59 4f 52 52 51 4c 4e 4d 52 52
 54 4b 4f 4b 58 4f 48 54 4f 55 5a 58 56 5f 56 52 5e 5d 5d 5c 5d 5d 5f 53 5e 5c 63 55 56 5a 55 62 58 5a 5b 5d 5a 61 63 5e 5f 5f 66 69 6c 6a 70 6f 6d 6f 74 6b 76 6d 72 72 6e 6e 71 67 61 64 66 68 5d 57 44 49 40 4e 40 3b 28 11 06 06 0a 02 0a 09 13 16 11 19 1d 21 28 30 35 46 42 48 4a 47 4f 54 55 52 58 5a 50 5d 5a 5d 7a 82 75 72 6f 71 71 6a 6e 6b 72 6e 6c 69 6d 6c 6d 67 63 68 63 5f 63 61 5e 60 5d 56 5f 5f 5f 64 6c 67 6a 6f 66 64 60 58 58 56 55 57 59 5e 5c 56 51 53 58 58 59 5f 57 62 6b 5f 53 44 42 49 4a 49 4a 46 4b 49 4f 60 50 4e 52 5c 5b 5e 4f 59 4f 47 52 47 51 46 4e 45 4f 50 4e 51 4d 50 45 3b 2d 1e 0f 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 04 06 05 03 08 13 1c 24 2b 25 32 32 3c 40 43 49 4c 52 4e 47 56 50 4a 55 52 50 4d 49 53 4a 4a 4d 56 52 51 4f 50 56 54 4e 50 4c 4f 45 49 47 53 4a 4b 4c 47 4f 52 4b 58 51 54 57 56 52 4a 5d 55 57 56 56 5a 5c 51 59 57 55 5b 53 54 4d 57 65 5d 5e 5d 54 53 67 60 64 5b 5f 64 6c 6b 68 63 6c 6a 71 6f 6d 72 6f 6b 70 71 6d 6a 6c 64 61 60 65 6a 66 4f 48 40 3e 38 42 3b 19 11 06 05 03 04 06 0b 0b 0a 13 14 10 21 2a 29 2c 39 34 3e 4b 41 45 44 45 4b 4c 4b 4a 55 51 5f 6d 77 71 6d 6a 70 71 64 6f 65 68 6f 67 67 69 60 5e 67 65 64 53 67 55 62 56 56 53 51 4d 56 5d 60 6a 74 6f 64 58 5e 4b 4a 59 4d 4d 57 52 54 55 57 5c 50 56 50 57 5a 5f 5d 57 55 4e 4b 42 45 44 49 48 4e 4a 4a 4d 43 54 4d 53 5c 57 51 52 4f 53 48 47 4d 4b 4f 4a 4d 57 4b 4a 4f 4b 4d 40 34 22 0c 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 13 1e 1e 1a 24 2d 2e 32 31 39 3a 49 43 3d 46 35 40 3c 3d 3a 38 3a 38 41 47 38 41 40 42 49 3e 44 40 3a 40 45 40 44 45 48 41 47 3e 39 40 3a 3e 43 40 4d 43 45 4a 45 4a 4c 4c 52 4e 50 42 4e 43 46 4c 49 47 45 41 4d 46 4d 4b 42 50 51 4c 4c 53 48 49 4c 50 55 5f 4f 55 55 59 54 59 5a 55 58 57 5e 56 4c 55 51 53 5b 4e 45 3e 36 3d 2e 2a 32 34 2a 1f 01 06 05 03 00 06 05 03 00 06 05 04 0b 06 11 10 1c 1e 25 24 21 28 2d 33 30 38 32 30 35 2e 3d 54 5a 52 54 59 5a 54 54 4f 5e 54 58 53 57 57 57 57 5a 5d 54 53 54 4d 4a 4c 4a 43 48 3e 4f 45 46 46 43 48 4d 53 4b 4c 4f 4d 4e 42 47 44 4b 47 42 51 41 4c 51 43 4c 46 4d 4a 4e 4a 46 47 4c 45 44 47 51 4b 4c 44 43 44 47 4b 4f 52 54 45 49 42 43 46 42 49 40 42 44 45 43 46 41 45 45 43 3f 2b 15 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 23 20 2a 24 2f 33 34 3a 3d 3f 46 45 40 40 3e 3e 38 3e 3d 3a 3d 44 40 36 41 44 3f 47 48 47 4c 41 42 43 45 3a 40 41 43
 3c 42 41 48 45 43 41 43 45 46 44 48 4c 45 48 49 50 52 4b 4d 49 4d 53 45 53 48 4c 47 41 46 47 4e 4e 43 49 4d 4d 54 4c 4a 52 50 4e 5a 59 50 55 55 5b 58 5c 57 59 55 60 57 56 56 5a 55 56 57 52 3f 47 40 3a 3a 32 34 2f 2f 1f 08 06 05 03 00 06 05 03 01 06 05 03 09 06 05 0b 0f 1b 19 20 1f 2f 27 31 2b 30 28 31 2d 32 37 4f 50 53 54 53 54 53 48 58 52 5d 5d 55 5b 5e 59 5b 5c 52 5b 52 4e 51 49 49 47 45 47 41 43 42 44 44 4b 4b 50 4c 44 4f 42 46 4f 49 47 45 4d 4c 4f 49 4e 4c 43 4a 4e 42 4e 49 48 4e 4b 4e 47 47 50 4c 52 4e 48 46 49 3f 4b 4e 47 54 4e 48 50 4e 4e 4a 41 4d 46 41 4b 42 49 4a 43 49 46 3b 39 29 15 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 11 21 25 2a 25 31 33 40 3f 42 3f 3e 3f 41 3f 40 3e 39 34 37 41 3a 35 3c 3d 44 46 44 41 3e 41 40 42 40 45 3e 44 42 42 40 44 35 41 3e 42 3c 40 40 3e 3c 3e 41 4c 45 4c 49 48 4a 4b 4a 49 49 49 4a 4c 52 48 3d 3b 48 4a 42 46 4a 48 4d 49 55 4d 52 52 50 53 50 56 5b 56 5a 53 55 56 55 5c 56 55 52 5b 5b 56 51 62 55 4c 41 3d 33 35 2f 30 2b 2f 20 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 0b 14 12 14 1c 25 24 2f 27 2c 2c 27 2a 28 48 4c 53 58 50 54 56 55 55 54 53 52 53 5e 52 54 5c 5a 54 50 4b 52 46 4d 49 3e 45 40 3d 43 44 3e 41 43 48 4d 4d 4c 43 44 4a 49 44 45 48 48 4d 4e 45 4f 40 43 43 4a 43 4f 42 49 4d 4b 4c 49 4d 4e 4f 4f 4c 49 46 42 49 4e 49 4b 4e 53 4e 4a 49 45 4d 4a 42 42 3e 3e 48 43 47 44 45 3e 3d 36 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 11 1f 17 1a 2b 28 30 36 33 44 3d 40 39 37 3c 41 41 3b 41 36 36 44 38 38 44 3f 43 3e 3f 38 35 44 42 39 47 3e 40 3e 44 41 3e 36 3d 3f 40 32 41 3b 51 3d 41 48 51 45 44 41 47 43 4b 4d 44 48 45 4b 4b 52 37 46 42 4b 4e 43 44 45 51 46 48 4a 4e 56 51 4f 56 52 5a 4f 5a 5a 53 54 58 4e 5a 53 56 5b 56 55 56 56 58 5e 50 44 3d 35 34 30 2d 36 2f 1a 08 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 04 06 08 06 10 15 17 1c 21 22 25 1c 26 22 2d 3d 49 50 4e 40 54 4b 4a 53 55 51 54 4a 50 55 55 58 50 55 56 4d 45 3f 48 40 47 4c 46 47 45 49 41 52 45 4a 4d 49 4a 46 46 46 46 4b 4b 3b 3e 45 3e 4a 3e 4b 48 45 49 4d 4a 43 45 49 5b 52 4d 49 44 4b 48 45 47 3e 41 43 41 4a 4b 4a 52 42 49 47 47 49 3f 49 49 3d 47 40 47 48 46 42 44 41 28 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 13 24 2a 2b 2c 34 39 42 36 3b 3a 41 3a 3f 40 3f 3e 3c 39 44 45 40 3c 41 3b 44 44 3d 40 3f 3d 3d 3f 45 37 37 38 42
 3d 41 3e 3e 3e 41 3d 4b 3f 41 4c 49 3f 44 48 4c 49 4b 41 54 4a 50 48 40 4b 49 47 4b 47 48 4b 4e 4c 47 3f 4a 41 4c 50 4a 50 4c 52 51 4f 56 51 57 54 58 59 5c 51 5f 56 54 55 50 5d 52 57 52 60 54 47 3f 41 38 41 36 2f 34 26 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 09 04 04 12 0e 13 17 1c 1b 1e 1f 1b 26 44 53 44 47 45 4e 4f 49 4d 4e 51 58 4d 4f 51 54 55 4e 47 50 49 51 42 45 45 43 43 4a 48 45 46 45 49 49 46 48 45 45 45 4d 45 46 4a 4e 46 46 4d 45 44 3b 48 44 3e 40 40 48 4b 4b 58 5b 52 4d 48 41 42 4b 4a 4a 41 44 44 47 41 46 49 47 47 4b 41 46 48 41 3e 45 43 49 3d 43 49 42 42 42 38 1d 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 11 1b 1e 2b 2f 2c 36 3d 30 3b 3e 3b 34 3d 46 41 3a 3e 3c 3a 3c 44 45 3a 42 42 39 38 37 3f 3c 44 3a 3e 3a 37 40 3a 3b 43 3e 3d 3d 35 36 44 3c 44 40 47 44 49 4d 45 4b 46 41 45 43 4c 4a 47 4b 44 42 4e 4c 49 4f 46 4c 4d 49 4b 4d 43 47 4a 53 4f 53 54 48 53 50 4e 5a 54 55 54 47 57 57 5a 4b 55 5b 54 57 58 5d 5b 46 47 3e 38 34 35 3a 37 23 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0e 0c 16 10 17 13 17 19 1c 37 40 40 47 44 4d 4b 46 47 51 47 52 51 52 4f 50 56 50 4d 50 4d 47 41 47 47 4c 49 47 45 49 48 45 44 47 48 49 46 45 44 45 45 49 47 47 44 40 4d 48 47 44 49 40 3f 43 41 40 4b 46 49 49 4b 49 3e 46 47 42 44 40 47 43 45 45 43 4f 4a 4d 3f 3e 47 46 40 46 45 48 39 4b 4e 44 46 44 40 35 21 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 15 23 27 28 3a 36 3d 35 39 3d 37 42 3a 35 3c 3c 3a 44 3a 43 32 34 3d 35 45 3d 3c 35 39 37 37 3c 35 3a 38 40 35 44 36 3f 35 31 37 39 38 3a 41 3b 41 42 3b 4e 43 46 47 4c 3f 48 47 49 49 49 3e 50 41 44 44 49 45 46 4e 4a 52 43 47 4e 4a 4f 49 46 48 4d 51 4e 57 4f 54 51 4c 55 50 4e 52 53 5a 59 53 4f 5b 5e 53 49 40 3b 38 35 40 2b 25 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 07 0e 13 17 16 14 29 42 37 4d 3c 45 41 41 49 47 4c 4f 4f 49 4f 48 49 49 43 52 49 49 47 44 4d 42 47 46 46 48 4a 43 45 41 44 51 49 44 4c 50 41 45 4a 4c 45 45 47 42 43 3f 4a 44 3e 41 3f 45 42 44 4c 4a 44 46 51 45 49 47 44 44 38 41 40 3f 45 43 39 49 39 3e 48 45 44 41 40 47 44 4a 47 3d 4c 35 35 32 1a 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 16 23 27 27 34 40 3e 3c 3b 3f 36 3c 40 36 40 3b 3c 44 3f 46 33 3c 39 38 3f 3f 37 32 40 37 35 39 34 45 3e 44
 33 39 39 3c 3f 3c 34 3e 43 3c 45 3e 3f 45 47 45 47 42 45 4a 4b 48 43 52 4f 48 49 43 49 4a 4d 42 4b 4c 45 4e 42 48 4b 4f 51 48 4a 44 4f 4e 4a 51 57 52 55 53 50 59 58 4f 52 5a 56 54 52 5e 64 62 51 49 44 40 40 3d 3c 3a 2b 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 0f 08 11 07 18 2d 41 3f 40 3f 46 4c 49 49 49 50 4f 52 4f 49 52 45 49 49 48 44 47 45 4f 45 45 42 42 4d 4c 43 49 46 40 48 4c 47 41 48 4a 54 4f 4a 46 46 42 4c 50 46 44 3b 44 42 40 3e 47 43 42 47 3e 3e 4a 4a 3d 42 4b 3a 47 45 4a 45 46 46 4b 3f 48 43 43 4a 43 45 46 44 48 43 45 4e 44 49 3f 38 25 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 0c 21 34 33 32 32 3f 3a 42 40 38 3c 39 3a 3f 41 3e 31 33 39 3b 38 3a 30 39 36 3e 35 43 3a 40 3e 3e 3f 36 3c 3d 38 3b 40 38 33 3c 38 38 38 40 40 38 41 43 43 44 52 46 48 4d 4d 4a 49 4a 49 48 45 43 4c 4a 52 4a 43 43 48 4a 52 4b 4d 4a 4f 4d 4c 4f 4d 4d 54 4c 53 5a 52 52 54 55 52 54 59 60 55 5b 61 5b 5a 49 42 3f 3f 38 38 3d 25 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 0f 09 09 1d 38 3b 42 42 43 4d 40 46 49 41 55 4c 48 45 50 4a 49 45 46 48 48 41 46 45 4b 45 43 4e 4f 48 4b 44 48 47 51 49 4b 42 50 4c 42 45 49 46 3a 41 44 3f 3d 4b 48 44 3e 3f 45 3e 3f 4a 42 39 3c 49 45 47 3f 43 49 38 45 40 43 44 4d 47 4c 3f 45 3b 3c 4a 3a 3d 41 42 45 41 41 45 36 2f 1a 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 18 26 31 34 40 3d 2f 38 38 3e 36 33 38 40 3f 35 3f 3b 3b 32 3f 3a 33 34 3b 41 38 36 41 44 37 39 37 34 37 37 37 3a 33 35 3e 36 41 3e 39 39 3f 3e 3b 42 44 45 47 46 42 54 55 4e 55 50 46 45 48 4b 4d 54 50 40 45 4b 4c 42 46 47 45 4e 4e 49 4c 4d 42 51 54 50 4f 4f 54 55 52 58 50 56 51 54 56 5a 5c 60 51 50 4b 44 43 42 3c 3c 24 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0a 21 34 3a 37 3f 41 42 44 45 44 4d 42 4c 4d 49 46 48 45 47 41 4b 42 47 4f 4b 4f 47 4b 4d 41 4d 47 3d 44 45 44 41 49 44 45 46 45 44 44 44 49 44 39 45 46 47 3d 43 4a 3a 4c 48 46 45 4b 45 43 45 40 48 41 44 43 3d 44 46 47 42 41 41 44 48 3e 47 3f 40 41 42 46 41 41 43 42 49 3a 22 12 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 1a 22 32 3a 38 35 41 39 3b 3c 30 33 3a 35 3b 37 38 3b 33 34 2b 33 33 36 3c 3f 3a 3b 3e 42 39 3d 3e
 35 3a 3f 2f 38 33 3a 3c 3d 36 3f 40 41 3d 39 3e 3d 41 42 46 42 4c 55 4f 52 4a 47 44 47 46 53 3c 27 34 51 4d 48 44 41 47 49 4e 49 45 40 45 45 4b 54 4e 55 4e 4b 4e 52 4d 5a 52 53 54 5a 62 58 58 5c 50 4e 48 41 49 37 42 2f 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 1d 2f 3f 43 3f 3b 45 41 3f 44 3f 48 41 49 4d 4b 3c 4b 4e 44 45 4b 48 48 41 4a 50 47 49 4c 42 42 48 42 4d 45 40 3a 3d 48 4b 41 3e 4c 41 42 48 46 47 48 44 44 42 40 42 4c 3e 44 45 46 49 41 42 40 3d 3d 49 44 46 45 47 4d 43 3a 44 44 44 45 46 41 43 40 42 49 49 44 49 44 3d 2d 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 13 27 2a 35 40 33 39 3a 39 3b 3d 36 3b 33 35 3a 38 39 39 32 39 36 3a 3a 39 39 3b 37 39 3e 39 3d 37 35 37 38 3b 3a 3b 3a 3e 39 3c 42 3a 44 3c 34 3e 3f 36 40 3f 47 4b 4c 4b 5b 4c 44 4d 43 4c 47 45 4a 4d 4f 46 43 49 48 47 4d 45 45 49 45 48 4a 44 47 47 48 52 58 59 55 5d 54 5a 59 59 50 5c 60 5e 56 51 52 4f 44 44 43 3a 37 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 33 36 3d 38 3f 44 34 43 42 3f 46 43 4e 4b 43 45 40 41 3f 42 49 4d 46 4a 4e 4c 45 49 4e 52 48 3e 46 4c 47 47 46 4d 4f 48 47 46 40 3b 49 49 44 3f 43 3b 4d 3e 3e 47 50 3e 45 47 45 4a 43 47 45 3d 41 3d 4f 3d 49 37 48 40 44 4d 47 48 49 4c 3d 41 41 48 41 3e 4e 42 3c 38 26 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 16 2b 2f 35 33 3c 39 3a 41 40 36 3d 38 2f 36 36 39 37 3b 39 38 32 3b 34 3b 2d 3a 3b 37 3d 35 39 36 32 36 33 37 41 34 3a 3b 37 36 34 3f 44 38 3c 40 3f 3f 3a 40 46 43 4d 53 54 47 4c 46 42 52 49 45 40 43 4b 3d 44 47 3f 4c 4c 49 49 41 4c 47 4c 52 4d 4b 49 51 51 4d 56 4f 52 55 52 5a 62 54 5d 59 51 55 48 40 49 3d 3c 30 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 29 38 46 39 40 39 3f 3b 42 3f 49 3e 48 42 43 44 45 48 45 44 4f 40 4a 4a 4a 4b 4b 41 48 44 48 46 44 4d 42 46 42 42 41 48 4c 3f 45 38 43 47 48 43 44 43 45 3f 3e 3f 48 3d 45 3f 42 3e 49 3b 46 39 42 45 40 42 46 42 44 41 46 47 47 3e 43 43 43 43 3a 45 45 3f 48 3d 3d 2f 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 30 28 30 30 3c 36 3b 3e 39 3c 36 34 2f 37 31 38 32 36 30 2b 35 38 3e 38 3c 37 35 38 30 3e 3b
 33 35 42 34 3c 35 39 36 37 3b 37 38 33 41 3f 41 39 3a 3c 47 36 3e 38 40 4a 51 48 41 49 42 47 49 4a 43 45 4b 42 41 41 44 40 47 50 4e 47 45 3e 45 4b 50 4d 50 4c 53 4b 54 56 51 56 5f 5c 5d 61 55 52 4e 46 50 4e 42 55 40 38 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 31 39 3d 35 40 3e 43 3e 41 3a 3e 45 47 46 43 46 4b 49 45 45 48 43 45 48 47 41 4a 48 4c 49 47 46 4a 48 44 3f 43 45 43 3b 47 47 47 3f 44 3f 3e 45 4b 40 43 4b 46 4d 42 45 47 46 45 3f 3a 43 46 41 41 48 47 3c 49 44 44 45 4a 49 4a 48 40 42 3f 48 44 47 46 45 44 3a 36 21 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 28 35 3a 3e 3c 38 3f 39 3b 33 38 3b 31 2e 36 33 32 31 2e 3a 35 3c 31 3a 37 37 3c 35 3b 3d 3a 35 3d 36 37 35 38 42 3a 37 3b 41 3b 3b 39 41 3d 43 39 3f 3f 3d 41 44 45 3d 4d 52 49 49 4b 4b 50 4d 55 4c 43 4c 47 51 54 46 4a 49 45 44 51 44 41 41 4f 51 55 55 55 53 57 53 56 5e 52 58 5e 57 54 59 4b 52 50 4c 4b 4b 39 21 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 2e 30 3f 3c 44 37 47 3e 3f 41 54 42 40 46 49 40 48 46 49 4c 50 4f 53 46 4b 4f 47 4a 47 44 46 49 4a 46 44 45 3d 47 42 41 4c 42 3f 40 47 3c 44 49 45 51 45 40 48 45 45 3b 41 43 45 41 46 47 42 49 4a 4c 49 41 4a 40 4b 45 49 43 43 45 4a 48 4b 4c 46 44 44 43 47 3a 2b 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0f 25 39 38 3a 3b 3b 35 2b 37 2b 33 3b 34 3a 33 3a 2f 39 31 37 33 38 35 3b 3c 39 3b 34 41 3d 32 35 39 36 3a 3b 3c 33 3b 3f 39 3a 3a 38 39 40 38 45 41 3e 42 41 3f 40 48 4d 57 45 3c 47 4a 57 57 52 4d 48 47 48 49 54 45 40 43 45 4d 49 4b 45 4c 50 4a 48 49 4b 47 4f 54 5c 64 5d 5e 52 59 56 56 49 55 53 4f 55 4a 3c 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 29 30 3d 3e 46 3b 3b 3d 3c 3e 43 44 44 43 52 47 48 49 4c 47 4f 4b 4c 42 4b 3e 49 50 4b 4f 4a 40 4d 45 40 47 46 48 48 48 46 40 47 47 43 4b 47 3e 44 45 4d 3f 40 3e 47 42 41 42 42 3f 44 40 44 42 44 44 50 45 47 49 42 4e 4a 43 4d 40 47 45 49 4e 49 43 4e 44 3f 2e 17 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 2b 33 3a 3e 3a 34 39 40 33 3a 2e 31 35 32 34 36 35 2b 39 32 41 31 36 3a 38 34 33 32
 34 36 3a 2e 3a 35 36 36 3a 36 39 3c 34 3a 38 3b 4a 3c 37 44 3d 3e 46 40 4d 3e 3f 44 47 46 45 47 59 50 54 55 54 48 4c 54 4f 42 4c 40 40 4a 3f 4b 46 43 4c 51 54 4f 51 52 58 52 52 59 5b 5a 51 58 56 5c 57 50 4a 43 47 45 3f 23 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 28 37 44 38 47 47 44 3c 41 44 46 52 4d 53 4e 4a 51 42 46 44 45 46 48 48 46 48 41 4d 46 3f 44 45 4c 4f 4a 3a 42 50 42 45 44 3a 47 43 3a 49 3c 47 44 45 49 3e 4a 45 47 46 45 4b 42 3f 41 3e 41 45 4c 3d 46 45 44 44 42 42 46 53 4c 49 40 49 44 49 49 4d 44 3d 35 26 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 0b 1e 37 2c 37 3b 3f 32 35 37 40 30 36 33 3e 2d 2f 37 2e 37 37 3f 3c 3d 3b 39 39 36 33 3a 3d 37 3e 3a 39 39 39 34 37 3c 36 37 40 39 3d 3a 39 41 45 3f 49 4d 43 44 40 44 45 4c 43 46 45 4b 4b 4c 4f 50 50 53 5c 5a 4b 4b 4c 45 46 47 50 48 4f 49 4f 4b 5a 52 51 4e 59 58 5b 5b 5b 57 5a 53 4f 53 54 57 4d 4b 48 37 26 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 2f 39 41 3c 3a 3c 3e 45 49 4e 4c 52 58 4e 4e 42 4f 4a 52 40 3f 4b 47 44 4c 4a 4f 4a 44 4c 4a 48 4d 47 4e 43 4e 41 49 4b 46 48 43 4c 44 41 44 4b 43 49 42 40 49 3b 49 45 42 51 44 38 3f 40 4f 4d 4c 45 44 3e 48 45 45 4b 46 49 4a 46 46 50 4b 46 44 45 48 3f 2e 1e 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 15 2d 32 34 3d 36 34 3c 39 38 35 2e 3b 38 36 36 31 3a 38 3c 3c 35 3e 3b 38 39 40 32 33 43 3a 3c 3d 3b 38 3b 3e 3a 3a 41 42 3f 39 42 3b 36 3a 3a 36 42 41 47 41 41 49 45 43 46 41 48 4f 50 52 55 59 4f 50 59 5e 53 55 46 49 43 47 47 45 4d 4f 4e 4c 53 4b 54 53 53 54 57 59 56 59 59 57 55 55 4e 4d 4e 55 4e 42 2d 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 27 3b 48 42 3f 42 41 4a 43 50 54 4e 52 4c 4c 41 4b 48 4c 48 3c 4a 47 45 44 45 4d 41 51 49 51 4a 4e 4c 48 4a 47 3c 44 45 48 45 47 3e 3b 4a 47 48 4a 45 3f 44 46 44 42 44 3b 39 45 42 50 3f 48 46 45 40 4b 41 3d 3e 44 54 47 4e 55 49 41 45 3f 40 3e 3d 3e 36 26 16 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 1c 32 2f 39 3b 30 38 35 38 38 39 2f 3c 30 35 33 3b 39 35 3d 38 3f 3f 3e 3b 34 39
 43 3b 37 3a 37 3f 39 3b 36 34 3d 42 34 36 3c 45 3a 40 3d 45 38 42 40 40 44 40 41 46 45 42 41 47 47 4e 4d 51 4b 4d 50 54 56 55 51 48 42 44 45 4b 4b 45 4c 4d 4b 4f 58 51 53 53 59 5d 58 5e 4c 55 4e 56 58 50 49 51 45 49 46 24 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 29 3e 43 42 3f 3f 42 42 52 4a 57 3e 47 46 45 46 41 42 42 41 4a 44 42 47 4a 45 42 40 43 4d 45 46 45 47 42 49 40 41 46 41 3f 41 41 44 3f 44 45 43 3f 3b 3c 3a 46 42 44 4c 45 47 48 3d 3e 3b 41 44 48 44 45 46 43 40 4c 4e 47 4e 46 47 4a 44 45 46 47 44 3b 2f 1f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 23 2f 37 38 36 35 3c 3a 39 3c 38 38 32 35 39 3a 38 3b 37 34 3d 3c 3b 3b 3c 44 38 35 39 35 33 3a 38 38 3a 40 3e 35 32 3f 42 40 40 36 3e 47 3f 3b 46 3d 3f 44 43 48 44 46 43 50 4c 4d 48 48 50 4f 4d 53 54 52 50 47 43 4e 3e 4d 4a 46 46 50 52 53 56 4e 4b 55 50 5b 57 58 5b 57 58 5a 53 55 4f 51 4f 46 3e 2f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 40 4b 40 3e 42 42 49 4d 49 44 3f 45 3e 45 45 46 4c 3f 44 4b 49 4d 48 58 40 45 47 49 4d 4e 46 44 47 3e 42 47 48 49 47 4a 3c 46 41 46 4c 47 44 4a 47 4c 44 43 42 4a 48 3e 43 43 3e 46 40 45 4a 4a 44 4e 43 42 4a 42 40 50 4d 51 46 4d 4f 46 4a 4b 37 3b 1e 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 11 1d 35 32 32 38 2e 39 34 3b 33 2f 3a 3b 33 33 3a 3e 35 3e 3d 3b 3f 36 37 41 42 45 34 37 3c 3e 38 38 3b 40 37 41 3f 40 41 42 43 3f 3e 44 39 42 43 3e 43 40 40 47 45 4d 4d 4b 49 4b 4e 46 4b 4b 4b 52 53 4f 50 4f 49 4f 41 4c 4b 49 48 4d 43 55 4e 54 4d 57 56 56 5d 55 51 49 50 4f 53 51 50 50 4a 4e 46 35 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 26 3d 47 44 42 4a 4c 44 45 3c 43 3f 44 48 44 43 42 48 4e 44 46 4d 48 46 50 48 4a 45 4f 46 4e 3f 4b 49 3f 43 40 3e 47 42 49 4b 43 45 43 49 47 3d 43 44 44 45 44 41 3e 48 44 44 42 3c 4d 47 40 49 46 3b 46 44 47 45 4d 4a 49 50 4f 48 4d 44 44 4c 41 3d 2a 11 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 21 26 2e 39 3b 37 34 39 38 38 37 33 38 2c 31 33 3b 37 36 3a 41 40 3b 3c 37
 32 3d 34 37 36 38 39 3e 3d 46 3b 3b 3e 3e 3d 3d 3a 39 46 45 3e 42 43 3c 3b 3e 38 41 3d 46 41 45 46 45 46 49 48 50 4c 54 4f 4f 4d 4a 45 49 47 4a 49 43 4b 46 4d 4c 4a 4d 50 53 59 51 54 58 59 4d 54 4b 5a 47 4a 4e 4d 43 3d 33 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 20 35 49 41 4b 47 4b 45 41 43 43 48 46 41 49 4a 46 45 44 41 47 47 45 4c 4b 3f 4e 49 46 42 48 48 46 44 45 40 40 47 3f 43 42 47 46 44 40 3c 51 40 3e 45 47 3e 41 42 48 4b 46 40 3a 3e 3b 45 44 42 43 3f 43 3a 43 47 47 47 43 49 54 4c 4c 46 41 3d 3e 26 1f 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 20 2a 34 2f 37 32 3b 30 34 39 39 36 3e 33 35 3b 39 39 41 42 36 36 39 30 3a 3b 34 34 34 38 3d 35 40 37 3a 39 38 3d 3d 39 3d 3c 44 42 43 3f 41 3d 3f 3d 45 44 42 45 4a 40 4a 4c 4b 4e 40 4a 4d 4f 51 4f 54 4d 43 49 52 4b 55 49 4e 4f 50 4d 4b 44 4c 5b 57 58 5a 53 52 54 4d 4a 55 4e 51 55 4f 4a 3d 36 15 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 2a 4d 51 4a 49 53 46 47 48 47 44 46 40 41 4a 44 43 45 45 44 47 40 45 42 43 4b 3f 49 44 4f 4c 3d 44 3e 4a 3c 3c 45 3f 45 41 4a 4a 4c 49 43 44 44 42 3f 42 41 4e 45 49 42 3b 45 3e 3e 46 42 40 49 4d 44 46 40 44 4a 47 47 4f 49 55 4a 4a 43 44 3b 3c 1d 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 16 24 2b 2c 35 37 36 45 3a 3e 3b 33 31 38 35 40 37 35 44 39 40 41 36 39 37 3f 33 41 38 38 39 3b 3f 48 36 3c 39 3d 41 44 42 3f 42 3b 3b 45 3d 3f 43 41 49 41 40 3c 40 4d 44 47 51 45 4d 47 46 45 4c 56 4a 52 44 46 4d 48 4d 52 4a 4d 4e 56 4e 4d 4c 47 55 4d 4f 55 4e 56 52 51 51 4d 4c 50 48 4b 3b 35 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 31 59 56 49 49 3e 44 45 47 42 3e 37 48 3e 47 45 4d 49 4c 44 49 43 48 42 4b 45 44 49 48 46 43 47 49 3e 44 44 45 4e 43 3f 47 43 43 41 3e 42 44 44 3e 3d 44 3a 41 45 42 3e 3c 43 41 44 4d 45 42 41 52 4b 47 45 45 43 45 47 49 47 4b 4e 4a 43 43 3e 30 16 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 20 29 38 3b 44 3b 34 35 33 3a 32 38 30 33 3a 35 39 34 3a 34 31 38 38
 3f 38 3f 39 3d 3d 36 3a 37 33 3e 42 3b 3b 3a 3d 4a 39 45 40 41 39 3d 44 3f 44 45 3f 3d 3d 3e 3f 45 3e 45 46 44 45 47 48 4b 53 52 49 47 42 44 47 45 43 4b 48 4b 53 47 46 47 4b 43 58 52 50 47 4d 50 52 51 4e 53 4d 45 4b 49 3a 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 56 57 50 49 3f 44 43 41 38 44 44 3a 45 42 48 49 3f 43 3d 49 4a 43 4a 4a 45 40 42 46 43 49 3b 39 44 43 42 3e 46 46 47 39 44 43 3c 42 43 3e 40 48 3c 40 3f 41 37 45 3b 46 43 3f 48 47 42 44 38 42 47 42 43 4b 4c 4f 4b 4d 40 4e 4c 3d 48 3d 30 1e 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 22 2d 34 36 3b 34 3b 43 3a 39 31 38 3a 3b 35 39 40 3a 41 3e 38 35 3c 36 3f 3b 37 3a 3c 37 36 42 3d 35 3f 41 3e 3f 41 43 45 3f 3a 47 41 44 46 3d 45 49 3b 41 4a 41 48 42 46 47 47 45 51 50 47 49 4c 44 4d 4c 46 50 48 4e 4e 47 4e 52 49 4d 4f 50 4e 54 50 51 55 4c 53 50 4d 48 47 4f 56 4a 44 32 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 44 45 3f 48 41 3e 40 3d 40 44 48 4c 40 49 48 43 46 44 45 4d 44 4a 49 4d 46 45 46 4e 48 42 3a 46 41 3c 45 40 4d 48 47 49 3b 3f 43 3c 41 46 41 41 41 3c 41 48 41 48 3f 39 4a 4a 47 40 3e 41 51 46 43 43 48 49 4c 50 49 4f 4d 4d 44 3d 3b 3c 26 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 15 2c 32 36 38 34 37 3b 32 33 32 36 36 35 3c 3d 36 38 38 3a 3a 39 3c 3e 37 3f 37 3f 36 3d 35 3f 40 3a 3f 43 3b 49 3d 3b 40 4b 36 39 4a 42 45 4f 3d 4b 44 40 3c 42 4c 41 4d 48 41 46 44 49 4e 49 4b 48 43 47 44 51 48 4b 50 43 4e 50 4a 47 4d 4d 4f 58 4c 5b 54 4c 4c 4d 4c 45 48 44 52 49 4a 32 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 3c 44 40 41 48 41 43 3f 40 41 40 45 46 49 46 42 40 48 40 4c 46 4a 49 49 49 44 4f 4e 49 4a 42 40 48 44 3e 39 43 40 3d 40 3e 3b 49 45 43 44 3e 3a 42 44 32 4a 41 44 46 3c 3f 46 41 41 42 45 49 45 48 44 49 45 4a 49 4b 50 53 4b 46 42 3c 27 1c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 22 24 2d 31 3b 43 31 40 39 3c 36 31 3a 34 36 32 30 31 38 3d 38
 40 35 35 35 3f 40 3a 34 3b 3b 3e 3e 3d 41 44 43 41 3f 3f 41 36 49 41 41 3f 43 48 44 41 40 48 43 3a 44 43 43 4b 45 43 4a 46 4b 48 4e 46 43 4b 4c 4c 44 48 4b 45 4a 4a 4b 4b 48 4c 4e 4d 52 4b 4a 4b 48 4a 4c 50 4a 51 46 41 39 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 17 37 44 3f 3e 4b 3b 3d 47 3c 42 47 44 4b 45 43 47 48 49 39 42 4a 4f 40 4e 46 43 47 43 42 43 3d 3d 40 44 44 3e 41 46 3f 4a 45 43 3c 45 49 45 48 3d 3f 43 3e 3e 46 44 44 3e 45 3d 3d 47 47 42 44 44 4d 45 41 45 49 43 4d 4f 49 50 43 31 2b 24 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0e 15 24 26 2f 39 3b 42 3a 3d 34 36 36 38 38 3a 3a 3c 3b 36 33 39 3e 3f 3b 30 34 39 39 3b 3a 3a 3e 36 3e 3b 44 44 3f 40 37 46 3b 49 3f 3a 3a 3c 39 40 3d 41 3a 44 41 3d 44 41 47 47 48 48 47 3c 4e 41 4b 4f 4c 49 4a 4a 43 47 48 40 47 46 4f 4d 4e 4e 4a 4b 4c 48 49 45 54 53 4d 4a 4c 46 47 33 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 35 44 35 3b 3c 40 42 3f 3f 4a 41 42 3e 44 46 48 3e 48 48 4d 45 4b 45 48 46 4a 48 4a 44 49 3e 3d 49 45 44 3c 44 40 3d 3f 40 44 3d 3b 42 3f 47 3e 3e 45 3e 3a 3e 41 41 3d 47 3f 3f 45 45 44 4f 4b 47 45 47 47 4c 42 45 4b 44 49 3b 38 23 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 27 35 3a 39 39 3c 3b 39 37 3a 37 39 3b 3f 39 37 39 41 3c 3a 38 42 3e 38 36 38 3a 3b 3c 3b 3e 43 3a 3e 44 47 3e 40 3e 43 40 41 3e 3c 43 39 44 3d 3b 41 43 46 3e 40 47 46 40 42 45 4a 4c 46 44 4e 44 3e 49 49 4c 44 47 4b 48 42 45 4d 4b 4e 4e 47 4e 48 43 49 4d 48 45 45 4b 45 48 48 3b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 2c 43 38 3c 36 38 3f 46 3d 45 3e 3c 47 48 50 44 4e 4d 44 46 43 4f 4e 4e 49 44 44 45 46 47 3f 3e 4a 44 3a 42 3c 44 45 42 46 40 3b 44 3d 49 42 44 3b 40 3d 40 47 45 48 4c 3f 43 41 4a 49 49 40 47 44 46 46 4f 45 4b 49 49 43 41 37 29 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 20 2d 35 3e 32 39 3f 38 3c 37 35 39 44 3f 37 42 39 38 3f
 42 39 3e 40 36 3b 3e 39 40 41 40 3e 40 3b 3c 44 48 42 3d 44 42 44 3b 37 48 40 41 3e 38 44 3e 3e 41 43 3d 43 3e 44 3f 44 4c 3d 3d 40 3d 40 41 49 3f 4b 47 44 4f 41 4b 52 4a 4d 49 48 51 4e 4a 48 48 4e 4c 4c 4c 43 4e 48 41 3b 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 2d 3c 41 3f 45 43 3c 46 40 46 3c 42 44 46 4c 46 50 47 4a 4f 48 49 48 4f 4b 44 4a 42 43 43 3c 3a 38 3d 44 46 3c 44 3f 3d 41 3d 43 43 41 45 3d 45 3d 3d 3c 44 3a 45 40 3b 41 3c 42 43 48 44 43 41 3e 3d 40 3d 4b 43 45 47 41 3a 2c 12 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0c 21 31 30 39 3e 3a 37 36 36 3c 41 3c 35 43 31 31 40 32 3e 3b 37 38 3e 34 3c 3d 39 3e 3b 45 36 43 43 45 3d 44 47 3f 40 42 45 3f 40 3d 35 3d 37 3d 3f 40 40 3c 41 42 3f 40 40 41 43 3c 49 44 41 4c 42 45 3d 41 3d 43 47 49 48 46 4c 46 4d 4d 46 45 4a 45 4d 42 49 42 46 46 44 44 38 3d 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 28 34 3c 3d 41 42 3d 3e 46 40 46 47 50 48 46 49 44 4a 50 50 46 45 48 49 44 42 44 4c 42 3c 3f 3c 46 40 3f 38 41 45 40 41 4a 46 43 39 3e 3c 3a 46 45 44 44 42 40 4b 3b 41 3d 40 40 47 43 41 45 49 42 45 39 4a 3e 3f 3a 48 3d 30 1e 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 15 22 34 33 3d 3b 3b 38 3f 3a 39 3f 3b 41 3e 3e 37 3c 3b 40 3f 3e 3d 3e 3e 3c 3c 40 42 44 39 49 40 47 44 3c 4a 44 3b 43 41 3d 45 3b 3d 47 34 3e 42 3d 44 45 42 3a 3c 36 46 41 40 42 43 3f 38 49 48 42 49 46 41 48 3a 47 4a 40 44 4d 52 47 47 4f 4c 49 4c 4f 4d 4d 4a 42 47 48 40 40 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 32 3d 35 41 41 3e 44 3d 50 4d 49 48 3f 41 4c 45 4d 4f 46 49 41 43 48 4c 4d 44 43 43 42 42 40 3d 3c 39 3b 3e 49 45 49 3f 3c 41 40 41 45 41 3f 43 45 3a 43 3e 40 40 3e 3e 40 45 40 47 45 42 43 4c 4a 4a 44 4d 4a 42 41 37 2a 20 0d 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 2a 34 3c 39 37 36 3a 35 47 37 36 3c 36 30 35 42
 39 41 32 36 38 3d 33 3f 3f 3a 40 3d 42 46 45 3b 3e 44 3c 3e 44 41 42 3e 3d 3a 36 3e 3e 3e 40 42 37 42 41 41 38 3e 42 3c 40 38 42 3b 3e 44 3f 3e 44 41 3f 45 43 46 45 40 48 42 4b 44 41 4a 49 48 4a 46 42 4a 46 42 49 45 41 37 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 29 44 3f 45 3e 40 48 44 48 3e 49 46 42 49 4a 50 48 45 45 4a 45 4a 51 3b 44 43 4b 42 3e 44 37 41 3e 36 3b 46 40 45 40 3d 40 49 3f 3e 3e 44 40 44 3c 44 3d 39 3f 3f 46 3f 44 39 41 47 42 3e 4a 42 45 46 52 4f 47 50 36 2f 1d 12 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 1d 2f 34 39 34 3b 33 3a 44 3a 36 39 36 41 3a 32 3e 3d 3e 3d 38 43 37 3b 3f 3b 3b 3c 3f 43 3d 39 3a 3a 3a 44 42 40 43 32 3d 3c 3c 3a 3b 3b 3a 41 3e 3c 43 40 3a 3e 44 3d 40 44 4a 44 3e 3e 43 43 3b 3f 40 46 45 4a 47 40 47 43 47 49 4b 41 46 46 47 45 46 3d 46 3d 42 46 48 3c 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 2c 42 44 4a 48 43 3b 45 4e 46 4c 47 44 4d 46 55 47 4c 45 44 4c 49 47 4a 39 3e 40 3c 36 43 43 41 3b 3d 42 41 40 3b 3e 41 3c 44 40 3b 3f 3c 41 3e 42 45 3b 3b 37 42 41 44 44 42 3d 3a 47 42 45 4f 45 4c 4f 52 57 3b 37 29 0e 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 2a 34 35 2d 36 3c 35 3b 42 3b 42 39 38 3d 3a 45 41 3d 3b 3a 41 40 40 3b 3e 3a 3e 3d 46 41 3a 41 3b 44 41 3b 40 3e 3c 40 48 35 3f 41 38 3f 3d 39 38 39 42 3a 37 3c 3f 41 3f 39 39 49 3f 44 47 4a 42 41 41 45 48 47 3f 44 3e 51 49 4b 44 41 46 40 46 45 44 3c 44 47 40 3e 3b 1e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 29 3f 3f 44 43 3a 40 46 42 4b 48 4d 56 4b 50 50 46 4b 46 44 4d 44 4a 46 3e 43 49 46 4a 48 46 3b 44 44 41 3b 3e 3c 41 43 3c 41 41 3d 46 3f 42 3e 43 3e 40 38 3b 43 45 3e 43 41 41 46 45 47 52 52 51 47 4d 4e 3a 34 24 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0e 19 24 35 34 38 3e 40 3f 3d 3f 39 3e 41 37 45
 3e 47 36 38 36 45 3d 45 3d 45 34 3c 37 41 43 39 40 41 3f 49 43 39 3d 3f 40 38 3d 3d 37 40 3e 46 49 3d 42 43 39 4a 40 41 43 42 3a 45 4a 42 39 3d 42 40 43 44 41 45 44 39 4a 3d 41 44 47 4f 48 44 3c 46 45 44 45 42 3f 3d 43 3d 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 29 45 3e 49 45 48 4a 45 4d 50 4a 4e 4d 4e 51 52 4c 54 44 4d 42 41 3c 48 3a 3a 40 3d 42 3f 40 41 48 44 41 3f 40 43 37 3b 44 2d 49 43 39 44 39 39 3b 45 3d 40 40 40 3d 40 43 43 3c 41 40 45 52 52 45 4b 4b 41 38 25 13 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 1b 2a 30 34 36 38 32 3c 3d 3f 3d 38 38 3a 42 38 34 3d 38 3e 3b 38 3f 3e 3e 44 3c 3a 3f 3d 45 44 3e 41 45 3e 3e 33 3c 3a 40 40 3a 3b 3d 3c 3e 3c 3e 45 42 3a 38 3f 41 44 3c 40 44 3e 3d 45 48 46 39 44 3e 42 41 39 42 4b 4a 4c 46 3f 43 43 42 3e 44 44 45 3d 3c 3c 3d 3d 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 2a 38 3c 44 45 3b 44 44 4d 50 4e 51 52 54 52 4a 49 3f 3f 44 43 3e 42 43 40 44 36 42 41 46 3b 3f 45 3a 3e 49 3e 3d 43 3c 43 46 37 3b 3d 3c 33 3d 37 3c 41 3d 3b 44 43 3f 45 4b 41 44 45 46 47 4c 3e 49 3a 32 27 14 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0d 1a 2d 29 38 36 44 42 3a 3a 3f 39 3e 3b 37 3b 3f 39 38 47 3c 42 3a 42 3f 3e 38 3e 39 41 44 46 3e 3d 3e 45 41 3e 39 3c 3d 35 3d 41 44 3c 3c 3e 40 45 40 3f 45 3e 3d 40 36 47 46 3e 3c 40 45 3e 42 44 45 46 42 45 3e 45 44 44 3f 49 46 46 40 3d 3e 48 3d 3e 49 49 44 39 26 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 27 41 41 3d 4a 3e 4f 47 44 52 4d 51 51 4d 4b 44 4a 47 41 4a 3e 46 3c 44 39 3c 3b 43 3e 45 48 45 49 42 3d 42 43 3d 3e 36 42 3d 38 3f 3b 44 44 39 43 3d 3e 47 3e 40 3e 39 3b 41 44 3e 3e 45 4f 45 42 3b 2e 20 1a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 13 22 2e 37 43 3d 42 3e 44 45 3b 41 39
 39 3f 3d 37 37 41 38 3b 3b 41 3d 43 41 3b 39 3c 40 3d 3c 43 37 3c 41 3c 45 38 3a 3c 3d 44 48 47 40 42 40 48 3c 3b 37 40 3b 39 3e 44 47 47 39 43 43 43 3e 48 4b 41 45 48 42 40 4e 44 49 4b 4a 42 45 45 3b 41 39 49 42 45 35 41 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1f 48 44 42 48 3e 44 4b 49 4a 4e 4f 47 46 44 43 45 47 41 43 3d 43 3e 3e 43 33 41 48 45 43 40 42 43 3d 47 42 3d 3c 39 3e 3b 46 40 44 40 38 40 40 3c 3d 3d 41 3d 3c 44 38 3b 3d 3d 47 4a 46 41 3d 37 2e 1d 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 15 1e 22 31 3b 36 44 3b 3a 3b 36 35 3c 37 40 36 3e 38 32 3f 44 3e 38 43 36 35 3b 3a 39 39 3d 47 35 3c 41 33 3c 38 3c 36 3a 35 3a 43 47 3a 38 41 3a 36 3d 3b 3c 34 43 3b 3d 44 38 44 42 42 3a 3f 43 44 43 43 4a 44 47 49 4b 4a 47 51 47 49 3e 44 44 42 43 46 3e 3a 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 3d 3e 47 49 44 3c 48 44 46 47 46 43 3e 48 42 3e 44 46 43 40 42 40 3d 37 3f 39 3b 3e 37 43 41 40 41 38 39 42 42 40 3c 3a 3f 40 38 3d 38 42 3b 3b 39 3c 38 31 3a 3d 3f 48 45 3e 46 3d 44 47 3b 25 20 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 16 28 2d 3f 3c 42 48 36 43 3e 41 3d 40 3e 3b 45 38 3e 33 34 4c 43 42 3f 3c 3e 3e 3d 3a 42 3d 42 31 3b 3b 40 38 44 47 43 37 3c 3b 3d 3a 3c 44 32 3b 36 34 35 3e 3a 42 3a 44 3b 44 3c 3d 4a 42 40 49 48 45 43 41 4d 4e 53 4b 43 46 44 43 48 49 40 45 4b 43 45 47 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 40 3f 4c 44 4b 41 47 49 4e 42 4d 3c 43 49 3e 47 3d 42 3d 39 46 44 4a 3a 41 43 39 3f 45 3d 47 39 45 3e 3e 42 44 45 31 3f 3a 40 41 43 3c 3b 45 3e 44 3e 3c 37 43 3e 41 3c 43 3c 3d 3b 43 32 2f 22 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 15 26 35 3a 38 3f 3e 37 3a 3f
 40 3a 41 3b 3b 40 37 40 36 35 3d 3d 36 43 40 3f 3d 3c 42 43 3b 41 3f 41 38 42 39 3b 38 32 40 3b 3e 3e 41 3e 3c 3e 3b 41 47 42 43 3e 41 48 37 41 44 43 3f 47 41 47 49 43 46 45 3d 49 49 49 4d 4f 4c 44 49 3d 42 46 44 47 41 44 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 42 42 4e 41 4a 48 45 46 45 41 46 4c 45 4c 40 45 4a 40 45 41 3f 41 45 37 44 43 3c 43 3f 3f 41 41 48 43 40 3e 39 3d 38 3e 3e 3e 45 39 3c 44 38 40 47 41 36 45 44 44 3e 42 42 3b 3b 3d 32 28 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 1b 22 36 37 3b 38 3b 3e 3b 3b 3c 37 40 3d 35 36 32 39 35 35 31 38 41 40 37 3e 3f 3b 3a 3e 30 3f 43 45 43 40 44 3a 3e 3e 3b 3b 44 41 3b 37 3b 3d 42 42 38 3a 3c 41 41 42 41 3d 3c 3d 45 47 45 48 43 3c 49 38 48 42 45 46 46 46 44 48 43 3c 41 49 3b 40 3e 28 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 36 33 4e 49 3e 3c 41 45 48 3c 3a 3b 44 47 44 3f 46 46 47 45 48 3d 3c 3e 3b 3d 35 41 4a 3d 41 40 44 40 41 38 3f 42 44 42 3d 3d 3b 43 3e 3a 3d 40 44 3a 3b 40 46 47 53 43 44 3b 37 32 23 16 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 15 24 32 3c 34 34 3e 38 3f 41 38 3e 38 3d 35 40 37 3c 3d 42 39 39 3c 39 3b 3c 46 34 3a 3b 2e 3f 3a 3c 3a 39 3c 3f 3f 44 3c 42 3a 3d 3d 43 3b 40 43 39 3e 46 3a 3f 45 3d 41 3b 3b 41 41 44 41 43 45 46 47 4c 3c 4a 3e 46 4b 41 40 44 46 3e 44 43 49 40 34 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 35 49 49 44 3d 39 3d 48 43 42 3c 44 3b 3f 41 3e 41 3f 49 43 4a 46 3f 41 33 3a 3e 46 42 41 46 40 3e 3e 43 4b 46 4a 3b 3b 40 36 39 39 44 37 38 44 3f 40 40 3a 3e 43 3b 40 39 33 2b 1e 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 16 14 26 37 37 36 40 40
 3f 43 3f 3d 39 36 3f 3d 3a 3e 35 3a 38 41 3d 3b 42 3f 3a 3d 44 37 39 3c 39 3b 44 3d 3d 3e 3b 35 3d 3b 3f 42 3c 3f 3c 3a 44 3f 3f 41 37 47 38 40 4a 41 41 4a 4a 43 3f 47 3e 49 42 3f 3e 3f 4b 4a 53 47 4a 42 3f 42 40 41 42 3e 30 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 14 40 4b 4a 47 3d 46 45 48 42 40 42 42 43 42 4a 3e 46 3f 3a 37 3e 40 3c 40 3d 3c 4b 40 41 4c 3d 44 43 3b 46 3d 3e 45 44 3d 43 3d 3e 3a 41 3e 43 45 3a 3c 36 3b 43 40 3b 3a 35 24 1f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 15 26 2a 38 3d 43 37 3f 43 3c 41 3e 37 39 3b 39 37 37 34 41 3a 36 3d 3a 3f 3c 34 3b 38 3a 37 40 37 3c 3f 44 3d 3b 38 41 3c 37 3a 39 3f 3e 44 3c 40 3b 3c 45 39 3d 44 41 3e 47 3a 42 4d 3e 44 46 44 45 3c 48 48 46 4b 44 3f 46 41 3f 45 43 40 3e 2a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3b 40 43 4a 48 47 45 42 2d 40 3f 40 46 3f 47 40 3e 47 4b 3f 4f 43 44 3e 3f 48 46 46 45 44 40 38 3e 43 47 47 3c 3b 3b 42 41 3d 3c 41 3b 3f 3f 40 3c 3b 3f 37 37 37 2f 20 25 0f 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 19 21 2b 36 37 3c 44 3d 37 3d 39 39 36 41 34 36 41 3c 3b 37 3a 3f 3a 3f 40 3a 35 3f 3e 3a 30 36 3b 3a 3b 3a 35 3c 37 38 40 39 3a 39 3c 40 39 3c 3f 3f 44 39 41 3b 3a 3d 3c 42 43 42 43 47 3d 45 4a 41 44 49 40 3f 3f 45 44 3f 4a 44 3f 3e 41 2d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3c 46 4c 45 47 38 3b 39 42 3e 3d 44 42 46 42 3c 47 4b 45 48 44 3b 41 47 3f 40 4b 46 39 41 41 45 3d 41 45 39 43 46 42 3c 3c 3d 40 3f 3e 3d 3a 3b 34 37 35 32 37 2e 25 23 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 14 1d 27 37
 35 3e 3d 35 37 3b 3c 36 3b 3f 42 44 3a 42 39 35 45 3e 40 40 3b 3f 38 34 41 3e 42 3d 3a 39 3c 44 45 42 46 3c 40 3b 3b 42 38 3a 43 3b 43 3d 38 3f 46 45 47 47 43 41 3b 46 3b 46 49 47 3e 46 47 45 41 42 4c 41 40 41 45 48 43 3b 2f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 35 3a 42 4e 43 45 46 4a 4a 43 44 46 49 44 4a 4c 4b 48 49 44 51 48 43 3e 3e 4b 41 44 45 48 44 41 3e 4c 40 45 44 3c 36 3f 43 3c 40 3b 39 42 3a 36 35 31 2d 35 24 17 11 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 04 1a 1a 25 2d 33 36 3c 39 41 3f 40 3d 3e 39 41 3c 41 3d 42 36 38 3a 3f 37 36 47 37 41 3b 3b 36 35 40 3d 3e 43 38 37 42 36 3a 3c 3c 3e 39 43 3d 3f 3f 42 47 42 49 47 40 49 47 4a 3f 44 45 43 4b 44 4c 42 42 45 44 45 3e 45 3b 4d 45 3f 35 33 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 36 3c 43 45 44 4a 4e 46 4d 4e 4a 4c 54 40 4f 54 52 55 4a 56 56 55 56 55 4c 55 4e 4d 4e 4b 4b 48 50 47 38 4c 45 4b 3f 3a 42 45 35 46 38 3d 3e 32 35 2c 2a 1a 17 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 0e 16 23 2d 32 32 3b 3a 35 33 3f 39 43 3d 3c 3b 3e 46 3d 3b 36 3b 41 42 3f 37 39 35 35 3e 3d 39 3d 3c 3d 3e 3f 3d 39 35 3e 40 3b 3f 42 41 47 3f 3e 3e 47 40 3d 3c 3c 40 44 46 47 40 42 42 42 4a 44 4e 45 40 3e 42 41 39 44 45 3b 41 32 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 3b 49 56 50 4c 55 55 4f 5d 5c 62 60 64 62 62 66 63 5f 62 64 6a 6d 6a 5c 65 58 61 5b 54 61 55 59 4b 51 50 4d 4a 4a 4d 4e 48 38 3f 3b 2f 36 2f 2e 26 1a 1b 0f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 12 20 25 2f 2f 3d 38 3f 3a 3c 3d 3f 3b 3c 38 40 3e 3e 3e 3c 3f 41 37 3d 3a 39 3f 3d 38 3e 3c 40 40 3a 41 45 3a 3e 40 39 46 39 45 42 3d 3f 3b 44 4a 45 45 40 40 44 42 48 46 41 46 46 42 51 45 48 3f 3a 46 44 42 46 49 42 49 3e 2a 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 48 52 5a 6b 67 65 68 6c 6c 74 6e 6c 74 73 7e 76 79 78 74 7e 79 7a 7b 75 77 76 77 72 74 73 6f 69 64 62 60 5e 56 5f 57 58 51 4b 48 3d 3a 29 20 1f 16 07 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 1f 21 25 33 3a 39 38 44 39 3a 3d 36 46 3d 3a 42 37 3b 39 43 40 3b 37 3f 3f 3f 39 3d 3b 3a 43 42 39 43 44 40 40 43 3e 3e 42 37 3f 45 43 42 41 41 47 45 3e 46 3e 42 49 4e 40 42 48 4a 3d 44 47 46 41 3c 42 43 40 45 3d 3b 2d 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 4f 62 69 7c 73 76 7e 77 7e 71 7b 7a 7e 82 82 83 77 7c 7e 7f 81 7c 84 83 7e 7f 76 7b 78 7e 75 77 75 76 75 71 65 67 60 59 58 47 3f 3b 2f 1d 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 11 15 22 2b 33 32 3a 35 36 3d 39 44 45 37 3c 39 44 3f 40 3b 30 3c 3e 43 3b 34 3f 3a 3e 3e 3f 3f 3e 3a 43 3f 3a 3f 40 46 42 49 45 3b 41 40 48 41 3e 40 3d 3f 45 42 37 40 46 4a 3e 4a 4d 41 44 45 42 45 3f 43 3d 42 41 38 31 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 4f 6e 7e 7e 79 6d 77 7d 7a 7a 79 7d 7a 77 80 7e 81 7e 7d 82 84 7e 81 80 80 7b 84 7f 7e 7e 7b 80 7c 7a 6e 68 68 67 63 5f 56 45 3d 25 1b 16 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 02 06 09 16 20 22 28 36 3f 3f 3f 40 43 3e 3e 3b 3e 43 3c 3b 3d 3c 3d 45 3d 3d 3a 33 41 3e 41 45 3d 42 43 44 42 40 4c 3a 3f 43 42 3f 3e 3d 40 47 46 4b 41 47 46 42 49 40 40 49 44 45 4a 47 4a 45 49 45 3d 45 3c 43 44 41 40 37 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 56 72 7e 82 7b 78 76 80 77 7b 79 77 7d 7f 80 7c 78 7d 7c 76 81 7f 7d 7b 7f 7a 80 7d 7e 80 74 77 6b 6c 6e 69 65 5f 53 51 38 33 1d 11 06 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0d 19 25 24 31 35 3a 39 3c 3b 3c 36 43 38 3e 3a 3e 40 41 40 3a 43 3c 41 41 41 42 41 3e 46 49 38 45 42 3d 3d 47 48 48 40 4c 3f 46 42 41 4b 47 40 4b 40 45 49 44 47 45 49 42 42 4f 40 4a 49 4a 43 49 4b 43 3a 41 38 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 46 6c 71 7e 6f 73 77 71 77 75 7a 7a 7c 7b 7b 78 7d 7c 76 73 74 77 7d 79 76 73 73 76 7f 74 6e 6a 69 6a 64 60 54 47 44 31 24 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 11 1d 2b 26 35 39 3a 44 37 36 3f 3f 44 3f 48 41 3c 49 45 45 3f 40 41 3a 45 40 4b 3f 44 4b 3e 40 45 40 43 48 47 4b 49 48 4a 48 46 49 45 4a 44 48 46 46 43 4e 4c 47 4e 48 49 4b 49 4f 4b 4d 4a 49 4b 47 4f 3f 24 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 45 68 72 72 6f 74 74 70 70 6f 72 71 71 76 71 73 75 71 75 70 72 73 70 72 68 6e 70 67 6f 6a 62 5c 56 55 4d 43 3e 35 24 18 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 01 06 0d 14 24 25 33 3a 3e 3e 44 40 3f 42 49 42 46 3f 44 47 4d 45 42 41 48 44 49 40 42 4a 4f 45 49 4d 49 53 49 4f 4d 48 53 4f 53 57 4d 55 50 4b 50 51 55 51 4b 55 58 5f 54 53 54 52 5a 53 56 52 5c 57 64 5d 53 4a 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3f 5c 6c 75 6d 66 6b 67 6b 69 70 71 76 6d 73 6c 6b 73 71 66 6c 63 6e 66 69 68 63 66 64 5e 5a 53 47 40 3e 2b 1f 1d 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 1b 25 36 3d 3b 4b 43 45 4a 47 47 4a 4f 4b 55 4f 51 47 4a 50 4a 51 55 57 55 4f 53 56 56 4f 55 53 56 5a 5c 5d 57 57 5f 60 59 5f 67 5d 62 5c 63 61 61 68 69 6f 65 64 68 67 64 66 6a 69 71 6a 68 5f 5e 28 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 38 5a 60 66 65 65 60 71 6b 5e 66 70 67 6b 6e 6a 6f 6f 66 65 68 63 60 64 58 5d 63 51 4d 49 4a 35 36 2b 1f 1a 15 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 16 21 34 37 40 3c 4a 49 4f 52 4f 55 56 57 5f 51 57 57 53 56 5b 5c 5d 5b 5f 65 64 5e 68 64 5f 5e 6a 65 6c 71 72 6c 69 67 6d 70 78 6e 6d 78 6d 6d 6d 75 76 75 74 71 6d 6c 6e 70 65 72 6e 68 6a 5b 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 32 52 5e 61 5d 5e 61 65 64 5f 5b 62 65 64 65 5a 64 62 60 5a 5b 5b 5b 4e 49 45 4d 43 3f 33 2f 1d 21 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 07 12 21 31 3b 42 4b 5b 54 5f 5f 5c 60 68 65 60 5f 5f 69 6f 6c 6b 69 6b 70 76 79 6f 6c 72 71 74 7b 77 76 6c 77 7c 79 7f 84 75 7d 76 78 7c 7b 73 72 75 76 79 79 74 70 6f 79 67 68 75 65 64 5e 55 2e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2f 56 5e 65 5d 5b 54 5a 54 5e 5f 5d 58 5e 56 4e 52 5b 5b 4d 4a 42 4d 42 39 36 36 2f 26 20 16 14 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 15 17 24 3c 3f 4a 59 59 63 61 6b 6d 6a 6c 6b 75 76 75 74 72 7b 77 7e 76 80 7c 7a 84 7b 81 7b 79 81 81 7b 81 78 79 7b 78 77 7d 77 76 7a 7d 7e 7a 79 76 6b 73 6c 6e 6c 6c 65 73 73 62 65 5f 2e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 4c 52 5f 5d 4f 5e 54 58 57 52 53 54 50 50 4f 48 45 42 45 41 33 2d 2a 2a 21 1d 17 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0f 22 21 3b 40 4b 51 59 64 62 6d 78 72 77 71 72 74 77 74 79 7b 74 68 7f 76 7d 7b 76 7c 7c 7d 77 7b 74 75 74 75 7b 73 77 77 6a 73 6e 6c 71 71 6f 64 65 6c 69 71 67 6a 5f 6b 69 59 60 5a 2b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 3b 5d 5c 4a 4c 4b 4b 53 55 4c 48 46 43 40 39 3c 3b 2e 29 2b 1d 1d 1c 0c 12 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 20 2a 3b 4e 56 5e 5d 60 66 6e 72 71 74 70 75 71 78 7a 7a 73 6e 70 75 75 7f 72 6b 71 6b 73 70 6d 69 6f 68 6e 6f 6d 64 67 6d 70 74 68 64 68 65 64 65 63 60 5b 62 62 59 5b 50 4b 30 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 3f 45 40 46 3c 3b 41 37 38 40 31 2e 32 29 2b 29 1e 19 0d 11 03 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 0e 18 2a 2f 42 49 51 5d 62 69 67 62 69 6c 75 71 70 72 72 71 6e 72 6d 71 65 70 6d 69 6d 6d 64 65 62 64 64 64 66 63 57 61 62 6c 68 61 66 5e 61 60 60 5e 5c 60 63 61 54 56 50 52 2f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 30 3b 36 31 31 2f 2c 29 25 1e 24 1c 1b 0a 13 0b 08 09 09 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0f 18 1b 2a 28 3b 4e 4f 5a 55 5d 5c 62 66 6c 6d 70 6a 62 69 66 6c 6e 67 62 69 65 5e 60 61 62 63 60 60 60 5f 65 60 5d 5b 64 5f 5a 67 5c 5a 62 58 54 5a 4e 5a 54 59 50 5a 50 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1b 24 25 17 1a 1e 12 14 0f 0d 06 09 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 0f 1b 22 20 32 36 3f 4c 54 4b 50 64 5e 60 62 67 63 64 5e 5f 62 60 5a 5c 5e 61 52 58 51 56 54 52 57 5d 5b 59 5c 5a 55 5b 5b 60 57 5f 52 51 54 53 57 53 49 52 47 4b 47 30 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 0d 05 0a 0b 06 09 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 12 15 1c 24 2b 38 47 4a 50 46 4d 50 5b 59 53 52 5c 5f 5a 59 59 53 4a 51 4a 4e 4c 4a 4b 4e 52 56 56 52 5b 4f 5a 57 50 56 52 57 4e 51 4b 4f 51 48 4c 47 44 3f 3e 31 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 10 12 24 29 26 35 3f 49 40 45 4a 4e 51 4f 49 4b 47 4b 47 44 3c 2d 32 3e 3f 3b 46 46 51 4d 4e 53 54 43 50 49 4c 4e 44 45 43 4a 45 3b 44 35 3b 38 35 37 24 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0b 19 10 18 25 31 28 30 39 31 35 38 38 41 3d 3a 38 2b 22 12 1e 1e 23 2f 35 3d 43 47 41 44 39 3f 40 32 3d 3d 3c 37 31 30 33 2c 27 2b 26 24 1c 1d 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0b 16 15 12 21 1c 2d 26 21 28 2c 29 27 27 16 11 06 11 13 15 19 26 30 29 30 33 29 31 2a 2b 25 27 2b 25 1c 1b 17 14 16 12 10 13 0d 03 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0c 0e 12 0f 14 11 13 14 12 10 0f 03 06 05 08 02 0b 05 0f 14 19 17 11 10 13 0b 03 0e 06 05 0d 06 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
