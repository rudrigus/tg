 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 07 07 07 05 05 05 06 06 06 07 07 07 07 07 07 05 05 05 04 04 04 04 04 04 06 06 06 0c 0c 0c 0c 0c 0c 09 09 09 0a 0a 0a 06 06 06 07 07 07 05 05 05 04 04 04 04 04 04 03 03 03 05 05 05 03 03 03 04 04 04 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 08 08 08 0d 0d 0d 14 14 14 1e 1e 1e 2d 2d 2d 38 38 38 51 51 51 36 36 36 29 29 29 1c 1c 1c 2d 2d 2d 56 56 56 5c 5c 5c 57 57 57 3f 3f 3f 3c 3c 3c 3b 3b 3b 32 32 32 35 35 35 36 36 36 23 23 23 1b 1b 1b 15 15 15 0e 0e 0e 09 09 09 06 06 06 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 04 04 04 07 07 07 0c 0c 0c 1d 1d 1d 37 37 37 63 63 63 89 89 89 89 89 89 ac ac ac bf bf bf a8 a8 a8 73 73 73 5d 5d 5d 5f 5f 5f 61 61 61 64 64 64 61 61 61 5b 5b 5b 50 50 50 48 48 48 4b 4b 4b 4f 4f 4f 52 52 52 56 56 56 79 79 79 9e 9e 9e 95 95 95 6f 6f 6f 51 51 51 49 49 49 38 38 38 1c 1c 1c 0e 0e 0e 06 06 06 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 0b 0b 0b 17 17 17 37 37 37 5c 5c 5c 6b 6b 6b 8b 8b 8b 93 93 93 bc bc bc c4 c4 c4 b5 b5 b5 9c 9c 9c 89 89 89 70 70 70 64 64 64 6d 6d 6d 74 74 74 73 73 73 68 68 68 65 65 65 5a 5a 5a 53 53 53 56 56 56 60 60 60 61 61 61 62 62 62 6f 6f 6f 75 75 75 74 74 74 6b 6b 6b 67 67 67 6a 6a 6a 7a 7a 7a 6c 6c 6c 5d 5d 5d 32 32 32 12 12 12 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 0f 0f 0f 21 21 21 4c 4c 4c 74 74 74 77 77 77 80 80 80 80 80 80 8d 8d 8d 95 95 95 ae ae ae bb bb bb b3 b3 b3 a2 a2 a2 9a 9a 9a 89 89 89 82 82 82 87 87 87 8e 8e 8e 8a 8a 8a 84 84 84 80 80 80 79 79 79 6d 6d 6d 67 67 67 6b 6b 6b 6c 6c 6c 68 68 68 73 73 73 7a 7a 7a 79 79 79 7b 7b 7b 7c 7c 7c 77 77 77 78 78 78 72 72 72 92 92 92 a1 a1 a1 6c 6c 6c 2d 2d 2d 0f 0f 0f 05 05 05 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 0b 0b 0b 1f 1f 1f 4f 4f 4f 99 99 99 a5 a5 a5 82 82 82 87 87 87 90 90 90 8f 8f 8f a0 a0 a0 a2 a2 a2 bb bb bb d4 d4 d4 c4 c4 c4 a7 a7 a7 a4 a4 a4 a0 a0 a0 a6 a6 a6 ae ae ae b2 b2 b2 ae ae ae a7 a7 a7 9d 9d 9d 96 96 96 8c 8c 8c 7c 7c 7c 77 77 77 73 73 73 6d 6d 6d 7b 7b 7b 8b 8b 8b 95 95 95 9a 9a 9a 98 98 98 91 91 91 8a 8a 8a 7d 7d 7d 7c 7c 7c 83 83 83 8d 8d 8d 6d 6d 6d 32 32 32 0a 0a 0a 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 06 06 06 13 13 13 33 33 33 74 74 74 98 98 98 9d 9d 9d 8c 8c 8c 90 90 90 99 99 99 ac ac ac ad ad ad bd bd bd cb cb cb d8 d8 d8 e4 e4 e4 d0 d0 d0 b0 b0 b0 a8 a8 a8 a7 a7 a7 b5 b5 b5 c2 c2 c2 c5 c5 c5 c2 c2 c2 b9 b9 b9 b3 b3 b3 ac ac ac a2 a2 a2 94 94 94 87 87 87 7f 7f 7f 77 77 77 87 87 87 a2 a2 a2 b3 b3 b3 b6 b6 b6 b3 b3 b3 a6 a6 a6 9b 9b 9b 92 92 92 89 89 89 8a 8a 8a 8d 8d 8d 85 85 85 79 79 79 30 30 30 07 07 07 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 08 08 08 1b 1b 1b 4a 4a 4a 83 83 83 7a 7a 7a 75 75 75 86 86 86 89 89 89 98 98 98 a7 a7 a7 ba ba ba c6 c6 c6 cf cf cf e4 e4 e4 ef ef ef ea ea ea d4 d4 d4 ba ba ba b1 b1 b1 a9 a9 a9 b7 b7 b7 c4 c4 c4 c8 c8 c8 c6 c6 c6 c0 c0 c0 bd bd bd b7 b7 b7 ac ac ac a5 a5 a5 9e 9e 9e 90 90 90 86 86 86 96 96 96 b5 b5 b5 c7 c7 c7 c7 c7 c7 c1 c1 c1 b6 b6 b6 b3 b3 b3 a5 a5 a5 9b 9b 9b 91 91 91 8b 8b 8b 8f 8f 8f 93 93 93 68 68 68 1d 1d 1d 05 05 05 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 28 28 28 5f 5f 5f 6b 6b 6b 6b 6b 6b 70 70 70 7a 7a 7a 88 88 88 94 94 94 9c 9c 9c ab ab ab b8 b8 b8 cf cf cf dd dd dd eb eb eb f7 f7 f7 ef ef ef d6 d6 d6 c5 c5 c5 c1 c1 c1 b3 b3 b3 ba ba ba c5 c5 c5 cc cc cc cd cd cd cc cc cc c5 c5 c5 be be be bb bb bb b7 b7 b7 b3 b3 b3 aa aa aa a0 a0 a0 aa aa aa c6 c6 c6 d6 d6 d6 d2 d2 d2 d0 d0 d0 c9 c9 c9 c3 c3 c3 b4 b4 b4 a3 a3 a3 95 95 95 8c 8c 8c 89 89 89 89 89 89 a6 a6 a6 52 52 52 15 15 15 04 04 04 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 20 20 20 73 73 73 86 86 86 77 77 77 7a 7a 7a 84 84 84 8b 8b 8b 94 94 94 a1 a1 a1 ad ad ad b8 b8 b8 c5 c5 c5 d0 d0 d0 de de de ec ec ec f3 f3 f3 ee ee ee d8 d8 d8 cd cd cd d1 d1 d1 c9 c9 c9 cf cf cf ee ee ee f6 f6 f6 f6 f6 f6 ef ef ef de de de d1 d1 d1 cd cd cd ce ce ce cd cd cd ca ca ca bf bf bf c1 c1 c1 d2 d2 d2 df df df de de de df df df d4 d4 d4 c7 c7 c7 b2 b2 b2 a1 a1 a1 94 94 94 8f 8f 8f 89 89 89 79 79 79 a5 a5 a5 94 94 94 3b 3b 3b 06 06 06 03 03 03 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 04 04 04 10 10 10 44 44 44 8c 8c 8c 88 88 88 83 83 83 86 86 86 8a 8a 8a 95 95 95 9d 9d 9d a9 a9 a9 b8 b8 b8 be be be c6 c6 c6 d0 d0 d0 da da da e4 e4 e4 ed ed ed e6 e6 e6 d8 d8 d8 d2 d2 d2 db db db e1 e1 e1 f8 f8 f8 ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb e9 e9 e9 e5 e5 e5 ec ec ec ec ec ec e1 e1 e1 cf cf cf ca ca ca d6 d6 d6 e0 e0 e0 e1 e1 e1 e2 e2 e2 d6 d6 d6 c3 c3 c3 a8 a8 a8 99 99 99 96 96 96 8f 8f 8f 7e 7e 7e 77 77 77 7b 7b 7b 9d 9d 9d 58 58 58 10 10 10 04 04 04 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0e 0e 0e 33 33 33 5a 5a 5a 6c 6c 6c 81 81 81 83 83 83 89 89 89 90 90 90 97 97 97 a3 a3 a3 b1 b1 b1 bc bc bc c5 c5 c5 ce ce ce d5 d5 d5 df df df e5 e5 e5 e6 e6 e6 e0 e0 e0 d2 d2 d2 d2 d2 d2 de de de ee ee ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc fd fd fd fb fb fb e7 e7 e7 d6 d6 d6 cf cf cf cf cf cf d9 d9 d9 e3 e3 e3 e4 e4 e4 e2 e2 e2 cf cf cf b7 b7 b7 a4 a4 a4 98 98 98 90 90 90 84 84 84 7e 7e 7e 78 78 78 73 73 73 76 76 76 7d 7d 7d 30 30 30 08 08 08 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 09 09 09 2d 2d 2d 51 51 51 60 60 60 6a 6a 6a 78 78 78 7d 7d 7d 87 87 87 92 92 92 96 96 96 a3 a3 a3 b3 b3 b3 c2 c2 c2 cc cc cc d6 d6 d6 df df df ea ea ea ee ee ee ee ee ee df df df d2 d2 d2 d3 d3 d3 e4 e4 e4 f0 f0 f0 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc f2 f2 f2 e1 e1 e1 d3 d3 d3 cf cf cf d2 d2 d2 d6 d6 d6 dc dc dc e0 e0 e0 e2 e2 e2 da da da c1 c1 c1 ae ae ae 9e 9e 9e 96 96 96 8f 8f 8f 88 88 88 7d 7d 7d 75 75 75 72 72 72 6e 6e 6e 7b 7b 7b 50 50 50 08 08 08 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0f 0f 0f 48 48 48 71 71 71 66 66 66 6b 6b 6b 72 72 72 7b 7b 7b 81 81 81 8d 8d 8d 9a 9a 9a a1 a1 a1 b0 b0 b0 c2 c2 c2 d0 d0 d0 dd dd dd e7 e7 e7 f2 f2 f2 f6 f6 f6 f5 f5 f5 eb eb eb dd dd dd e0 e0 e0 f6 f6 f6 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fb e3 e3 e3 dc dc dc d7 d7 d7 d5 d5 d5 d7 d7 d7 da da da df df df e2 e2 e2 de de de d0 d0 d0 b9 b9 b9 ab ab ab a0 a0 a0 9a 9a 9a 8f 8f 8f 83 83 83 79 79 79 73 73 73 69 69 69 67 67 67 69 69 69 5c 5c 5c 0b 0b 0b 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0d 0d 0d 52 52 52 6d 6d 6d 67 67 67 69 69 69 6f 6f 6f 7d 7d 7d 86 86 86 88 88 88 96 96 96 a2 a2 a2 af af af bd bd bd cc cc cc da da da e5 e5 e5 f0 f0 f0 f5 f5 f5 f6 f6 f6 ec ec ec e3 e3 e3 e6 e6 e6 f9 f9 f9 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f9 f9 f6 f6 f6 f8 f8 f8 ef ef ef ea ea ea e7 e7 e7 e8 e8 e8 e6 e6 e6 e2 e2 e2 d9 d9 d9 c8 c8 c8 bb bb bb ab ab ab 9d 9d 9d 92 92 92 87 87 87 7f 7f 7f 77 77 77 70 70 70 64 64 64 5e 5e 5e 68 68 68 63 63 63 0f 0f 0f 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 10 10 10 4e 4e 4e 75 75 75 65 65 65 67 67 67 71 71 71 7d 7d 7d 85 85 85 87 87 87 92 92 92 a1 a1 a1 ab ab ab b7 b7 b7 c3 c3 c3 cd cd cd d6 d6 d6 e2 e2 e2 e8 e8 e8 e8 e8 e8 e5 e5 e5 df df df de de de e5 e5 e5 f8 f8 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc fa fa fa f9 f9 f9 f0 f0 f0 e9 e9 e9 e4 e4 e4 e2 e2 e2 dc dc dc d4 d4 d4 cd cd cd be be be b3 b3 b3 a8 a8 a8 95 95 95 8c 8c 8c 84 84 84 7a 7a 7a 75 75 75 6a 6a 6a 63 63 63 5a 5a 5a 66 66 66 63 63 63 0e 0e 0e 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 18 18 18 59 59 59 89 89 89 67 67 67 68 68 68 74 74 74 7e 7e 7e 7e 7e 7e 82 82 82 8d 8d 8d 97 97 97 9b 9b 9b a6 a6 a6 b0 b0 b0 bc bc bc c5 c5 c5 ce ce ce d6 d6 d6 dd dd dd e2 e2 e2 d9 d9 d9 d1 d1 d1 d4 d4 d4 f6 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc e4 e4 e4 e2 e2 e2 dd dd dd d8 d8 d8 d1 d1 d1 cb cb cb c5 c5 c5 bf bf bf b8 b8 b8 b2 b2 b2 a9 a9 a9 9f 9f 9f 8e 8e 8e 85 85 85 7e 7e 7e 79 79 79 70 70 70 6d 6d 6d 63 63 63 59 59 59 63 63 63 62 62 62 0d 0d 0d 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 17 17 17 64 64 64 96 96 96 66 66 66 67 67 67 6a 6a 6a 74 74 74 7c 7c 7c 86 86 86 8f 8f 8f 97 97 97 92 92 92 94 94 94 a0 a0 a0 ab ab ab b2 b2 b2 bb bb bb c4 c4 c4 c1 c1 c1 c3 c3 c3 bd bd bd bd bd bd c2 c2 c2 f7 f7 f7 ff ff ff ff ff ff f9 f9 f9 f6 f6 f6 fe fe fe ff ff ff fe fe fe d8 d8 d8 ce ce ce c9 c9 c9 c4 c4 c4 bd bd bd b4 b4 b4 ad ad ad a6 a6 a6 a0 a0 a0 9a 9a 9a 92 92 92 8e 8e 8e 84 84 84 80 80 80 7e 7e 7e 75 75 75 71 71 71 6b 6b 6b 61 61 61 5a 5a 5a 64 64 64 62 62 62 1a 1a 1a 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 10 10 10 5f 5f 5f 99 99 99 65 65 65 65 65 65 67 67 67 6c 6c 6c 6e 6e 6e 7e 7e 7e 84 84 84 83 83 83 8d 8d 8d 92 92 92 96 96 96 9c 9c 9c a2 a2 a2 ac ac ac b1 b1 b1 ae ae ae b1 b1 b1 ab ab ab aa aa aa b3 b3 b3 f7 f7 f7 fc fc fc df df df b0 b0 b0 b6 b6 b6 ca ca ca e5 e5 e5 fe fe fe e3 e3 e3 d1 d1 d1 c3 c3 c3 b3 b3 b3 a8 a8 a8 a0 a0 a0 96 96 96 8e 8e 8e 88 88 88 7e 7e 7e 7b 7b 7b 7d 7d 7d 7a 7a 7a 78 78 78 7a 7a 7a 73 73 73 6e 6e 6e 67 67 67 60 60 60 5a 5a 5a 5f 5f 5f 66 66 66 2a 2a 2a 04 04 04 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 16 16 16 4b 4b 4b 8e 8e 8e 61 61 61 63 63 63 68 68 68 66 66 66 67 67 67 76 76 76 7e 7e 7e 7b 7b 7b 84 84 84 8c 8c 8c 86 86 86 8b 8b 8b 98 98 98 b2 b2 b2 a2 a2 a2 a5 a5 a5 a8 a8 a8 a0 a0 a0 9e 9e 9e a5 a5 a5 e9 e9 e9 a9 a9 a9 7e 7e 7e 82 82 82 97 97 97 ba ba ba d7 d7 d7 fd fd fd fd fd fd ee ee ee c8 c8 c8 b1 b1 b1 a2 a2 a2 96 96 96 88 88 88 80 80 80 7b 7b 7b 71 71 71 6a 6a 6a 6c 6c 6c 6f 6f 6f 70 70 70 7a 7a 7a 75 75 75 6a 6a 6a 62 62 62 5d 5d 5d 59 59 59 57 57 57 6e 6e 6e 30 30 30 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 05 05 05 21 21 21 3d 3d 3d 66 66 66 5d 5d 5d 5b 5b 5b 5f 5f 5f 64 64 64 64 64 64 6e 6e 6e 71 71 71 72 72 72 76 76 76 7d 7d 7d 77 77 77 77 77 77 86 86 86 9b 9b 9b 9a 9a 9a 9b 9b 9b 9c 9c 9c 95 95 95 91 91 91 9a 9a 9a e3 e3 e3 6c 6c 6c 64 64 64 89 89 89 c8 c8 c8 f3 f3 f3 fd fd fd ff ff ff ff ff ff fe fe fe d5 d5 d5 a9 a9 a9 9d 9d 9d 91 91 91 82 82 82 7a 7a 7a 74 74 74 6c 6c 6c 69 69 69 68 68 68 6b 6b 6b 78 78 78 7f 7f 7f 78 78 78 6d 6d 6d 63 63 63 59 59 59 57 57 57 57 57 57 73 73 73 30 30 30 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 27 27 27 48 48 48 58 58 58 58 58 58 59 59 59 5b 5b 5b 5e 5e 5e 60 60 60 67 67 67 6a 6a 6a 6c 6c 6c 6c 6c 6c 72 72 72 6d 6d 6d 6f 6f 6f 79 79 79 85 85 85 91 91 91 96 96 96 97 97 97 8e 8e 8e 89 89 89 8c 8c 8c ca ca ca 55 55 55 65 65 65 b8 b8 b8 fb fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e0 e0 e0 a5 a5 a5 97 97 97 8a 8a 8a 7a 7a 7a 73 73 73 70 70 70 6c 6c 6c 69 69 69 68 68 68 6b 6b 6b 78 78 78 77 77 77 71 71 71 6c 6c 6c 5e 5e 5e 53 53 53 51 51 51 56 56 56 72 72 72 20 20 20 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 23 23 23 6c 6c 6c 6c 6c 6c 59 59 59 5a 5a 5a 5a 5a 5a 59 59 59 5e 5e 5e 64 64 64 62 62 62 65 65 65 65 65 65 69 69 69 67 67 67 6b 6b 6b 6c 6c 6c 7a 7a 7a 89 89 89 94 94 94 8f 8f 8f 88 88 88 83 83 83 84 84 84 8f 8f 8f 4f 4f 4f 73 73 73 dc dc dc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dd dd dd a7 a7 a7 93 93 93 83 83 83 72 72 72 6d 6d 6d 6d 6d 6d 69 69 69 65 65 65 64 64 64 69 69 69 6f 6f 6f 69 69 69 64 64 64 61 61 61 5a 5a 5a 51 51 51 52 52 52 58 58 58 65 65 65 0d 0d 0d 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 04 04 04 16 16 16 6a 6a 6a 7b 7b 7b 63 63 63 61 61 61 67 67 67 5d 5d 5d 5e 5e 5e 63 63 63 5f 5f 5f 5d 5d 5d 5d 5d 5d 64 64 64 60 60 60 64 64 64 65 65 65 71 71 71 81 81 81 90 90 90 88 88 88 83 83 83 7c 7c 7c 76 76 76 70 70 70 4c 4c 4c 71 71 71 d7 d7 d7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe cb cb cb a1 a1 a1 8e 8e 8e 76 76 76 68 68 68 63 63 63 64 64 64 62 62 62 5e 5e 5e 60 60 60 65 65 65 64 64 64 5f 5f 5f 5c 5c 5c 5c 5c 5c 58 58 58 55 55 55 55 55 55 5d 5d 5d 3a 3a 3a 04 04 04 03 03 03 03 03 03
 03 03 03 02 02 02 04 04 04 04 04 04 10 10 10 47 47 47 74 74 74 57 57 57 57 57 57 57 57 57 59 59 59 5f 5f 5f 6e 6e 6e 5f 5f 5f 5b 5b 5b 5c 5c 5c 5f 5f 5f 63 63 63 62 62 62 62 62 62 69 69 69 73 73 73 80 80 80 81 81 81 7e 7e 7e 73 73 73 64 64 64 5b 5b 5b 48 48 48 5f 5f 5f aa aa aa f9 f9 f9 ff ff ff ff ff ff ff ff ff ff ff ff f8 f8 f8 b0 b0 b0 99 99 99 87 87 87 6d 6d 6d 61 61 61 62 62 62 63 63 63 5f 5f 5f 5e 5e 5e 60 60 60 5b 5b 5b 59 59 59 5a 5a 5a 58 58 58 58 58 58 59 59 59 59 59 59 53 53 53 51 51 51 17 17 17 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 04 04 04 11 11 11 27 27 27 65 65 65 5c 5c 5c 55 55 55 54 54 54 58 58 58 59 59 59 63 63 63 69 69 69 67 67 67 63 63 63 6a 6a 6a 6a 6a 6a 67 67 67 67 67 67 67 67 67 6f 6f 6f 7b 7b 7b 79 79 79 79 79 79 6d 6d 6d 5a 5a 5a 4c 4c 4c 3b 3b 3b 4f 4f 4f 7e 7e 7e c9 c9 c9 fc fc fc ff ff ff ff ff ff ff ff ff e6 e6 e6 9a 9a 9a 8e 8e 8e 79 79 79 65 65 65 5d 5d 5d 64 64 64 63 63 63 60 60 60 57 57 57 56 56 56 53 53 53 57 57 57 59 59 59 58 58 58 56 56 56 56 56 56 54 54 54 54 54 54 37 37 37 05 05 05 02 02 02 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 0d 0d 0d 20 20 20 4b 4b 4b 6a 6a 6a 51 51 51 54 54 54 59 59 59 5a 5a 5a 5c 5c 5c 65 65 65 64 64 64 5d 5d 5d 5f 5f 5f 62 62 62 63 63 63 64 64 64 6f 6f 6f 78 78 78 79 79 79 74 74 74 73 73 73 67 67 67 56 56 56 45 45 45 2b 2b 2b 39 39 39 66 66 66 8a 8a 8a c6 c6 c6 f8 f8 f8 fd fd fd f7 f7 f7 b9 b9 b9 86 86 86 7c 7c 7c 6a 6a 6a 5b 5b 5b 5b 5b 5b 60 60 60 5a 5a 5a 53 53 53 52 52 52 55 55 55 57 57 57 5a 5a 5a 5d 5d 5d 54 54 54 53 53 53 51 51 51 50 50 50 46 46 46 12 12 12 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 0a 0a 0a 23 23 23 3c 3c 3c 6a 6a 6a 52 52 52 52 52 52 55 55 55 55 55 55 56 56 56 57 57 57 56 56 56 59 59 59 5f 5f 5f 60 60 60 61 61 61 61 61 61 66 66 66 6c 6c 6c 6f 6f 6f 72 72 72 71 71 71 67 67 67 57 57 57 42 42 42 22 22 22 1c 1c 1c 44 44 44 69 69 69 83 83 83 ab ab ab c4 c4 c4 ba ba ba 8f 8f 8f 7b 7b 7b 72 72 72 66 66 66 5a 5a 5a 5e 5e 5e 5f 5f 5f 5b 5b 5b 58 58 58 59 59 59 58 58 58 57 57 57 53 53 53 5a 5a 5a 55 55 55 50 50 50 4e 4e 4e 4b 4b 4b 2f 2f 2f 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 04 04 04 04 04 04 06 06 06 1e 1e 1e 34 34 34 4e 4e 4e 51 51 51 50 50 50 4f 4f 4f 54 54 54 51 51 51 50 50 50 52 52 52 55 55 55 5b 5b 5b 5e 5e 5e 5c 5c 5c 59 59 59 5e 5e 5e 61 61 61 69 69 69 6e 6e 6e 70 70 70 6b 6b 6b 60 60 60 45 45 45 22 22 22 0a 0a 0a 1d 1d 1d 3f 3f 3f 53 53 53 62 62 62 70 70 70 80 80 80 74 74 74 6d 6d 6d 68 68 68 64 64 64 60 60 60 66 66 66 64 64 64 5d 5d 5d 58 58 58 57 57 57 58 58 58 4b 4b 4b 4c 4c 4c 56 56 56 55 55 55 4d 4d 4d 4e 4e 4e 48 48 48 17 17 17 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 0b 0b 0b 26 26 26 3c 3c 3c 42 42 42 3e 3e 3e 40 40 40 45 45 45 43 43 43 42 42 42 41 41 41 44 44 44 49 49 49 4d 4d 4d 4c 4c 4c 48 48 48 4c 4c 4c 50 50 50 56 56 56 5a 5a 5a 5b 5b 5b 59 59 59 52 52 52 36 36 36 1b 1b 1b 04 04 04 05 05 05 0e 0e 0e 20 20 20 2f 2f 2f 37 37 37 57 57 57 57 57 57 59 59 59 58 58 58 4d 4d 4d 47 47 47 4c 4c 4c 4c 4c 4c 49 49 49 4b 4b 4b 4a 4a 4a 4c 4c 4c 49 49 49 49 49 49 4b 4b 4b 4c 4c 4c 46 46 46 46 46 46 3e 3e 3e 09 09 09 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 19 19 19 35 35 35 3b 3b 3b 3c 3c 3c 3d 3d 3d 3c 3c 3c 3b 3b 3b 3b 3b 3b 3c 3c 3c 3e 3e 3e 44 44 44 47 47 47 48 48 48 47 47 47 48 48 48 4a 4a 4a 4d 4d 4d 52 52 52 54 54 54 54 54 54 55 55 55 3c 3c 3c 20 20 20 03 03 03 03 03 03 03 03 03 05 05 05 0e 0e 0e 1a 1a 1a 43 43 43 4a 4a 4a 4f 4f 4f 4c 4c 4c 47 47 47 46 46 46 46 46 46 48 48 48 47 47 47 45 45 45 42 42 42 48 48 48 47 47 47 44 44 44 44 44 44 44 44 44 43 43 43 45 45 45 28 28 28 04 04 04 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 2a 2a 2a 39 39 39 39 39 39 37 37 37 36 36 36 3b 3b 3b 39 39 39 38 38 38 3a 3a 3a 3d 3d 3d 42 42 42 4e 4e 4e 48 48 48 46 46 46 47 47 47 49 49 49 4c 4c 4c 52 52 52 55 55 55 5a 5a 5a 47 47 47 24 24 24 03 03 03 03 03 03 02 02 02 03 03 03 04 04 04 08 08 08 38 38 38 42 42 42 48 48 48 45 45 45 47 47 47 49 49 49 46 46 46 46 46 46 44 44 44 43 43 43 42 42 42 45 45 45 43 43 43 42 42 42 43 43 43 44 44 44 41 41 41 40 40 40 0f 0f 0f 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 37 37 37 37 37 37 34 34 34 34 34 34 37 37 37 38 38 38 37 37 37 38 38 38 3a 3a 3a 3e 3e 3e 42 42 42 47 47 47 4c 4c 4c 48 48 48 47 47 47 48 48 48 4e 4e 4e 55 55 55 58 58 58 4e 4e 4e 2f 2f 2f 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 34 34 34 3f 3f 3f 45 45 45 47 47 47 48 48 48 48 48 48 47 47 47 43 43 43 43 43 43 43 43 43 44 44 44 43 43 43 41 41 41 45 45 45 46 46 46 45 45 45 46 46 46 2b 2b 2b 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 22 22 22 37 37 37 36 36 36 35 35 35 3a 3a 3a 39 39 39 39 39 39 39 39 39 3c 3c 3c 3d 3d 3d 42 42 42 44 44 44 4b 4b 4b 51 51 51 4c 4c 4c 48 48 48 4f 4f 4f 54 54 54 56 56 56 51 51 51 33 33 33 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 04 04 04 37 37 37 44 44 44 4a 4a 4a 46 46 46 46 46 46 47 47 47 49 49 49 45 45 45 44 44 44 44 44 44 42 42 42 44 44 44 43 43 43 45 45 45 47 47 47 49 49 49 40 40 40 11 11 11 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 2f 2f 2f 37 37 37 35 35 35 3a 3a 3a 39 39 39 39 39 39 3b 3b 3b 3d 3d 3d 3f 3f 3f 3f 3f 3f 42 42 42 47 47 47 4a 4a 4a 4c 4c 4c 49 49 49 4c 4c 4c 50 50 50 51 51 51 4f 4f 4f 37 37 37 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 3e 3e 3e 45 45 45 42 42 42 46 46 46 46 46 46 46 46 46 44 44 44 42 42 42 44 44 44 42 42 42 41 41 41 42 42 42 43 43 43 44 44 44 48 48 48 49 49 49 29 29 29 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1a 1a 1a 37 37 37 36 36 36 38 38 38 39 39 39 39 39 39 3a 3a 3a 3e 3e 3e 3f 3f 3f 41 41 41 41 41 41 43 43 43 47 47 47 48 48 48 49 49 49 49 49 49 4d 4d 4d 4d 4d 4d 4b 4b 4b 39 39 39 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 34 34 34 40 40 40 43 43 43 45 45 45 47 47 47 47 47 47 42 42 42 42 42 42 41 41 41 41 41 41 40 40 40 42 42 42 43 43 43 46 46 46 4a 4a 4a 3d 3d 3d 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 2b 2b 2b 39 39 39 3b 3b 3b 3a 3a 3a 3b 3b 3b 3c 3c 3c 40 40 40 41 41 41 3f 3f 3f 3d 3d 3d 40 40 40 40 40 40 42 42 42 44 44 44 45 45 45 49 49 49 49 49 49 48 48 48 3a 3a 3a 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2b 2b 2b 40 40 40 44 44 44 49 49 49 48 48 48 46 46 46 3f 3f 3f 40 40 40 41 41 41 41 41 41 3f 3f 3f 41 41 41 43 43 43 45 45 45 42 42 42 1a 1a 1a 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 10 10 10 34 34 34 3b 3b 3b 3b 3b 3b 3b 3b 3b 3c 3c 3c 3e 3e 3e 40 40 40 3d 3d 3d 3c 3c 3c 3e 3e 3e 3e 3e 3e 40 40 40 41 41 41 43 43 43 44 44 44 45 45 45 43 43 43 38 38 38 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2b 2b 2b 44 44 44 4b 4b 4b 4b 4b 4b 45 45 45 40 40 40 41 41 41 3f 3f 3f 3f 3f 3f 3e 3e 3e 3d 3d 3d 41 41 41 43 43 43 49 49 49 27 27 27 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1b 1b 1b 3c 3c 3c 3b 3b 3b 3c 3c 3c 3c 3c 3c 3c 3c 3c 3e 3e 3e 3c 3c 3c 3c 3c 3c 3f 3f 3f 3b 3b 3b 3e 3e 3e 40 40 40 43 43 43 45 45 45 47 47 47 42 42 42 3b 3b 3b 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 29 29 29 45 45 45 49 49 49 44 44 44 41 41 41 3e 3e 3e 41 41 41 3f 3f 3f 3d 3d 3d 3e 3e 3e 3d 3d 3d 3e 3e 3e 40 40 40 26 26 26 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 26 26 26 3a 3a 3a 3c 3c 3c 39 39 39 3b 3b 3b 3d 3d 3d 3b 3b 3b 3c 3c 3c 3d 3d 3d 3d 3d 3d 3e 3e 3e 3f 3f 3f 43 43 43 43 43 43 46 46 46 42 42 42 3c 3c 3c 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 26 26 26 43 43 43 41 41 41 42 42 42 42 42 42 3e 3e 3e 41 41 41 40 40 40 3e 3e 3e 3d 3d 3d 3e 3e 3e 3e 3e 3e 20 20 20 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 23 23 23 39 39 39 3a 3a 3a 3d 3d 3d 3c 3c 3c 3b 3b 3b 3a 3a 3a 3d 3d 3d 3b 3b 3b 3e 3e 3e 40 40 40 42 42 42 44 44 44 44 44 44 41 41 41 3d 3d 3d 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 23 23 23 48 48 48 4b 4b 4b 4f 4f 4f 51 51 51 4d 4d 4d 4a 4a 4a 45 45 45 41 41 41 3b 3b 3b 2d 2d 2d 14 14 14 04 04 04 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1b 1b 1b 35 35 35 3d 3d 3d 3c 3c 3c 3c 3c 3c 3c 3c 3c 3f 3f 3f 40 40 40 40 40 40 42 42 42 42 42 42 44 44 44 46 46 46 42 42 42 3d 3d 3d 06 06 06 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 33 33 33 74 74 74 77 77 77 7c 7c 7c 7c 7c 7c 7b 7b 7b 77 77 77 69 69 69 50 50 50 1f 1f 1f 06 06 06 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 14 14 14 37 37 37 42 42 42 48 48 48 47 47 47 4b 4b 4b 4d 4d 4d 51 51 51 55 55 55 55 55 55 57 57 57 5a 5a 5a 59 59 59 56 56 56 09 09 09 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 2c 2c 2c 6a 6a 6a 6c 6c 6c 6e 6e 6e 6a 6a 6a 63 63 63 54 54 54 33 33 33 10 10 10 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 04 04 04 10 10 10 3d 3d 3d 60 60 60 6c 6c 6c 72 72 72 74 74 74 76 76 76 74 74 74 74 74 74 72 72 72 6d 6d 6d 68 68 68 5f 5f 5f 0b 0b 0b 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 1f 1f 1f 4f 4f 4f 4b 4b 4b 41 41 41 30 30 30 1e 1e 1e 0c 0c 0c 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 0a 0a 0a 29 29 29 4a 4a 4a 5e 5e 5e 60 60 60 5c 5c 5c 54 54 54 58 58 58 59 59 59 58 58 58 52 52 52 4a 4a 4a 0b 0b 0b 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 08 08 08 13 13 13 0b 0b 0b 06 06 06 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 16 16 16 1f 1f 1f 1e 1e 1e 10 10 10 21 21 21 22 22 22 1d 1d 1d 16 16 16 10 10 10 04 04 04 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 02 02 02 03 03 03 03 03 03
