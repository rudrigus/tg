 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 0d 05 03 00 06 05 03 00 06 05 05 01 06 0e 0a 0b 09 05 0c 05 0d 07 08 14 19 24 27 22 18 1a 1e 28 29 17 2e 2f 38 35 2f 2b 34 39 49 44 33 42 4c 49 3e 48 45 45 4a 42 43 4e 4e 4f 53 54 49 3e 3d 49 5a 34 2a 22 21 28 21 25 29 2a 3a 3f 3b 42 35 36 1a 1f 25 1f 1b 1d 1d 23 1b 0f 19 12 11 13 06 07 12 14 0d 02 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 00 06 05 06 03 06 05 12 16 14 09 05 08 06 0a 09 14 06 0a 0d 05 0d 13 13 1a 25 23 20 11 19 19 13 25 24 31 31 3c 3d 2c 33 3f 3f 34 42 43 50 43 47 4b 43 44 54 49 54 54 53 5b 52 59 54 58 5c 69 62 63 6b 62 67 62 50 54 57 73 6c 54 48 43 3c 3b 35 38 3e 47 47 61 65 62 69 63 43 31 3e 45 43 37 28 2a 2b 2a 24 2c 19 1b 15 0f 1a 22 1a 1d 11 15 17 14 0d 07 0b 05 0f 06 06 0f 12 05 04 02 06 12 0a 00 06 05 03 07 09 05 03 00 06 05 0f 0e 08 05 07 00 06 05 03 05 06 08 05 05 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 0d 1a 15 11 00 06 05 03 09 06 17 0e 10 0e 13 1f 1f 13 0b 0c 10 15 1c 19 25 45 49 2d 0f 10 1f 1e 22 28 33 46 48 44 3d 38 4b 4f 45 46 56 54 4c 45 55 6d 69 64 61 56 5e 66 67 66 68 68 6e 81 92 8c 92 8e 8b 80 78 70 70 79 94 97 7e 73 63 59 5f 52 4a 56 54 54 63 69 89 7c 69 4f 4e 53 54 4d 4e 43 44 33 3b 38 37 41 36 32 27 29 34 2d 2f 22 25 28 25 16 1c 14 18 0f 05 09 0b 0a 0f 13 09 06 11 03 02 06 07 09 00 06 0a 06 02 08 0b 03 0f 06 05 0a 01 06 06 07 04 09 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 06 05 0a 16 2c 27 24 13 12 06 03 0b 06 09 14 10 06 0b 10 1a 15 10 0f 14 0d 1e 19 23 36 35 2d 22 1f 25 1b 2b 46 64 56 50 4f 42 43 50 54 57 66 71 72 77 76 89 a6 9b 97 8d 92 8e 91 97 9b a2 a7 af be d4 e1 dc d1 d0 c4 b9 ba b4 bd c4 c8 bd a4 a0 9c 8d 7f 7a 80 79 76 79 7b 8b 7c 72 77 76 6f 72 71 72 68 58 50 4c 4c 54 52 46 3c 3b 35 40 3a 49 4b 46 53 49 38 3b 34 32 34 21 26 1e 1a 19 11 13 08 14 0b 18 0e 0f 11 08 0b 0c 08 0c 08 11 09 0e 0f 0e 0a 0d 06 06 06 03 09 05 03 05 0a 0d 03 06 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 06 0e 23 1f 1f 12 11 0c 06 00 06 14 0f 0c 0e 0e 07 19 1b 22 26 1c 1a 1f 24 1e 25 22 25 2a 36 34 30 41 5b 70 6c 61 56 56 69 7c 7e 89 a9 b3 b5 c1 d4 e7 f5 f5 eb d7 d8 e2 e3 e2 e6 e1 ea f0 f0 ff ff ff ff ff ff ff fd fa f9 e7 ea e6 d4 d6 cf c9 c7 b7 b9 ad aa a3 96 8a 92 8e 95 92 9a a8 a7 a4 a1 90 80 76 6b 6c 61 62 43 3c 3b 44 47 49 45 4d 53 55 56 5c 4f 54 50 44 3f 41 3d 39 2d 25 1e 20 21 1e 1c 1e 16 11 12 10 06 10 09 10 0e 0a 0b 0c 0f 08 0b 0e 11 10 07 09 03 07 06 07 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 0b 21 17 0b 0b 0f 05 03 0b 12 07 12 10 0e 16 18 12 19 21 1c 19 2e 2b 2e 26 25 2e 46 42 55 4b 51 5f 6b 89 98 90 93 8d 99 ae b6 d3 e3 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 fd ff ff fd fa f0 e4 d2 de c0 b9 b9 b5 af ab b3 bb c6 ce cd bb b8 aa 97 7f 6f 60 4d 54 4b 45 3f 4f 45 4e 51 56 38 60 5e 5c 62 58 5a 59 5a 52 54 4d 4f 46 44 42 35 34 2c 1d 25 1a 1e 18 1a 18 14 18 11 1f 0e 1a 0d 0d 0f 0b 09 0e 03 0c 0b 05 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 10 12 1a 33 29 0d 0b 0c 07 14 13 0d 0b 11 14 17 1c 23 29 27 26 34 37 32 36 38 40 3d 43 52 5a 6e 6f 79 80 94 a3 b5 ce d1 c0 cf d2 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f2 ed e0 de d3 d5 d9 d0 d8 d5 d3 cc c3 b7 99 8c 7f 75 61 5a 4f 4f 50 4f 52 4c 5c 60 6f 67 60 59 64 61 59 5a 5b 59 5a 5e 67 64 64 65 66 57 57 51 3e 40 39 35 35 24 23 23 16 17 13 1c 14 0a 15 0d 09 0e 07 03 06 05 0b 14 09 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 07 06 18 06 15 20 1b 15 0f 09 15 20 24 25 18 1e 20 21 38 36 31 34 48 5f 64 58 50 4c 53 5a 63 75 82 89 95 ac ba c6 d1 e0 f0 e8 e6 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ee eb ec ec e8 e3 e1 d2 c7 be a0 8c 82 7e 6a 66 62 61 5d 60 59 54 5a 64 69 6d 73 68 6b 6b 65 5f 60 5b 5d 5f 67 63 6a 67 68 71 7b 6f 76 6d 68 65 57 4a 48 39 33 34 1b 25 1e 20 1f 1d 18 0d 10 0e 12 0c 07 12 08 07 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 08 0b 0a 07 11 0b 12 14 11 16 16 19 2f 30 25 24 2e 35 3e 40 37 46 52 6c 99 9f 77 64 6d 71 7a 91 9e aa c4 d3 e2 dd dd ed df e9 eb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff fc f8 f1 e8 df da ce b8 a5 a3 8b 81 6f 65 70 67 65 63 65 64 6a 6c 6d 6c 6d 67 66 62 5d 68 59 57 5c 55 60 68 63 7a 71 6e 75 83 84 8d 82 85 84 73 68 61 52 42 37 2a 27 28 21 26 1c 12 0f 0a 0e 0a 0c 08 09 03 00 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05
 03 02 0b 07 05 09 06 05 07 0f 06 0c 09 0a 0a 06 0e 08 0a 07 0e 22 22 20 25 2d 28 2c 3b 36 40 40 51 5a 54 52 4f 5e 6a 99 ae a5 93 92 8a 98 a2 b0 c4 d3 d9 d9 d4 d0 c4 d0 e0 e5 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ee ed e4 d4 ca b2 9d 8d 82 81 79 77 7c 7b 6e 6a 76 6d 72 71 74 76 65 68 66 60 64 62 5e 54 61 5c 68 6f 6e 6d 70 90 9d 9d a1 9b 9e 9f 99 9e 8f 81 79 67 5c 44 3f 38 27 1b 1a 1e 18 0e 11 11 11 0a 0f 08 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 09 06 09 09 00 06 0a 0a 08 07 0a 05 0c 15 05 0a 0e 11 18 1b 29 3b 3e 49 43 3f 3b 38 45 43 59 5f 6c 76 72 70 72 85 92 9f a3 a3 9d a1 a9 9e b2 c1 c2 bb c0 b8 b3 b6 be cf d6 e0 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f7 e0 c7 ad a8 9c 95 8e 84 87 89 82 7a 7c 77 7f 79 75 70 6b 67 6c 6c 69 6d 58 68 5d 65 67 6b 61 6e 73 85 a5 b8 b4 be bc b8 b8 b9 b2 b4 b3 ae 94 7d 76 5d 48 46 39 26 1e 12 12 17 0d 0c 0f 06 09 0c 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 03 05 06 05 03 02 06 05 03 08 09 05 08 04 06 0c 0b 0b 10 10 09 13 1c 29 33 3e 49 4e 62 5d 52 54 59 60 61 67 66 6b 7c 84 87 81 93 97 98 9f 97 9c a3 9b 9f a5 a8 a9 a3 a1 ae af af af c6 d3 d5 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e1 cc ba af a7 9f 9e 96 88 8a 8b 8d 87 80 81 74 72 72 77 73 6e 6e 6e 6e 65 6d 6a 6a 72 6f 69 75 81 99 b2 b8 c2 c6 ca c7 c0 d4 ce d3 ce cf c0 b5 96 87 75 65 4b 35 2d 15 08 05 0c 10 09 05 05 0b 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 06 05 0d 14 14 05
 07 07 06 07 03 0a 0d 0e 0a 0c 0e 13 1b 1f 28 24 28 30 31 3e 43 49 61 68 6c 69 6c 6a 6a 6f 73 75 7a 7c 87 88 85 8b 8a 94 95 94 96 98 91 8f 97 95 9c a7 a6 b2 aa b3 b8 b7 ca d2 d6 e9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd e6 ca c7 ba ab a9 a7 99 a0 92 9c 91 8d 8d 8e 8b 83 7f 7b 7b 78 7c 72 72 75 6c 6f 71 73 76 77 77 8b a3 c1 c6 cb d5 da dc e5 e9 e0 e9 e0 de d3 c6 b8 a5 a1 84 62 45 2e 24 15 18 15 16 0f 08 01 0b 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 11 0e 0e 05 08 06 0b 0d 10 13 16 0a 10 1f 1c 32 3a 40 38 35 42 38 44 4f 5d 6a 74 75 70 78 75 70 74 7a 7d 84 83 86 84 88 94 8f 8e 95 96 9e 98 95 9f a2 ad a8 b6 b6 b1 bd b6 c1 c6 d3 d4 dd e0 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e2 d0 c9 bc bc b4 a1 ac a0 9f 9d 9d 93 95 95 89 8f 88 85 80 87 7a 71 75 79 7b 81 80 7e 7e 86 81 8d ad b7 c9 db db e7 ee f8 fb f2 f5 eb df d9 d2 c2 b8 aa 94 6a 51 46 3c 2f 27 13 15 0e 07 09 0c 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 04 04 06 05 0b 0c 06 0c 09 0e 11 1e 1c 28 32 3d 3f 48 46 45 46 4c 47 4d 57 5b 65 62 6f 70 65 6a 6c 74 81 87 8b 8c 8a 8f 8f 91 94 90 9a 9b 9f a2 9d a2 ae ae b7 ba c3 c4 bf c9 cc d4 dd df dc de f2 ed f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 db d5 c2 c1 b6 af ae a7 a9 aa a1 a2 9d 9a 98 95 87 8c 89 7b 7a 89 7a 83 80 80 83 84 89 8b 8d 99 ab b5 ca dd de f1 fb ff ff ff f9 ec e8 e0 d6 d8 c2 ad 97 8f 7d 72 63 51 35 1b 0b 0b 08 05 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 06 03 0a 0c 06
 09 18 11 14 12 18 1d 2a 3c 3c 41 49 4a 50 4f 54 5e 5f 61 5b 5b 5f 6a 62 66 66 6a 75 7c 83 85 88 97 94 9b a4 a7 a0 a4 a6 a4 9c a5 a3 b4 b2 af c2 c7 cd d6 d0 d8 e1 e9 e8 f1 e2 e4 ed ec ea fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 de cf c6 c4 b7 c4 bf ac b2 ad ab af a5 a4 94 8b 93 96 82 87 86 92 8c 8d 85 8e 8f 91 8d 93 9e a3 a6 c6 d2 e8 f9 ff fc ff ff fe fd f5 eb dc d6 d1 c7 bc b0 a7 9d 8f 8a 6f 51 2c 15 0e 05 03 06 06 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 09 0a 09 11 0c 08 14 16 1b 19 25 2c 30 45 51 50 61 5f 67 5f 66 68 61 63 6d 62 64 5e 5f 69 6a 72 6d 7d 84 87 92 86 94 94 9f a1 be b0 ba b1 bb b3 ae b5 af bc ba c6 cd d0 d6 e0 df ef e4 f7 f2 fa ff f9 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e4 d9 c8 ca c9 c4 bc ba ae af a7 b1 a7 9f a2 9a 9c 94 92 89 8d 97 95 91 8c 93 95 92 98 94 90 ab b5 c3 e2 f3 fa ff ff ff ff fc f1 e6 e4 e5 da d7 ca c2 be b6 a6 9f 98 84 5d 2b 0a 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 04 06 05 03 00 0a 05 09 04 06 0d 0e 03 0a 18 22 34 3b 4b 50 49 62 6a 76 86 7e 7e 73 73 75 6b 6a 6b 6d 64 5e 5f 75 75 75 86 8a 8c 8d 8e 94 a3 a7 ae b9 be bc c1 bf c4 c0 c3 bd bc c5 c5 ca d4 d3 e2 e7 ef ef fd f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e6 e1 db cd ce cb ca bf be b5 a1 a7 9d a1 a2 9a 95 99 93 8f 94 9d 9d 95 93 95 9b a2 a2 ad b4 c9 e3 f1 ff ff ff ff fc f8 f2 ed e4 ed e6 de cd cf be b8 a7 a3 a9 97 7b 55 26 0c 03 05 06 05 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0c 0e 08 18 13 1a 1e 2e
 3e 50 5f 6d 6f 73 79 84 8d 8c 88 8f 85 87 80 7e 75 6a 6c 65 6f 70 79 70 78 86 90 9a 99 9d a5 a6 b3 be cd c7 c5 ca cd cb cc ce cc cd d0 d0 d2 db e0 e6 f2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ee ea e6 d9 e0 d9 d3 d7 ba be af ae a9 ae 9b 9d 9b a0 9f a2 9c 9d 98 9b 9a 9e a6 a7 ad b5 bf d8 ee f4 f5 ff fd f3 ed eb ea ec f1 f1 e4 dc d7 cf c5 a9 ad ae a0 84 78 3b 16 03 00 06 05 03 08 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 07 05 06 05 07 08 07 10 0d 0b 10 19 20 33 3b 52 6e 80 8a 99 93 96 89 8e 92 95 94 8f 8f 8f 8d 84 7d 78 74 72 76 78 7f 84 8b 91 9c 98 a1 a3 b0 b1 ba be c7 cd d1 d6 d7 cc d6 ce d8 dd d9 df e2 e2 e7 ef fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f4 ea ef de e3 d5 c9 be b2 b1 a6 a9 a5 a7 a0 a0 a9 a6 a0 a3 a1 a5 a9 af a1 ad bd c4 d3 df ec f0 f6 f2 ef e0 f1 ef f2 fa f9 e4 e7 dd d3 cb b9 b5 b1 a1 8a 7c 54 1a 0d 06 06 05 03 00 06 07 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 08 03 0c 08 07 12 1b 1e 2f 3e 3c 58 6d 92 a4 b3 b4 b8 ab 9b 8f 93 9a 97 8b 8d 8d 97 8b 85 71 72 77 74 7d 80 89 8e 95 99 a6 ae ac b2 b4 b4 bb c8 cf db d7 da dc da e1 de dd e1 e5 ea ed f3 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fa f2 ec db d3 c9 c3 b6 b1 a8 a1 ad a9 ab ae a9 a3 a8 a6 ab ad aa ae ad b5 ba be d1 e5 e7 e7 e8 ea eb eb ea fa fa f5 ee e1 e0 cf ce c3 b7 b3 ac 96 8c 5b 2f 13 0a 0a 05 05 0b 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 03 01 06 08 0a 0a 13 1e 27 36 36 45 47 54 6a 85
 a6 c1 cc c8 be bd a1 8e 88 92 96 93 92 90 90 95 8d 7c 82 86 85 8a 88 8d 92 9c 96 a8 ad b0 b2 c1 c4 c9 ce dd d7 df e1 e9 ec e9 e6 e7 e3 ef ed f2 f9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f3 ec e2 dd d2 c8 bf b9 b6 ae b5 b0 af af b2 a9 a3 a7 ae a5 b1 b6 b4 ba c5 c8 d4 da e1 da e4 e3 ee f5 f5 f3 f5 f0 ea ef e8 dd d5 cb c1 b3 aa a0 92 7d 49 1a 11 08 05 03 07 06 07 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0a 06 05 0c 07 0e 0c 1b 22 2f 3c 40 3f 42 45 52 58 6e 82 a3 be cc cf bd b0 9e 9a 96 9d 94 90 97 96 9d a4 8f 85 86 84 89 92 94 97 a0 a5 a8 ac bb c4 c2 ca cd d0 d9 db d8 e1 e4 f1 f3 ef fe f2 f4 f4 ff f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f6 e9 e3 e2 d5 ca c2 bd af b1 b7 be b8 b6 b4 b5 b5 b7 b6 be ba c1 c5 c0 c8 c4 d7 d9 dd e6 f2 ee ea f1 e2 f7 eb e7 e5 ea dd ce ca c3 bf ac b0 a9 a0 72 41 1f 07 0b 0d 0a 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 07 08 06 0c 0f 15 22 2c 36 42 42 44 3b 44 43 51 55 5f 76 75 96 ab b0 c4 b4 a6 a6 a2 9a 9c 90 91 a0 9e a3 99 8c 8e 88 93 8a 99 9b 9c a3 a4 a7 b6 bc c7 d2 cb d7 d7 dc df e2 e4 ed f1 e9 f4 fb f9 fd fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 f4 f8 f7 ec f0 d4 cf c0 bf c1 ba c1 b6 bd bc c1 c2 c2 c9 bc c7 ca c8 ca ca d2 cf de e3 e3 f2 ef ef e9 eb ed ed ed e7 e5 d4 d5 c6 be b9 b5 be b6 af 90 5d 2e 19 09 09 0a 07 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 04 05 0e 05 0a 11 15 19 24 3b 51 41 4d 50 45 48 48 4b 49 52 60 6a 6d 81
 89 9b ac b2 ad aa aa a1 98 9f 92 9a 99 96 93 8c 8b 8f 8e 9c 9e 9e 9b a6 a6 ac b5 bd c8 ce ca d5 d7 d5 d3 df e3 e1 f0 f0 fb ff ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 ff ff f8 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff ff ff f5 e4 e1 e9 f7 ff ff fa e8 e3 d7 c3 ca c0 be c8 c1 c4 c6 bb c0 c1 c7 cf c8 c2 c9 c8 d4 d7 dd db db e7 ec ec e5 ec ed e7 f0 e0 df db d1 c4 ba ba b6 b7 bf bc a4 7b 48 1e 0b 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 07 0e 19 15 1b 31 35 44 54 5b 5e 58 55 52 53 46 4c 4f 51 5d 6b 65 7a 84 87 95 a2 ac b9 b2 aa b0 a6 a4 9e 95 9b 9b 92 95 9d 9d a1 aa a0 ab b3 b9 bb bf c1 cd d1 d0 d6 d7 d8 d2 d5 e0 e1 df dd ef f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc f9 f9 ff ff ff ff ff ff ff ff ff ff fc fe ff f8 ff ff ff ff fa e7 e7 e6 f1 fb fb f6 ec c1 e0 de e1 d6 cd ca c7 cb cb c4 c3 d1 d2 ca ce d4 ca d6 d4 db e4 e5 dd e3 e7 e9 ed df e0 e5 e9 e4 df dd d1 c0 bb bf b5 c0 cb c5 b0 98 6c 3b 20 10 0d 06 05 03 07 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0e 05 0f 12 21 3c 40 4d 5b 5d 69 6f 68 5f 54 50 51 55 54 5a 5b 66 5f 66 7e 86 8e 98 a1 ae b5 b3 b6 b0 a7 a2 a6 a1 a3 9a 98 9c a5 a8 ae bc b5 bc c2 c0 d6 ca d3 cf d1 d9 d2 d5 d3 db d6 e3 e2 e0 ee f5 f8 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fd fd f7 f5 fc ff ff ff ff ff fd ff fb fb fa fa fa ff ff ff f8 ef ec ed ea ea f8 ed e9 f8 ef fc fb f6 ea e0 d1 d2 d5 d2 d6 d6 cb cb d7 d2 d2 d7 d5 df dc df da df e3 e5 e3 e2 e0 e2 e4 e1 d7 d4 c0 bd b4 b0 be c4 c6 c4 bf a3 87 5d 2e 1f 05 06 0d 03 05 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 0d 20 43 4c 55 60 5d 73 77 70 68 63 59 51 54 4c 58 5f 5b 60 69 6e 81 90
 9c 9c a3 b5 b7 b4 b4 ad ae b1 a7 b4 a3 a6 a6 ab ae ad c1 c7 cb c9 d9 da d7 d0 d9 d5 da d5 d7 d4 d4 d3 d9 d8 d7 e1 df f0 f7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff fe f7 fc fc ff ff ff ff ff fd fb fa ff ff ff ff ff fc fe ff f8 f4 ee eb ee ea ed f2 eb ff ff ff ff ff ff ff f9 e2 db d5 d0 cc ce cf de d9 d6 d4 ce d0 dd d6 d7 de df e4 dd d1 da db e4 e1 d8 ca bd b5 b1 b4 c5 c7 cb d7 c6 b5 92 75 55 26 10 06 05 08 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 01 06 05 05 05 0a 12 18 2b 44 58 64 6c 71 78 80 79 66 5b 5e 60 5f 61 64 66 66 70 6f 74 90 9f a0 ac b0 b0 b5 b9 b3 b3 ac b2 ae b6 b2 af b5 b5 c2 c3 cc de d9 e0 de e4 e3 dc dd e1 de e4 db d1 d8 d6 d7 dd d4 db e5 e8 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fe ff ff fd ff ff ff ff fc fa fc fc ff fa fe fa fa ff fa fc fa fc f3 f3 ed f4 f5 f6 f5 fc ff ff ff ff ff ff f1 dc d2 d3 d1 d7 d7 df dc d7 e1 d5 d3 d9 d3 df e0 db df e0 d5 da d9 d4 c8 c6 ba b0 bb c3 d0 cd d9 dc d0 b4 9c 7f 66 3f 21 10 09 03 07 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 0f 0c 11 1b 29 53 65 6f 72 7d 83 7d 79 7a 5f 66 6f 63 6c 6c 70 71 74 78 75 94 b3 b5 b5 b8 c0 c1 c3 b6 c1 b0 b6 ba c2 c4 c2 c5 be ca cf dd de e8 ee f1 e3 f3 e7 e7 ee e8 e1 e3 e4 d9 d2 da d8 e1 e5 e8 ec e9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff fd fc ff ff fe fc ff fd ff f5 fd f9 fe ff ff ff ff ff ff fb f9 fb f1 f4 f4 f4 f1 ee ef f1 fe f8 ff ff ff ff fd ea d7 d1 cd d9 e8 dc d5 d6 d5 d9 ce d6 d5 da d8 dd d7 da d6 cc d1 d2 cb be ba bb c1 c9 d2 ce d5 d3 d0 b9 98 7e 74 4a 25 1b 0c 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 06 0f 13 15 2d 4b 64 6e 69 7b 79 86 92 8c 7e 77 78 77 6b 6e 6a 6b 6a 79 80 89 a1 b7
 c2 ba c1 c3 c1 c3 c9 c1 b7 c4 c6 c4 ce d0 ce d3 d1 e1 de e8 f2 e9 f6 f1 f3 f1 ef eb ec e4 e4 e5 df da d8 dc d9 df e8 ea f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f8 fb ff f9 ff ff fc ff ff ff fd f9 fa fb f9 ff f9 ff ff ff ff f6 f3 f4 f5 f9 f6 e6 f6 f5 f8 fa ff fc ff ff ef dc ce da dc e5 de dc d4 d7 d9 d5 d1 d7 d7 d6 d6 d8 d2 d2 cc d3 cd c5 cc c4 c1 cc ca c6 c5 cf db c3 a9 99 84 7d 58 3e 25 0f 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0c 06 05 0c 19 20 37 62 78 6f 66 76 7c 81 8e 8e 92 85 77 74 7b 79 7a 75 71 7a 7e 78 91 a6 c1 c1 b9 c7 cc cb ca cd cd ca ce d6 d0 dc d0 d6 d5 e9 e9 f2 eb f5 f6 fe fe ff ff f5 fd f4 f1 f0 ee ed e0 e3 e0 e2 e7 ef eb f5 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff ff f7 fc fc fa ff fa ff f9 f0 fc ff fb fe fe ff ff ff ff fc fa ff f4 fe f9 f9 fd f9 ff ff fd fb fd fa e3 da e8 e2 e3 e8 db e0 ec e3 df d6 d8 e0 d9 d3 d4 d1 dc d3 d3 cc c7 cb cd c9 d3 c8 c4 c5 cf d2 ba 9d 86 85 84 7a 51 37 1c 0d 01 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 16 29 34 64 8a 80 80 76 7c 81 91 97 9a a0 99 83 7e 7d 82 7f 85 7d 82 84 92 9d b8 cb d1 cd ca cb ce d2 dc d3 d7 dd df dc e1 e8 e4 eb e5 e9 e9 f2 ff ff ff ff ff ff ff ff f8 fc f3 f9 f5 e7 e5 e5 e2 ec e5 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd ff fd ff f9 fd ef f7 f7 f5 f9 f9 ff fc fd ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff fe ee e1 e0 e9 ee e6 e5 ed ee e5 e5 e6 d7 db de da da d9 db d9 d5 ca d4 ce d3 d5 d0 c7 b9 c4 c5 c5 ac 97 8a 83 95 98 72 4b 21 07 00 06 05 06 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 0b 0f 08 07 11 12 2a 5b 8f 93 7f 79 84 89 92 90 9a 99 9c 9a 8e 86 85 93 8f 8c 8d 87 91 97 a9 d4 e3
 df d2 d3 d3 d2 d3 d5 d6 da e1 de e9 ea e2 f3 e9 e6 ed f6 f8 ff ff ff ff ff ff ff ff ff ff fd f5 fb f3 f2 e4 e8 f4 ec fd fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f9 f6 fb fd f5 f5 f0 ee f1 f6 f5 f2 f1 fe f9 f3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee e3 e9 e9 f8 fc fe ff ff ff ff f9 e8 e7 e0 e2 dd e2 df d1 d3 d0 d0 db db d9 d9 c0 bb b9 b7 bf ad 95 8b 84 98 af 95 59 25 14 06 06 06 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0b 06 05 0a 0f 19 0e 22 47 7d 98 95 7f 7e 8c 90 9d 90 96 92 9e 90 94 97 8e 93 98 92 92 8e 9b ab c0 f0 f9 e7 d9 d3 d0 d3 d7 d9 dd dc e4 e2 eb ed ef ed f0 f7 f6 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f6 f7 f6 f0 f4 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fb fe ff fc f8 f1 f4 f0 f2 ec ed f2 fa f1 f6 f8 f6 f6 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f8 fc ff ff ff ff ff ff ff ff ff ff f3 ec eb e7 e4 dd cc e2 df e6 db de d7 d3 c4 c0 b4 b8 ac 97 97 91 8b aa bb a0 69 35 19 0e 06 06 06 04 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 02 06 10 16 14 1e 25 32 52 8f 95 91 8a 8a 9b 99 98 98 9d 9a 9f 95 9a 9d 9a 9f aa a6 aa ab aa b9 e1 ff ff fa e6 da da dc d8 de e4 e2 e8 e8 e8 f2 f1 fb ff fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb f4 f2 f3 f6 f3 f2 ee ec f8 f0 f0 f5 fc ff ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f0 e3 f0 e4 e9 ea e1 d0 cd c3 b8 b3 a7 aa a8 9b 8f 92 a5 c6 b3 89 50 24 12 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 08 0f 11 12 19 1a 24 40 70 8a 96 90 89 8e 99 99 98 99 9b 99 95 9e 96 a4 a2 a2 aa b0 af b5 ae ca ef ff ff
 fe e3 df de dd dc e6 e6 e8 ee ed ef ee ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fb f5 f6 f5 f4 ee ef ee ea ec e7 ef f2 f6 fb fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f5 e8 ec ea e1 ca cd bd b5 b0 ab a6 a5 9b 92 a1 c0 c1 b1 a1 62 3c 1c 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 06 09 03 0d 10 10 12 1a 23 35 5d 8a 8e 96 97 94 95 97 a4 9d 98 98 9d 9d 97 a3 a2 a8 ab b7 b1 b3 b7 bd d5 fe ff ff ff f0 ec e2 e4 e4 e7 e7 f3 f5 ef f5 f4 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fb fd f8 f1 f3 ed ec f1 e5 eb e5 ea ed f5 f8 f6 ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ea f5 f2 dd d6 cf cd bc b8 b0 a1 9a 9f 9a 92 9f bc c1 b6 a9 76 46 2d 0b 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0d 0d 13 27 2c 38 55 86 96 8f 92 a4 a4 a1 a5 a3 a0 9f 9a 9b a0 a1 a0 a5 b4 b9 c0 bf bb b9 c8 e2 f7 ff ff ff f1 ec e6 eb f2 f4 f5 f6 fd f7 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 ff fd fd f9 fc f1 f0 ec e5 ea ef e8 e7 f5 f1 f6 ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e2 d6 cb c6 bc b3 ab a0 a6 9a a0 99 a2 b5 be b4 b6 93 5f 3c 10 0f 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 0b 0b 0c 1a 1a 25 30 52 74 8e 90 98 9f a8 a9 a0 a2 a0 a4 9e a1 8f 9d ae ac a4 b2 b4 b1 c4 bc d2 f7 fe ff ff ff
 ff f3 ed e8 f5 f6 fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fe fa f7 f9 f5 f7 f2 f1 eb e5 f0 f0 eb f2 f6 f9 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 e6 dc cc cb b6 ad af aa a6 a3 9c 9b b5 c5 c8 c9 c4 b3 7c 49 22 09 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 06 02 0a 06 0c 0b 13 28 32 47 75 8d 95 95 9b ad ab a5 9a a0 a6 9e 97 9a 9e a1 a5 a4 ac ad b6 c0 c7 e6 fc ff ff ff ff ff f3 f8 f5 f5 fe f5 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ff f3 f5 ef fe fa fa ef f0 ed e6 ea ec ef f1 f9 fe ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 d4 ca cb b1 b0 ae a8 9c a0 98 9e bb c5 d4 d7 d3 c6 9e 5b 1a 0a 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0d 08 0e 21 1b 30 4b 6d 8f a8 a7 9c 9e a4 b2 a4 a5 a2 a8 9f a5 93 9c 9e ac ae b3 b2 be d1 eb ff ff ff ff ff ff f9 fa fc f9 f4 f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f5 f0 f8 ff fb f6 ec ed ee e9 eb ee f6 f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e2 c0 be b5 b5 b2 a8 a3 a2 a0 aa b7 c4 d8 dd db cc a1 70 30 0c 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 06 0a 09 0b 19 1e 2f 3f 6a 88 a7 b5 a2 9d a4 a5 b3 ab a4 a8 a4 a9 9e 9d 94 a3 aa b5 b3 b4 c2 ce f6 ff ff ff ff ff ff ff
 fb fa fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff ff f3 f9 fc fd f4 ee ea ee eb f5 f3 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 d3 c9 b8 b7 aa b3 a6 a4 9f a2 af b7 b0 c6 d1 d7 c3 aa 73 31 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0d 0d 0c 0c 1b 26 41 61 89 a1 bb b6 93 a0 9f ae bd ad aa a5 aa a2 a3 9a a1 ad ad b2 b8 ba c7 d3 fc ff ff ff ff ff ff ff ff ff fc fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f8 fe ff ff fd f2 ed f0 ef f5 ef f4 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb d4 c2 ba b1 b4 ab 9f 9f a3 a6 ac b1 b0 b0 c6 c7 bc a1 73 30 0e 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 06 05 11 0c 1e 44 57 7a 9d b5 d5 c1 a4 9e a6 b3 bb b2 b0 a5 a7 ae a3 a6 a9 a7 a9 b7 bb bf d0 e4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f0 f5 f0 eb ff fb fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff eb db c3 ba b6 b0 aa a9 9d b2 b8 b4 b2 b5 b1 ac bf ba a5 79 36 10 09 03 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 06 0e 0e 0e 13 14 30 4f 7b 95 ae cb e3 c5 ad a5 ab af ba b9 b2 ae ac b0 ac b3 b3 b7 af b5 b3 bd d5 ec ff ff ff ff ff ff ff ff
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f3 f6 f9 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 dd c3 cc c0 c3 be af ac ac b5 b0 b8 bb af ab b2 ac a8 78 33 15 09 01 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0c 0d 1f 31 5b 8e a5 be d8 f1 d4 af af ad af bf c1 ba af b0 b5 b4 b2 b3 b2 b9 b4 b6 be d9 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec e3 e2 da de de d2 b9 b5 b3 ab b9 be b2 ac a2 9d a5 9a 74 3b 14 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0d 0e 17 25 3b 6f 97 bc d4 e9 fa d3 b2 b2 b0 aa c4 c5 c4 bb b5 b2 b7 b6 ba be c1 bb c2 cc d9 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ff ff fa f8 df c9 be b6 b2 c3 b3 b8 b8 a9 9e a5 93 73 34 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 08 07 10 18 1f 35 4c 81 a3 d1 eb fa fd d0 bd b0 a7 b3 bc ca c4 bc b4 bd b7 c4 bc bd c2 bf c6 cf da f9 ff ff ff ff ff ff ff ff
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea d6 c5 c0 bf c0 b8 ba b5 a5 9a 9b 93 67 32 0c 05 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 07 11 10 25 32 5f 8b bc db f2 ff f4 d2 bf b8 b0 af b9 c7 c3 bf bb bd c2 be c6 c0 c6 d3 d1 d9 dc fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dd c7 c2 c0 b9 b6 b5 ab a4 a4 9a 85 51 1f 16 0b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 13 15 1d 36 5c 8a c6 e5 f8 ff e6 ce b8 bd b5 b2 b7 c3 d1 be c0 c7 c3 c5 c8 cf d3 d5 e0 de f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f6 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e0 d6 ca b8 b8 b8 a9 ad a0 a5 97 73 48 20 13 08 01 06 05 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 09 06 0e 11 19 1a 3b 62 8a cb ec ff ff e8 c8 bc bc b5 ba bb c6 cd ca be d0 d5 dd d9 e9 eb ea ea e4 f1 ff ff ff ff ff ff ff ff ff
 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff fe ff ff ff ff ff ff ff ff ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 fe ff ff ff ff ff ff ff ff ff df d9 c0 bf c5 ba b3 a7 a6 a0 90 6b 33 14 0e 0f 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 09 12 11 20 33 5e 8d ce f0 ff ff db cd bd c2 b9 bf c1 c1 cf cb c9 d5 e1 ec fa f8 fb f5 f5 eb e9 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 fc ff ff fe fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fd f9 ff ff ff ff fa f9 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f5 e9 ff fd ff ff ff ff ff ff ff f4 db d5 c4 bf c1 cb b7 a9 a7 97 84 50 28 12 11 0f 06 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 01 06 0a 08 14 27 4b 6a 93 ca f7 fe f0 d5 c0 be c5 c1 be bb c2 cd ce cb da e3 f3 ff ff fb f4 f3 ec f0 f0 ff ff ff ff ff ff ff ff ff ff fd ff fe fa ff ff ff ff ff ff ff ff ff ff ff ff ff fb fa ff ff ff ff ff ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f6 f4 f0 f1 ee ed eb eb e2 e9 ea f4 f1 f0 ec f1 ee f6 ff f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f4 f1 eb f5 ff ff ff ff ff ff ff ff ff f8 d7 c7 bd bf cb c2 a8 a1 93 85 6f 33 1a 14 07 0a 05 0a 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 08 03 0c 06 10 12 15 2b 4b 75 8f cc f5 ff f1 d6 c1 c5 c0 c6 c4 cd cb ce ce d7 de ed f0 ff ff f5 e9 f3 ee ee f0 f9 ff ff ff ff ff ff ff
 ff fd f9 fa fd ff fc ff ff ff ff ff ff ff ff fd fb f4 fb fd f7 fb fa fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f5 f4 ee ea ef ea eb e3 e1 da e0 dc db e3 e1 e4 e0 e2 e6 e5 e4 f3 f4 fa f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fd f8 ef f2 f9 ff ff ff ff ff ff ff ff ff ff e9 cf cc c4 c7 b5 a6 9d 9a 8f 86 64 3d 26 11 0c 06 01 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 0e 0c 13 1c 24 3a 54 76 8a cc f0 f3 e1 d5 bd c1 c7 c2 c7 cd cf cf d5 d9 e2 f5 fb f4 fa f5 f4 eb ed e6 ed f9 fd ff ff ff ff ff ff f7 f9 f5 f7 fd f9 fc fc fc ff fa f5 fd fe fd f6 f0 f7 fa fd ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f4 f1 ee ed e7 e0 db d9 d2 d6 d9 c9 d0 d2 c9 d2 d4 ca cc d0 d4 d4 e1 db e0 db ea f3 f9 f9 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f5 ec fd ff ff ff ff ff ff ff ff ff ff fa e8 d6 d1 c3 b9 a5 9b 94 92 8a 73 4d 33 24 15 14 0f 08 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 04 03 06 09 16 1e 38 65 74 93 c3 f4 f0 e2 c4 b3 ba bf c8 c5 d0 cc d0 da d9 e5 fd ff fc ff fe eb f5 ea e1 e4 e6 f4 f6 ff ff fb ff f7 f8 ec fa f6 fa f5 f6 f0 fa f8 f6 f8 f5 f8 f9 f8 f7 f7 fd f6 fd ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f6 ed ec e2 e0 da d8 da d5 cc cc ca c8 be c1 c5 c1 bc be c1 c6 c2 c6 c5 cc cf d1 d0 d6 dc e3 ea ec f1 f7 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fb fb f6 ff ff ff ff ff ff ff ff ff ff fb f4 e3 d9 ca b8 a1 9b 98 91 90 87 66 4c 2e 31 23 19 10 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 10 13 17 28 42 67 87 95 c7 e5 e7 d7 c5 b4 b7 bd be ce d5 d9 d2 d5 e3 e9 ff ff ff f8 fe ee e9 e5 e3 e0 e0 e7 e8 f0 ed f3 f2 ec
 f1 f0 eb f5 f8 f7 f0 f3 f4 f8 f5 f5 fc f3 fb f2 f9 f2 fd ff ff ff ff ff ff ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 eb e4 db d1 d4 d2 cf ca c0 b7 c1 bd ba b2 ba bd b9 b9 b4 bc bc b4 b8 b6 c2 be c5 c9 c8 d1 dd e5 e1 e8 eb ed fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 ec df db cf b7 ab a4 8f 90 93 8e 86 78 51 47 3a 2b 19 0e 04 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 0d 08 12 1e 21 45 68 8e 97 c4 e2 e1 d1 c6 be bd b9 c6 d1 da dd d3 d9 e1 f0 ff ff ff f0 ee ee eb e5 eb e1 df de e4 e5 ea ee e9 eb e8 ef e6 e9 ef f4 f3 f2 f1 f4 f6 f5 f5 fd ef fd fc f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f1 f0 e2 df df d0 d3 cf c3 c5 c0 ba ba bb b2 ab b0 ad b1 ab b1 ae b4 b6 b0 b0 b5 b6 be b5 ba be d0 cd d5 cb d9 e5 e9 f0 f2 f9 ff ff fe ff ff ff ff ff ff ff f8 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef eb ed db cd ba b3 ab 99 9b 92 8f 8f 89 7c 66 52 46 28 22 17 05 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0b 1b 29 3e 6a 8e 9c b9 d5 d9 cf c5 bc b6 b8 c4 d3 d8 db d6 e2 ec f9 ff ff ff f0 e7 eb e6 e4 dc db dc db da e6 e9 df d9 e6 e6 e7 e6 e4 e7 ef e9 f2 f3 eb f6 f1 ef f4 f2 f4 fc f5 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ef df e2 d7 d4 c6 cf c3 be b6 af b9 b2 ae af ac ab ab a2 a6 a2 a7 a2 ac ad ac a9 ab a7 ad b3 ad b5 b5 bd ce c6 d3 d5 df e3 ea f4 f2 f7 fa ff fe ff fc ff fa fc f4 f2 fa ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f2 e6 e8 d3 d4 c3 b9 a6 a5 9c 96 8b 8a 8e 8b 82 75 57 40 32 27 18 10 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 07 0c 13 1a 29 45 65 8b 9f c1 d0 d6 d3 c6 bb b2 bf c2 d5 e8 e4 f4 fd fa fe ff ff ff f2 f2 e5 d5 db dd da d7 d5 de df de df e3 e2
 e3 e3 e3 e0 f2 e7 ed ef ed f3 f3 f0 f9 fa f6 fd fb fb fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e8 dc da d4 c9 c5 c4 c4 b5 af ad b0 b0 ae b0 ae a3 a6 ac a7 a7 ac a9 a2 a8 a2 a5 a4 aa 9f a9 a5 ac af b2 bd c5 ba cc cc cd d5 e9 ef eb f2 f8 fc f8 f8 ff ff f5 fb f9 f9 f7 fe ff fb fe fe ff ff ff ff ff ff f3 ed e1 e4 e1 d8 cb be b5 a8 a3 a3 94 90 96 88 91 95 92 80 5f 56 40 2a 21 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 0b 08 09 06 15 21 21 3e 61 89 9d b6 d9 db d0 c7 c0 bd bb cb d9 e3 f0 f3 ff ff ff ff ff ff ff f4 e1 de db dc d6 d3 d4 d6 dc db e0 d6 e6 e6 e2 e0 df e9 e4 ec e4 f2 f0 f4 ed fa f6 fb fd fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 eb db dd ca c8 c4 b9 b7 ae ab b3 b0 ac aa af ac b4 aa a0 a6 aa a8 a9 a9 a2 a0 9f a1 a2 9b a0 a4 a6 ac af aa ad bd b2 bb c6 c4 c8 d5 db e3 eb e0 e9 f0 ec f4 f1 fa f1 eb f4 f3 ee f3 fb f6 f0 fe ff ff ff f7 ea e9 e7 e5 df d2 d1 c2 b6 ac a6 9b 9d 95 8e 85 8b 8f a0 9a 8e 6c 4c 3c 31 1a 10 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0e 0b 16 26 40 6c 88 9f b9 d0 d3 d4 c2 bd be c5 cc d8 ea f8 ff ff ff ff ff ff ff ff f5 e3 e0 e2 d6 d9 d7 d1 d6 d7 e3 de e0 e6 e2 de e5 e8 ec e6 ee f1 f2 ea f3 f5 f5 f8 f7 ff ff fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc e7 d5 d8 cc c1 c2 bf b4 b2 b1 ae b1 a8 a6 aa af ae a9 ab a0 a1 a9 a7 a4 a1 9d a3 a0 a2 9e a0 a0 a1 a7 a6 9f af af a9 ae af be b2 c5 c4 c7 cc d4 e0 e0 e3 ea ec ee ee ea f2 ea e3 e1 e6 e6 f5 ea ed f2 eb f0 ee e9 e3 df d7 cd ce c7 ba ac ae 9d 9a 99 92 8f 85 93 93 9b 9f 96 6f 5b 40 29 1b 11 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 08 07 0a 22 2c 3d 60 8c a1 b6 d4 d6 cb c4 c1 b8 c4 d5 e5 fa f0 ff ff ff ff ff ff ff ff ff f1 e3 de d2 d9 d5 d2 cb c4 dd da e5 eb
 f0 ee eb eb f2 f0 f5 ec f4 f5 f0 ff fc f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f7 df d4 ce c5 bf b6 b4 b3 a9 ad a1 ab b2 ae aa ad b1 a8 a9 a6 9e a8 a2 a0 9d a5 a6 a0 a8 9d a4 a3 a1 9f aa 9e ae a5 aa aa b0 b4 b0 b8 bc bc bb c6 c6 d8 d5 d9 dd e4 ec e8 e5 ea e3 e1 de dc e3 d9 e9 dc db e3 e3 e0 d3 d8 ce d1 c4 ba b0 b3 a5 9c 9c 90 83 84 89 88 92 8a a9 96 80 66 46 3e 22 0f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 06 09 15 24 2a 3f 65 89 a3 b6 d5 cf bc bf c5 be d1 e1 ef f6 ee f3 ff ff ff ff ff ff ff ff f7 ee e3 dc df d6 d0 d8 da de dd e5 d9 e3 ed ea ec fb f2 f5 fb ff ee fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee eb d3 cc c7 b9 ad ad ae b6 af ad a4 a5 a5 a3 a8 a9 a4 a5 ae a0 9d a5 aa ac a2 a5 a1 a4 a2 9f a4 a5 a5 a5 a0 a6 a4 a4 a5 9f ad a9 a9 b6 b0 b8 be b5 c4 be c8 ca d5 dc d2 df d8 da d9 d4 dd e2 df de db da cf d7 d1 d6 d8 c3 c4 c0 b5 b1 a9 aa a2 9d 95 99 81 85 87 84 83 9a a4 a5 7a 5f 52 36 25 1f 0b 06 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 0a 10 1a 25 33 59 83 98 b4 d9 d9 bf c2 c0 d2 dc f1 f5 f7 ef f9 fd ff f7 ff ff ff ff ff f9 ec ea e5 e1 d9 d2 d2 da d9 e5 e6 e2 e8 e3 e7 eb fb fc ff ff ff f9 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 e6 e1 d1 c9 bd c0 ae a4 a8 9f a8 a6 a0 aa a1 a0 a8 a0 a1 a7 a3 9f a2 a9 9e a3 aa a2 a3 a2 a6 99 a0 a5 9e a0 9c a3 9b aa ab a4 b1 aa a4 ae ac b4 b1 b2 b7 ba c2 c6 cb c8 ce d8 d4 d1 d0 ce d1 cd d1 d3 ce d6 cc cd c4 c5 bc c0 b9 b1 ab a4 9f a3 98 9a 8b 88 81 81 87 88 84 8f a5 a3 7a 63 56 30 27 14 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 09 07 10 18 20 38 4e 7d 9c a7 c0 d0 cb ce ce da e7 f3 f7 ef f9 ff ff ff ff ff ff ff ff ff ff e9 eb e6 e9 e0 dd da db e0 df e9 e3
 ea e3 ec f3 f0 f4 f5 fc f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 eb e0 d5 cf c3 b9 b2 b3 ab ab a0 a0 a7 a1 a6 a1 a7 a3 ad 9d b2 a8 a0 a2 9f a6 a6 9c a0 9e 9e ab 9c 9b a0 a0 a2 a6 aa a1 aa a1 a7 ad a9 a9 aa b2 b2 ae ae bb b9 ba c1 c0 bf c6 d0 c7 cf cc cb cb d0 d0 cd cb c8 be c2 bd b9 bc b1 a9 b1 ae a4 a0 a2 93 96 90 8e 8a 87 82 81 87 87 a0 a2 88 69 4d 40 23 1f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 04 06 09 0b 18 2a 36 52 77 98 a2 b4 c7 bd bb c5 ce d9 e3 f2 ff ff ff ff ff ff ff ff ff ff ff ff f7 f0 ec e7 df dc d4 d4 da e3 ea ea e8 e9 ea f5 f8 f1 f5 fb fd fb f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e3 dd d9 c8 c6 bc b4 b6 a7 a6 aa 9e a3 aa a0 a9 a1 a3 a6 99 a6 a4 9f a0 a2 a1 a4 aa 9c a7 9c a3 9e 9e a0 a0 a7 a6 9e ab a6 ac a8 a3 a9 a8 ae ad b8 a9 b4 b8 b4 b3 ba b7 c1 bc bb bd c0 cc c5 cc c4 c4 c3 c3 be bf bb b6 b6 b7 b5 aa b2 a9 a7 a1 a0 97 91 8e 85 81 89 89 8a 86 92 a0 aa 85 73 4b 41 33 13 0f 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0a 13 1e 33 4f 76 97 a3 a2 bc c1 b9 be c6 d0 da e7 fb ff ff ff ff ff ff ff fd ff ff ff fc ea e5 e7 d5 da de de e0 dd df e0 f0 e7 f1 ee fa ed fa fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e8 de db ca be bd b9 b5 b2 b3 b5 a5 aa ae a0 9a 9c 9a a4 a0 a4 9f a2 9a a5 9d a5 9c a4 a2 a1 a0 a2 9c 9d 9c 9d a2 a7 a5 a6 aa a6 a8 aa a3 ac a9 ac aa ab b1 b5 b2 bb b1 c0 b9 b8 c2 c5 bd bf c3 c1 bd bf bf c2 bd b9 b3 af ae b1 af ac a6 a6 9e 9c 96 8a 89 8b 87 85 7a 81 8a 93 a5 a5 7f 6b 48 44 24 18 0e 05 07 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 03 0b 06 12 1e 21 2f 4b 65 8c 9f 9b a1 bd c1 c1 ce d4 dc e8 f3 ff ff ff ff ff ff fc f1 f0 ea ee f4 eb ee e4 e1 da e3 df dd e6 e6 e1
 e5 e7 ef f2 ee fe f4 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f7 fe ff fd ff ff fa f9 ff fe fc f8 f7 fb fd fc fa fe fc f9 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd e2 d8 cc c4 c6 be bc b9 bc b3 ad b4 b4 b3 ac a6 9c a1 9f 92 9c a0 9c 9c a0 9c a5 9d a0 9c 9b 9e a5 9f a0 9a 9f a5 a1 a3 a1 aa aa a5 ac a9 a5 a6 a9 ab aa af ac af ad b1 b2 b3 b6 c0 c0 bb b7 c2 b7 bc b1 af b3 ad b2 ab ab aa af ad aa 9d 9f 98 95 96 90 8d 8b 88 8a 8b 84 8c 91 a9 99 86 6a 54 3f 27 10 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 08 06 0a 18 1f 35 41 6a 80 95 9e 9a b3 be c0 ca d1 dc e4 ed f2 ff ff ff ff ff f5 e8 e7 e4 e7 e2 e6 e1 e4 e0 df e2 e3 e4 e7 eb e6 e7 e7 f5 ed fc f6 f9 fe ff fd ff ff ff ff ff ff ff ff f6 f5 ed f1 f3 fb f3 f8 fd ff ff fd f7 f9 f5 ed f6 f5 f8 fa e7 f7 f6 f3 f3 f6 f4 f4 ee f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e1 d9 cd d1 c5 c2 ce be bd b6 ba ad bb c0 c0 b0 9f 9f 9e 98 9f 9b 9a 9f 9f 9c a6 9c a1 a2 a7 a1 a3 a4 a0 97 a4 9a a3 a8 9c ae a2 a2 ab a9 a6 a6 ab a7 ac b0 a7 b1 a9 a9 b1 b5 b4 ba af b7 b3 bc b0 b6 b3 b6 b2 b2 ae af a5 a7 ae a3 ac a4 a4 96 87 95 90 94 8e 8c 8a 86 82 8c 90 a2 a2 85 66 57 46 29 16 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 07 00 07 11 19 19 29 42 58 73 92 99 8f a7 bf c8 d4 d2 d6 d8 e2 ef ea ea f6 ff ff ec d9 d2 d2 df dc de e6 de df da e1 e5 dc e1 eb ed f2 ec f2 f8 fc f8 ff fd fc ff f7 fc ff fe fd f8 f8 f8 f1 ec e5 ea e9 f4 fb fc ff ff ff f8 f5 f5 f8 eb eb ed ec ef e6 e4 e5 e9 e9 eb e2 e7 eb ef fb fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc e5 dd d6 ca cf c9 ca c6 b9 b7 b3 ae b1 b3 c1 bb aa a3 9b 9b 97 99 a7 9b 9f 9f a5 98 9b 9c a0 9b 9d 9a a2 a5 a2 a1 9c 9b a5 af 9e a6 a7 a4 a5 a9 a8 a6 ac a6 ad ad aa ac ac b6 ae b9 b3 ad ab a9 aa b1 a9 ab ac a3 af a4 a6 ae ae ae ab 9b a3 a1 94 93 8e 8e 8d 8d 8e 85 85 79 9d a6 9b 86 6f 51 3b 2c 17 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 09 14 1f 25 3d 52 77 91 91 90 91 b2 c1 c8 d1 d8 de e0 df e2 e6 e3 e3 fa ed d3 d4 d5 cd dd d5 e1 de db df dc e4 e7 e5 e4 ee
 ec eb f2 f0 f7 f9 f5 f9 fa f2 f5 f6 f5 f6 f1 eb ea e3 ec e3 e2 e8 eb ed f7 ff f5 f1 f5 f1 e5 e5 e5 df e6 e0 e0 e1 e3 dc e1 e0 e5 e5 e3 df e5 f0 ea f3 fb ff ff ff ff ff ff ff ff ff ff fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb de d7 dc d4 d8 d8 d1 c6 bd c0 b6 b5 ac b0 b1 bb b6 a0 9b 8e 93 96 97 a0 9a 9a a0 9b 95 97 9f 94 9f 97 9f 9d a2 a6 a3 a5 9a a6 9f a1 a8 9d a6 a5 a4 a9 a6 a1 aa a8 ab aa a9 b2 a6 aa b0 af aa ac ae af a6 a5 a5 a3 a9 b2 a9 b3 b0 a9 a5 a7 9e 96 90 92 8b 89 8b 8a 7d 7e 7f 7d 91 a5 9b 84 6a 4c 37 22 1a 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 09 18 15 26 3c 51 6f 8d 96 8d 8d a0 bc c1 cb d7 e3 e0 e3 de dc eb ea ec e6 db d6 d7 dc dc dc e1 d5 df df e5 e6 e6 e1 eb e9 ed f0 ea f3 f5 ef f3 f4 f3 f0 f2 ef ef e8 e6 eb e7 e2 e7 e4 de e6 ed ed f7 eb f4 e9 ee e8 e0 df e3 de df e3 d8 df e0 dc e9 df e1 e1 e1 e2 de e7 ed e9 f0 fa ff ff ff ff ff ff ff ff fd f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e1 db df df e6 de d7 d6 c9 bf c0 ba b2 ac b3 b1 ab a2 a5 9a 94 96 9d a1 97 94 a2 9a 9e 9c 9f a4 a0 97 9c a0 a3 9d a0 a1 9e 9c a7 a5 a7 a3 a4 9e a0 ad a9 a1 af a7 a5 a6 a5 ae a8 ad af b0 aa b0 a6 af a9 ad b0 a9 b0 a6 ab a7 ae ab a7 a8 a2 9a 96 92 93 89 8c 88 7e 79 7a 7f 91 a1 99 7f 68 54 46 22 1b 0d 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 03 06 0d 12 1b 29 34 4d 6f 85 a0 8a 86 95 a5 b7 c7 d2 d3 e2 df d9 e0 eb ef e3 df d3 d0 d8 d3 dc dd d7 da e1 e0 e1 e9 df e2 e3 e4 ec ee ea ec ec ef ed e6 e7 ea e6 e8 e3 e9 e0 e5 df d5 e0 de d7 da e0 e2 ef ee e8 e7 e3 dc df da da e1 db e0 d1 dc e2 d8 df e4 e4 e4 e5 e4 ed ec ee ee f8 fc fe ff ff ff ff ff ff ff fd fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 e5 e3 db e2 e6 e1 da df c9 c6 c5 b5 b6 af b1 b3 b3 ad 9e 9d 9d 92 92 8f 97 93 9a 98 95 9b 97 9f a1 9f a0 a2 a4 a2 9f 9d a3 a8 a3 a2 a5 a3 a5 a9 a0 a9 9f a0 a5 a5 a2 aa a7 ad a9 ac b8 a8 a6 aa ad b0 a6 a9 ae ac ae b0 ae ae aa a8 a6 a5 a0 a3 a3 91 94 92 8c 8b 86 71 75 80 93 a0 99 7f 69 4e 36 28 14 07 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 09 1c 22 36 52 65 87 90 90 85 7f 8a a4 bc bb cb cd ce cf d1 f1 f6 ec db cf d1 d7 d5 df d9 d8 e1 e1 dc e0 e2 e1 e1 e4 e4
 ee e5 ea e3 e1 e7 e4 e7 e8 e5 e7 e2 e6 dc de e0 d8 da db d5 d5 db d9 de dd e1 e6 dd d3 dd db d7 d7 dd dd d9 da db de dc e2 d6 d9 e1 de e1 e1 ea e7 f0 f7 fb fe fb ff f6 ff ff f4 fc f3 fb ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef e4 e1 e3 e6 e4 e0 de e2 da cf c4 be b0 af a8 a4 a7 ae a1 9b 9c 98 92 92 96 9a 93 9a 97 99 9d 9d 9a 9b 99 a0 a3 9f 9c a6 a5 a1 9e a1 a1 99 a0 9f 9b ac a3 9b a3 a2 a3 a1 a7 b0 a7 a9 ac a5 ab a6 aa b2 af ae ad a3 aa b0 a8 b0 aa ac ae a2 a8 98 9a 99 95 8f 7f 87 80 74 6b 7e 90 9e 8f 78 65 53 43 2f 19 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 06 0e 14 2f 39 4c 61 80 8f 93 89 7e 8b 9d aa b0 bb c0 bd ca ce e9 f2 e1 d7 cb cb d1 cc d8 d9 d6 d9 e2 db df e8 df e6 ed e4 e5 e3 e7 e4 e0 e1 e3 e4 e1 da de de d8 d9 d3 d8 e0 d5 d7 d4 d0 d5 d6 d4 d7 d6 d6 db df da d6 d3 dd e1 d8 de d6 d4 d9 d4 dc d9 d6 e1 dd e2 e4 e2 eb f6 f8 fd f3 f4 f5 f8 f2 f4 f5 ee f5 f4 e9 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 e8 e2 da da e3 fa f5 e3 e8 e5 e8 ea e6 ed e1 d9 d0 cb be bf b5 b4 af aa b0 a9 a1 9d 97 9e 92 96 93 97 8d 9e a1 9b 9d 9c 94 99 9d 9b a4 97 93 a5 a5 9d a8 9d a0 9b a4 a8 9f a3 a1 9a a3 a4 a4 a5 ac 9f a6 ae a4 aa ad a6 ac a5 ad ae ac ad ab ad af ac a9 ad a5 a0 a2 95 99 8f 86 8d 7b 76 71 77 83 8f a3 92 79 69 56 3d 32 16 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 03 00 06 05 0f 16 2c 35 4b 5f 76 90 8d 85 82 7d 90 9b a5 ad b9 bc c2 c6 dd e0 d8 ce cd cf d4 d9 d9 df d0 d3 d3 d8 de e3 e4 e2 e3 e2 e9 e0 e1 dd dd da dc da dc db d6 d6 d4 da d6 d0 d1 cb d1 d1 ce ce d1 ce c9 d0 d6 c6 d1 d7 cd e0 df da d7 e0 d8 db db d7 e0 db e3 de da df de ed e7 e5 f1 f1 f7 f9 f1 e4 ee e7 e9 e3 e3 e3 e2 e4 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 e0 d0 cf c5 c1 b8 bc bb c3 c3 de e6 e3 e6 eb ee f3 ea e1 e5 d4 cf d1 c4 b9 b2 b1 b0 a5 a8 a2 a0 a6 9f a0 a2 a3 8f 9e 8d 89 91 95 95 9d 9a 9e 9d 9c 9c 9d 9f 9d a4 9c 9f a0 a2 a0 a4 a1 a1 a3 a0 a4 a2 9e a6 a3 ab af ad b7 a9 a3 a9 b0 a8 b2 ad ae ab b2 ad b4 ab af ab b0 a4 a4 9f 8d 92 91 84 85 84 74 70 73 7b 8e 9d 91 78 6c 52 3c 20 16 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 06 05 12 14 24 34 4a 60 6c 86 8c 7b 7f 75 83 8d 99 a7 b0 b3 bb c4 ca d2 cf ca ce d2 cc d1 d4 d8 d8 d6 d6 df df de d9 d8 de d2
 df dc d3 d6 d6 d7 d7 d4 d1 d4 cf c8 ca ce cb c9 d3 cf c8 c5 cd c9 cf cd d5 d2 ca ce cd cd cf cf ce cd d5 df dc d9 dd d5 d3 d7 d8 e6 de d6 e1 e5 e7 ef f6 f1 ee ef ec e4 e2 e2 dc de d5 d8 da df ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef f4 ff ff ff ff cf ac 9a 97 99 86 85 83 8c 94 9a 97 ac c0 df df e1 e2 ec ea e6 e2 df de d2 c7 bc b1 b3 a5 ae a3 9f a8 a2 99 9d 9d 99 9b 9a 99 95 8c 8f 94 91 95 99 9a 92 97 94 97 a5 9a a0 98 98 9f 9e 9f a5 9b a1 a0 a2 a5 a5 a2 a8 a7 a6 ab a2 a5 a6 a5 ad 99 a5 a3 ac ac a8 ad ae a6 aa af b1 ab a6 9b 9a 94 93 91 8a 7d 70 6d 6f 6b 7a 8e 99 8e 71 5f 50 2f 23 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0b 0c 20 1f 35 46 5f 73 89 89 79 76 7e 7d 8b 95 9f a8 af b9 bf c1 cf ca c6 c3 ce c8 d0 ca d1 d2 d4 da da db db d7 db e5 dc d8 d3 d1 cc d2 cd c8 cb cc c6 c4 cf c7 c6 ca cc cd d0 be c9 bc c5 cb c7 d0 ce c6 c9 d1 d0 d3 d1 da d1 d8 d6 db d5 da d7 d5 d6 da d5 e1 e4 db e5 e2 e0 f0 ed ec ed ee e3 dd db d6 d0 cf d2 d7 d6 da ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff d2 a9 9a a3 a8 9e 8c 84 76 76 69 64 67 69 65 6c 68 74 7f 92 b1 d1 d5 dc ea e5 eb e9 e1 eb d9 d5 cb c4 ba af ab a2 a8 a6 a2 a4 9d 9a 9f 97 93 91 a1 98 96 8c 8d 8b 8d 96 9a 94 9d 97 93 94 94 9d 95 95 99 9c 99 98 96 a3 a0 a3 ab a9 b6 ab b3 ac a7 aa a6 a6 a9 a9 a8 af 9f a7 a7 a5 ad a8 af b1 ab a7 a8 aa 9e 92 96 8b 88 83 7a 6c 70 6d 75 74 8b 93 91 70 64 4d 36 24 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0b 10 11 29 31 46 5f 75 86 80 7c 79 71 77 85 86 9a a5 af b3 af b5 c1 c2 c7 ce cb ce cc ce cf dc d8 d8 d9 df dc d1 de d6 ce cc cb d0 cb ca c7 cb d0 c7 c5 c9 c4 c4 c4 c7 c2 c4 c9 c7 ca c5 c7 cc c7 cb c5 cd cc d2 ce d0 d6 ce d9 d4 d4 d9 cf ce d5 df d9 da e2 e2 e1 e2 df e9 e4 e8 ef f0 eb e5 dd e1 d4 ce ca c4 cc cd d0 db ee ff ff ff ff ff ff ff ff ff ff ff f9 dd c0 a3 8f 7a 70 6e 6e 66 5e 5f 57 56 53 4f 4a 55 60 60 5a 61 67 82 9d c9 d4 d7 e6 e4 e1 e3 e2 e6 dc d3 d0 c4 b7 b3 ae a5 a3 9f a2 9d a0 99 96 94 96 9b 98 98 8f 94 8b 91 96 90 99 93 93 9c 95 8d 9a 9c 95 91 9e 9a 99 93 94 98 a0 a6 a7 ad af b0 af ab af b1 ae a0 af a4 a4 a4 a9 ab a7 af a4 a8 ac ae a4 a9 a1 96 97 96 8d 8a 80 84 79 73 70 71 70 76 8b 99 91 75 5f 4d 37 2d 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 15 1b 1e 33 44 61 6d 82 8b 7e 76 73 7b 75 80 84 96 a4 ac ab b5 b5 bb c5 c7 c1 ca cb c3 c5 d3 ce d2 d3 d6 d6 d6 d0 d4 ce
 d4 cb c6 c6 c5 c2 bc c4 c1 c7 c5 cb bf c5 be c4 c4 be be c4 c7 c1 c6 cb c9 c2 ca cf cd cf d5 c9 d1 d0 cc d8 d4 cf ce d4 d1 d3 d9 d5 d3 d7 dc dc df e5 e1 e7 e8 e9 e5 db d5 cc cf d0 ca c8 c2 c2 c5 dc ff ff ff ff ff ff ff ff ff e1 b1 9e 7c 6d 64 61 54 59 55 49 4b 4e 47 47 4a 3a 47 48 48 4a 46 4b 53 62 71 92 be c6 d4 da df e3 dc ea e3 dc d2 cb bb bd b5 b1 a7 a2 a2 98 98 a2 97 98 95 8c 9a 9b 9b 8b 90 9b 8b 98 85 8f 90 92 8f 96 93 95 95 91 92 93 9b 9b 95 9a a0 a2 a8 a7 aa ae ab ad a9 a4 a9 a3 a0 a1 a8 a9 9f a1 a4 a2 a7 9e a6 a1 a3 9d a0 a1 94 96 87 8d 87 86 79 76 70 6e 6b 6b 73 87 8e 8e 73 5f 4a 34 20 0b 15 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 11 0f 26 36 3f 5d 68 7c 8a 76 77 78 78 80 82 85 93 99 a1 ac ac ae b6 b9 c0 c4 c2 c7 cd c9 cd c9 ca c7 cc d8 c6 cb cd c4 c9 c1 c1 c1 c1 be c5 c7 c4 bd c2 bc c4 ba c0 c4 bf be bd c1 c9 c3 c4 bb c9 cb c0 ca c5 c8 c5 cf d1 cf d0 d2 d1 ca c8 d3 d5 d1 d6 dc d3 d9 d9 d9 dc e0 dd e8 e2 df e1 d5 d4 c7 d1 cb c5 c0 c4 ba c5 cb e7 ff ff ff ff ff ff e0 b5 8f 71 69 56 51 4f 46 47 48 44 43 3f 3f 35 37 32 35 33 36 3a 33 45 46 4b 52 69 86 ad c9 d5 d3 d9 e2 d9 de e2 dd d8 cd c2 b5 b8 b0 a3 a6 9c a2 96 9c 93 95 92 98 99 8f 8d 93 8e 95 90 97 93 8f 96 92 88 8c 92 97 96 8f 99 88 93 95 92 97 97 a6 a5 aa ac ad ab a4 a6 9b a5 a6 a9 aa ad a5 9c ab 98 a5 99 a0 a4 a0 a7 9a 98 96 95 92 8b 84 81 71 76 74 6d 6c 70 72 6b 7c 8c 84 6d 5f 45 31 20 16 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 00 07 07 0c 1b 21 2e 46 55 69 80 8a 7c 7c 79 78 78 7d 78 89 94 9d a5 a9 ad b2 b8 b5 ba be c5 c6 be c3 c2 c4 c0 bd c7 bd bb c0 c1 c0 bb c3 c2 b8 bb b9 c4 ca be bd bb ba b2 bf c2 c6 be bd c2 c1 bb c2 c6 c3 c7 c9 c5 c9 cc c9 cb cf ce cf d1 d4 cb d2 d0 d3 d4 db ca d6 d0 d3 d9 da dd dd e1 dd e2 e1 d6 d3 c7 c7 c4 c0 be b7 bc c3 c3 d3 ff ff ff ff dc af 93 77 61 52 46 43 44 46 45 3b 3a 3c 3b 36 3d 34 30 2e 34 2f 34 38 42 38 3d 39 4f 5f 86 b2 cb d0 d4 d1 d9 d3 d7 e3 d8 d0 cd c1 c8 b3 ad a9 9b 9c 9a 9f 9b 9b 98 95 93 93 91 8e 94 90 86 86 88 8c 89 8b 90 81 88 8a 89 95 89 88 91 94 90 91 9b 9a 99 a2 a5 a2 ac aa a5 a5 9e a7 a2 a3 a5 9a 9e a0 9b a1 a5 97 a6 99 98 9c 9f 9d 95 89 90 8b 86 83 73 75 74 71 6d 6f 6f 78 7d 8a 84 67 64 46 33 25 0f 13 06 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 0e 19 1c 3d 47 55 6a 77 80 7b 79 78 79 7c 7d 80 86 8b 8e 99 a3 af b3 b5 bd b9 b9 be be c4 c1 bc bc c1 b8 be b6 b9 b7 be
 b9 b1 b7 b6 b4 be be b9 be ba be b9 bc ba b7 b9 b6 b4 c3 c2 be ba bb bd c5 c5 ca c3 c9 c7 ba c8 cd cd c5 d0 c5 cc c8 cf db d0 d5 cf d3 c6 d7 d6 d9 db e2 db dc d9 d5 d7 cc c9 bd bd bc bb ba b6 ba b7 b9 e2 f8 e0 c5 9d 75 5f 49 44 41 3d 3b 3c 34 3e 3a 29 35 27 29 26 2a 2c 21 24 24 2d 27 39 33 2d 32 40 5e 79 ad c1 c8 cd d1 d2 ce dc d5 d4 cc d7 c6 be be b0 a4 a1 9d 90 92 96 93 92 8f 97 95 91 8b 8d 8b 8c 85 8b 88 89 87 8d 8d 8e 8e 8e 8a 8e 95 8b 86 92 90 99 9e 9c 99 a5 98 a5 a1 a5 ad a2 9d 9a 9a 9f 99 94 9a 99 9b 99 9b 96 9a 94 94 90 97 8d 92 8b 85 7c 7f 75 70 75 6f 6c 69 64 6c 7a 8a 84 69 5b 47 31 16 14 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 16 1f 34 41 4f 6d 77 7e 7c 73 73 75 78 76 77 83 86 83 91 9a 9f aa b2 b7 b5 be ba b5 bd ba b8 b6 af ac b2 b9 a9 b2 b5 b3 af b5 b5 b1 b5 bd b3 b7 b1 bc ba b3 bb ba b9 ba b9 bd bf bf bb be c2 c6 b6 c1 c4 c4 bb c1 c9 c1 c6 c6 d2 cd cc c8 ce cc c2 c8 c6 d5 ca ce c9 d7 d6 d5 d5 cf d1 ce cb c5 c2 bd c1 b6 c0 b9 b4 ae b0 b5 bc cd ac 92 73 55 44 46 38 37 30 34 2f 2f 2f 2c 29 28 25 25 22 1f 21 22 21 25 1f 25 26 2d 27 2d 36 50 80 aa c5 ce d0 d0 d6 cf d4 d4 da d3 d5 ca bd b3 a6 ad 9d 9b 98 93 95 9a 8c 91 8c 8b 8e 8e 8e 8a 84 84 7d 7e 87 7f 8c 8f 93 8f 92 8e 86 89 8f 8a 8c 92 95 8e 92 9e 9a a1 9b 9e a3 a4 9b a1 9d 95 93 94 91 93 91 92 8e 93 95 91 8f 8d 92 8e 93 8f 85 78 79 77 70 71 6a 5f 63 63 6d 68 69 83 78 6a 5b 39 2b 21 07 0d 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 01 06 0a 05 16 28 2a 44 51 64 7b 78 74 6a 71 73 78 76 7a 73 85 85 8b 97 9d a2 ab b5 b6 b7 bc bd b5 b5 b6 b8 b3 ab aa af ae b6 b8 b3 b2 ad b4 b7 b3 ab b8 b4 b7 b9 ba b6 b7 b6 b8 be bc b0 b8 ba bf be bd c1 bf ba c0 bf b6 c3 c8 c5 c7 ca cf cc c2 cb cb d3 cc cb c1 cd d1 c7 cc d0 c9 d0 d0 ce cb c6 ce ba c0 b7 b1 b1 b7 b0 b0 b6 b4 b2 b5 b6 90 7a 67 51 33 30 2a 2b 29 2f 32 29 27 2d 27 27 26 25 19 1d 20 20 21 16 14 1d 29 2b 2b 33 2c 44 69 a5 c0 ca ce cf d4 cf d8 d5 d9 cd cb ce c0 ad a8 a4 a0 99 93 8f 9b 84 8b 92 92 8d 88 8e 84 83 85 82 84 7d 80 79 82 89 86 91 8c 88 8c 8e 8a 93 87 8b 95 9c 99 9b 9f 9b 9f 9d 9e a4 9b 9b 8e 98 92 9a 9b 8d 92 8b 93 8d 94 92 94 92 94 7d 8d 81 7d 80 76 72 71 6e 6b 69 60 5f 63 61 69 7b 7f 6c 5d 3d 2b 23 19 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 0a 0d 11 1d 33 47 5c 65 76 7b 77 6e 69 69 74 73 7e 80 80 84 89 8d 97 98 a5 b0 b0 ba b4 b8 b4 ac b4 b5 aa ae b6 ae af ad b3
 b2 b1 b4 b0 b4 ae ae b3 b8 ba b8 b5 b7 b5 b4 b4 b4 b6 b6 bb bb b9 bf b9 b8 c0 b9 b7 bc b7 bc c0 c4 cb c7 c9 c0 c6 c9 c1 d0 c9 cb ca c4 c4 c4 b9 c7 bc c8 d1 c9 c7 c7 be bf bf b6 b5 b3 ac ab aa a9 ae b8 ab b0 8c 6b 61 3f 31 32 29 2d 24 22 2b 1e 1f 1e 1f 1d 27 24 21 18 18 14 19 22 21 1f 27 23 24 25 2c 39 5f a5 bb cb cf cc cb d4 d1 d9 d3 d0 cf bf be b7 a9 ae 9e 9a 92 91 92 8c 8e 87 91 82 8b 85 86 86 86 82 82 82 82 7a 74 7d 7b 94 99 93 8a 8e 8a 90 89 97 8e 95 94 9b 98 a1 a3 95 a1 96 92 97 91 8c 92 8c 8c 8d 95 8e 8a 8c 93 92 92 92 99 90 92 80 80 77 75 75 69 6d 6c 68 6b 62 5e 62 61 71 7a 67 58 44 3c 23 12 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 10 14 2b 31 42 4a 63 6e 73 79 6e 6b 6d 66 6f 72 7f 7d 81 8e 85 89 93 97 a6 a6 a7 b3 b1 ae b6 b0 b1 a7 a0 a9 a5 ab ac ad a6 a5 a6 aa ad ad af ad a4 aa aa b4 a7 af b7 b1 b5 b4 b1 b5 b4 b4 b6 b9 bb b4 bd b9 bb bc be bd cd bd bf bf c0 bf c4 ca c6 d0 c6 c4 c0 c6 b5 bd bf c0 b7 c1 bd c4 b6 c1 ba b2 b1 b5 aa ba aa ad af a8 ac ab a1 85 6b 5d 38 29 29 1e 1a 20 1a 1e 19 13 1e 20 1a 18 12 1a 15 1c 11 0f 19 11 16 10 1c 21 22 2d 34 50 9b b9 c4 ca cf d4 d7 d0 d5 d4 cc ca c6 c2 b1 ae a0 9b 98 91 8f 8f 86 89 8b 88 8b 8a 81 84 82 85 87 77 7d 79 81 7d 76 76 89 92 92 92 90 92 86 89 87 97 9c 98 95 8d 93 98 95 96 92 90 96 88 8b 83 8f 8e 8c 90 8a 92 8c 86 8f 89 8f 94 90 8c 85 7c 77 75 6c 62 6b 61 66 5b 63 5b 62 5b 6a 6c 66 61 45 39 20 14 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 06 11 19 1c 2c 3b 55 63 79 77 7a 73 6c 62 68 70 77 79 86 7d 82 80 8d 8c 9b 9a a6 a8 b0 af ab ac a7 b1 ab a1 ab a5 ac a9 a5 b1 ab a3 a9 a9 aa ad ae ad b2 a9 af ac ad b2 af b9 b3 a9 b6 b1 ae b6 b3 b8 b4 b0 bb ba bd be be c1 b7 c0 c2 c5 bf c5 c3 c4 cc ba bc b8 b1 bb b7 b4 bc b7 bc b7 b7 b5 b3 b1 b1 b5 a5 a6 a8 a5 a5 aa aa a6 a9 a3 8b 6f 64 32 23 21 17 21 1f 20 17 15 0e 19 1b 14 14 17 0e 15 15 19 15 0f 15 19 14 1a 21 1a 2a 29 49 95 b1 c9 d1 cd d5 d0 d5 d6 d5 d2 c6 c3 b6 b2 a7 a8 a3 98 99 8b 83 93 83 89 8b 8c 8f 7f 84 89 7f 7e 7f 81 81 7d 7e 78 7c 86 95 a5 97 94 96 88 8f 96 9d 9c a2 9a 95 90 8f 92 8d 8b 87 8a 8f 8a 89 8b 8d 88 89 8c 8b 91 8f 95 8d 90 8a 89 88 7e 76 71 6d 6a 67 65 68 66 5f 64 5b 57 56 64 6c 68 5a 45 37 25 1c 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0a 17 20 33 3c 59 5b 6c 7f 71 67 64 60 6e 6a 72 76 7b 87 80 7e 89 92 90 9f 9d a3 ac a5 a7 ab ac ae a3 ac ac a1 ab ae a5
 af a9 a9 a7 ac a6 aa a9 a6 b2 a7 a9 ae b4 af b4 ac b2 aa b0 ae b1 b4 b4 b6 ae af b7 b2 af b8 c0 b4 bd bb bf c2 c1 bd c0 c8 b7 c0 b9 b3 b5 ab ad b3 b6 ab ae b4 ad ab b3 aa a6 ab a0 a4 a9 a6 ae a6 a9 ad a4 95 8f 78 55 35 23 16 13 11 1e 1f 16 10 00 0e 15 19 0e 13 10 0c 0c 09 15 0f 15 17 17 1c 13 18 26 2c 48 90 bd c2 c8 ca cd d3 d8 d9 d4 c9 d1 c1 c0 b9 af a4 a7 97 9c 92 8c 88 8b 85 8a 8b 86 83 7f 88 84 7f 7b 7e 7e 7f 7d 79 80 85 93 9b 8f 97 99 8c 95 9b 9c a7 a1 8e 94 91 8e 8f 8d 8f 8d 89 89 85 82 8e 84 83 84 89 97 8d 89 90 93 94 8d 82 80 78 6d 67 6f 6a 62 66 5f 5c 5d 59 58 5b 5d 61 66 6d 5e 4d 33 2d 0e 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0e 17 24 30 42 48 62 6a 7b 6d 68 65 5d 67 66 6c 79 78 85 80 81 82 85 94 97 96 9f 9c a0 a2 a1 a5 a1 a5 a5 a1 a5 9c a6 a0 a8 a8 ae a5 a2 a3 aa a5 af b0 a6 ac b1 aa ae ae a7 ac a9 a9 a2 ac ae b1 af ad ad ad aa ad b7 b4 bb b9 b5 c0 bc bb bd b9 b9 be b4 b5 ae af ac ae ad aa a5 aa a4 a5 ac a9 aa 99 a7 a4 a3 a5 9e a0 a0 a8 a0 a6 98 8a 74 47 2f 19 0b 12 16 11 10 14 12 0d 13 0e 08 07 0b 0e 0f 13 0b 0c 10 16 0c 15 18 13 1c 1c 20 3d 83 b8 c4 cf c6 d2 ca d9 dd d9 cd c9 c0 bc b5 b0 9e 9a 9d 91 8e 8f 84 83 86 7f 83 86 7f 86 8b 83 80 7f 7a 78 7d 7d 81 7f 85 8c 8c 93 8b 91 99 9d 9a a2 9b 9d 95 8f 84 81 7e 92 87 8a 8c 83 84 83 84 86 8a 8d 8c 92 86 8b 90 88 91 83 7d 84 6c 6e 6e 64 62 62 5d 5d 62 58 66 58 5b 5b 5d 71 60 5b 52 3b 22 15 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0b 17 21 2a 3d 54 62 6e 72 71 60 5a 62 5f 6a 66 74 75 7d 83 84 82 86 86 90 92 94 9b 94 9d 9e a5 ac ab ae ab a3 a2 a3 a5 a5 a0 a2 a8 a3 ac a7 a8 a2 a0 a7 a5 a8 ab a8 a4 a6 a6 b0 b1 a8 a9 af a5 b8 ab b0 b0 b2 af aa b3 af b4 bb b6 bc b7 b6 ba b9 b6 b8 b2 af a6 a8 a9 a6 9d a2 a4 a2 a0 a0 99 9c a5 9e a1 98 9f a6 a3 97 a2 9e 98 92 8d 75 4b 23 12 0d 14 15 14 14 16 15 12 15 10 15 0c 0a 0e 11 0f 06 14 0f 14 15 11 0d 0f 15 20 25 3b 7a b6 c6 ce c9 d1 d4 d7 d3 cd d3 cd c1 b9 b2 af a5 a6 99 90 83 8b 90 81 85 87 81 80 78 82 79 84 82 82 80 7b 7e 83 84 79 7f 88 86 84 8c 88 86 94 a6 99 a5 a4 95 8a 82 87 91 82 84 80 80 83 84 86 89 88 7f 88 8e 94 97 90 9a 86 8a 7e 7e 74 6a 6d 6a 6f 67 66 56 57 58 60 5d 57 57 51 61 64 64 62 4a 41 2e 1d 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 0b 11 20 33 3d 50 62 6e 6b 77 65 5e 5d 5f 6a 65 69 77 77 7d 7f 85 8a 92 92 8c 94 94 92 96 98 9d 9f a5 ae a7 ae 9e a3 a8
 a5 a3 a6 a6 ac 9b a7 a0 a5 a2 a6 a5 a1 aa 9c a7 a3 a5 b1 a4 a8 b0 af a5 ac ab a8 a7 ad b5 ab b5 b1 af b2 bb b4 b7 bb b9 bb b2 b5 a9 a8 a6 a6 a4 a5 97 9e 9b 9b a1 9d a5 a2 9e a0 9f 92 97 a0 a2 9b a0 a0 8d 8f 89 75 46 21 10 11 12 12 0f 07 14 14 0f 0e 13 0c 0d 0f 0e 0c 07 06 12 15 07 17 15 10 14 0d 1a 1d 2a 74 ba c5 cc cd d3 d4 d3 d7 d4 d0 ce bd b6 ba b4 a7 a1 95 94 8c 8d 8b 89 85 84 89 7d 86 80 81 80 84 83 80 83 83 82 81 82 85 8a 88 8e 89 8d 88 8b 9c 97 a0 9a 8c 8d 86 90 8d 8d 8c 85 85 84 85 80 86 8b 7d 92 8c 94 97 97 89 89 7f 80 74 70 6a 6c 60 5d 5d 60 5b 5b 5a 56 60 52 54 51 55 5f 68 5f 58 46 35 1e 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0f 1b 2a 37 4a 5e 63 6b 71 5d 56 53 56 5e 64 66 69 6d 6e 6d 74 83 8c 98 8c 8d 89 8d 8e 8f 93 97 95 a5 a4 9b a8 a0 a2 a4 a4 a9 a2 9f a1 9e a3 ac a0 a8 a4 a1 9e 9c a6 9f a2 a0 a2 9f a7 a9 a2 a5 a0 a9 a6 b2 a7 a5 aa b1 af b2 af b6 a7 a6 b3 ae ab b0 ab a7 9e a5 a2 9a 99 95 9a 8e 9c 92 8c 95 92 96 91 9b 9c a0 9d a4 a5 99 91 88 83 68 42 27 17 12 0f 07 10 12 0b 0f 0d 09 0f 0f 07 09 0b 0a 03 0b 09 08 11 08 14 11 0f 11 17 17 2f 7c b8 c5 cf cf cf cd cf d0 ce c5 cc c3 ba b6 a7 a7 a3 9d 91 8b 8b 87 84 85 85 88 84 85 79 7e 86 85 83 79 81 81 79 7a 86 7d 84 85 81 7e 88 7e 84 8e 90 95 95 92 8d 8b 84 90 82 88 86 82 81 83 87 85 7c 87 87 95 98 8c 92 7d 84 7c 72 79 67 62 63 63 64 5e 5d 60 60 5e 58 55 5c 56 56 52 5b 61 5d 54 43 32 1b 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 14 24 2d 40 4d 62 6d 6e 74 60 56 56 59 62 60 64 69 65 79 70 75 7f 84 88 84 90 8f 8e 8f 93 94 94 93 9d 9e 9f a4 a5 a0 a3 a3 a2 9b a7 a4 9e 9f a2 a1 a4 a0 9b 9f 9b a1 9c 9e a1 a0 9e a1 a9 a8 a2 9f a4 a7 9e a2 a8 b2 b2 af b0 b0 ac ae a6 b3 ab aa a3 a6 9b 9f a0 9f a2 92 92 97 93 90 8d 98 93 95 98 99 98 96 99 96 9a 97 8e 93 89 84 74 4c 28 15 0b 0a 07 0e 0e 13 0d 0a 0b 09 0d 04 0e 09 05 0c 06 05 07 11 0a 0b 18 12 13 14 1c 2e 71 b6 c6 d1 cf d4 ca d6 d2 ce c8 c7 c1 c4 b2 af a1 a0 97 93 8d 8a 89 84 86 85 7c 80 7f 79 7e 7e 81 87 7d 7e 89 83 86 85 8a 8b 8d 7d 81 88 7e 7c 8a 8c 95 90 89 8d 81 8a 83 89 86 82 89 84 81 82 85 84 88 86 8b 90 8d 8a 81 7a 7d 72 6f 65 63 60 5e 5c 5e 62 5c 61 59 54 5b 5b 59 4f 5a 54 55 60 51 4c 33 21 15 0f 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0a 0c 19 17 24 45 4d 56 6b 74 6a 69 53 53 58 5e 5e 66 68 65 69 71 74 7e 84 85 83 8e 8c 8a 85 92 91 90 90 93 9b 9a 99 a2 a3
 a1 a2 a1 9f a6 9b a1 a7 a0 a6 a2 9c a0 a2 a5 a4 9f 9a a2 a1 a1 9b 9b a0 a0 9e a6 a2 9a a7 a0 aa ab a2 a9 ab a4 a6 a5 a5 a5 a3 9e a2 a3 9b 95 97 98 98 94 91 90 8b 8f 8a 92 93 95 98 95 9d 97 9b 9c 91 92 8f 8f 85 6d 4d 29 13 0b 0c 08 0e 14 05 04 0b 0b 0b 0f 07 0a 05 0c 0c 08 05 04 09 06 09 10 14 17 14 1f 2c 64 b0 bf ca cd d8 c9 d4 d4 c6 d0 c8 c6 ba b9 af a4 a2 95 8b 8b 8c 82 84 7e 7c 76 7d 81 79 74 7d 81 8a 83 82 80 84 84 84 8b 86 8d 7d 7e 80 78 86 7e 83 8a 90 92 8c 8a 91 8a 8b 88 88 85 8c 7e 88 88 8d 8a 91 8c 8f 82 82 7f 76 69 67 6d 72 65 62 5f 5f 65 60 5f 5f 67 5d 64 54 52 50 51 5f 5b 61 4f 4e 40 2a 1b 0c 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 0c 14 20 28 3e 4c 4f 66 6d 72 64 56 4e 56 58 5b 63 62 5f 68 6b 6e 77 81 84 7d 86 88 8a 8f 93 92 86 82 8f 8b 94 9c 9b 98 a2 9b a8 9a a1 9f a5 9f 99 9e 96 9a 9f 9d 99 a0 96 94 a1 9c a0 97 9d 96 9a 9e a4 99 a2 a0 a5 b2 ac ad 9f ae a8 a2 9d a0 a0 a0 98 9d 94 9d 9a a3 9b 94 94 94 8c 87 91 92 8f 90 90 94 92 9b 93 8f 99 91 8a 92 85 85 68 4f 25 12 09 05 11 08 0b 0b 09 06 06 06 03 0a 06 05 06 00 06 05 06 06 0d 0a 10 0e 07 15 1a 1c 66 a5 be cb ce d5 d0 c5 cd d0 cd d0 c0 c0 b0 ad aa 9b 93 8f 87 8a 82 86 7f 7d 7b 78 78 7b 7e 7b 77 79 85 7f 85 86 7f 85 8b 81 7e 7f 82 87 7d 82 88 85 87 8d 93 8e 95 8f 8a 8e 8a 8d 88 84 83 80 84 81 89 8e 88 8b 7b 75 6c 70 62 65 6c 5f 60 63 5e 60 5e 60 60 64 5f 59 5d 5c 56 4f 50 53 5b 5f 58 4c 3a 29 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 20 2a 34 3f 43 50 60 69 66 56 56 49 51 5a 5d 65 6d 62 67 5e 66 6c 71 79 7f 80 84 86 87 8d 8a 8d 8f 84 8b 8f 93 96 9c 9a 9f 9e 9b a2 ab a1 a3 9f a0 9e 97 9e 9d 9b 9d 92 9b 93 9e 90 9b 9d 9f a5 a1 95 9c 9e a1 a0 9d a8 aa a2 9f 9a 9a 9e 94 a1 9f 97 94 97 96 99 9c a1 98 8f 87 8b 8f 8b 8f 8d 8b 8e 91 91 8f 97 94 8d 90 90 93 8d 89 72 59 2a 12 08 07 0a 07 06 0b 06 08 09 05 0a 03 06 05 03 07 07 05 03 09 09 0e 06 07 09 06 14 1f 61 ac c0 c7 cc cd c8 ca c8 c9 c7 c4 c8 c2 a5 a9 a5 99 99 8d 87 82 84 78 7b 7d 7a 78 79 79 7e 7d 80 80 82 8b 85 84 81 86 89 86 86 83 7f 7b 7c 86 84 84 88 89 95 9c 94 93 8f 8d 85 82 7c 85 7b 80 8a 8c 86 80 7d 7f 79 79 6a 67 63 66 65 62 60 57 62 63 62 5d 64 63 5f 60 59 5b 4b 52 51 50 5a 5e 5e 48 41 22 1c 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 26 35 42 4b 5b 66 68 60 5c 52 50 59 55 64 5e 67 68 69 6b 6b 6c 6b 73 7d 81 84 7e 83 82 8a 8e 91 91 94 91 92 91 94
 a0 9f 9a a4 97 9e a5 9f a2 9d 9a 9b 9a 9b 96 98 9e 96 9a 97 95 98 a1 9a 9e 97 97 9a a3 9d a1 a4 a6 a2 a5 ac a6 98 98 92 9c 94 95 90 93 99 94 99 a1 93 93 8c 92 83 92 96 88 87 89 8f 93 97 8c 90 8c 96 92 88 8d 87 77 59 27 0f 08 05 07 0b 0a 0d 03 00 06 05 07 09 06 09 07 04 06 05 03 07 06 0c 0f 0f 0e 0e 17 20 5b aa c1 ce d0 cf c8 d0 cd ca cb b9 bb b7 ba a6 a6 9a 9a 94 87 8a 8a 84 7d 86 78 7f 82 7b 7a 7c 84 7c 85 82 86 82 8a 8a 89 84 84 86 8b 8d 8e 84 8c 88 93 93 8d 99 93 92 85 88 88 87 83 80 7b 86 85 81 82 81 80 7f 6d 6f 6d 67 73 62 67 63 5e 66 67 60 67 60 60 65 68 65 64 51 4e 55 56 4d 53 5f 5a 47 43 2e 1b 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 12 1a 1d 3b 39 4d 58 58 63 65 59 4d 53 50 52 5f 64 60 66 6c 60 67 6a 6e 6d 74 77 80 80 8a 85 8b 87 83 8c 8e 8b 8e 89 91 9b 9c 9e 9a 96 99 97 9f 9b 9f a2 9a 94 9c 92 95 9c 95 9a 90 95 90 95 8e 9b 98 95 9d 93 9a 9f a5 a4 a1 9c 99 9a 90 98 97 98 96 91 8e 92 91 96 9b 9a 90 8c 88 89 8d 8a 90 8a 8c 90 93 8b 8d 8b 91 93 97 96 8b 91 86 81 5b 2c 0d 06 05 05 0a 06 05 03 07 07 0a 05 00 06 05 08 00 06 05 03 05 0d 0c 03 06 0d 17 0c 23 54 a8 bb d0 cf ce c9 c9 c5 bf c4 c2 bd b9 b0 ad a4 9c 99 8b 8a 87 81 80 74 84 79 7d 7d 77 83 86 85 89 85 8e 8e 8d 88 86 89 8a 8c 87 8f 90 8f 8d 90 8a 83 8a 8e 95 87 8a 84 82 7b 7a 7e 7b 7a 7d 7f 82 81 7b 6f 6e 6c 63 6a 65 69 5c 5a 67 5a 63 67 64 60 60 61 60 5a 58 57 53 52 4c 52 49 4e 5e 59 4b 44 2a 20 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 1f 26 2d 39 4d 4c 57 6a 60 57 4b 46 54 56 5d 64 65 74 65 6a 6d 68 68 68 6d 70 70 72 7b 7e 89 89 8f 92 8f 88 91 8d 90 92 8f 95 93 92 91 8c 9b 9c 96 8d 99 93 92 95 93 97 91 93 95 90 94 92 9a 9b 9d 8d 9c 99 99 a2 a3 9c 9e 98 a1 96 96 8e 90 97 88 91 8b 8a 9a 97 9b 8f 8b 87 8b 8d 8b 86 92 89 8d 89 96 95 97 9a 8d 99 92 88 94 81 83 79 65 24 10 06 05 03 06 08 05 03 05 06 05 03 00 06 05 03 03 06 05 03 06 07 07 08 0e 11 11 19 20 53 a8 bf ca c9 c9 c0 c7 bb bc ba c4 b9 b6 ab aa a6 a1 9c 8d 8b 8a 89 85 81 7f 79 79 7d 7a 7f 7b 83 87 8e 8d 89 9a 94 8c 8f 7e 90 86 8b 88 8c 8c 89 80 7b 8d 87 88 7f 83 85 7e 7e 72 7f 7b 78 7a 78 7a 72 6f 6a 62 60 6b 65 61 65 60 66 61 65 67 71 65 6b 5f 60 5d 54 56 4f 49 4a 45 4c 52 54 58 56 4e 3e 32 1b 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 0c 18 2d 37 41 4c 4b 54 5d 55 5d 4f 4a 53 4d 5a 5e 70 74 73 71 6a 5e 63 60 66 6c 69 78 75 79 7c 88 83 8a 90 8a 91 87 8d
 8c 8c 8b 93 92 95 9c 93 90 96 98 97 98 93 92 95 8c 87 8e 95 8d 91 97 89 93 90 96 95 98 95 98 a0 9c 98 9c 94 92 92 8f 94 92 8b 8e 92 8c a2 96 96 93 84 86 8c 84 8b 85 88 83 8f 92 90 93 96 90 91 8d 90 95 87 87 86 7b 64 36 0b 06 05 03 0a 06 05 03 09 06 05 03 07 06 05 03 00 06 08 03 09 09 06 09 07 0e 08 0e 17 52 a3 c5 c8 ca ca c5 c1 bf bc b8 bd b5 b8 a8 a7 9e a0 96 94 95 81 89 89 83 85 7b 7d 76 7c 85 8d 8b 8b 8c 8f 94 91 90 90 92 90 94 80 8b 8f 85 88 83 88 83 83 85 85 7c 82 7d 7c 7c 76 7d 75 6f 75 7e 79 6e 6a 5f 65 64 63 63 62 65 5f 5e 68 64 65 69 66 6d 61 5c 51 53 46 56 4c 4f 4b 52 4b 4c 5c 5d 4a 40 2b 16 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0d 16 13 2a 41 37 4c 53 5a 5c 54 4c 51 4d 52 55 50 5c 64 69 68 6d 6f 66 6c 5d 5d 69 64 63 6f 72 78 87 89 8c 8f 8f 8a 8a 95 92 94 92 8b 93 96 98 8a a1 95 8b 94 99 94 96 9a 8a 8e 90 94 90 91 91 91 96 8f 8a 92 94 96 98 98 9a 9a 8f 98 94 94 8b 8a 91 99 8d 95 97 98 8c 8f 8b 81 86 84 88 8b 84 8d 8e 89 91 91 97 96 97 9a 9b 91 88 8f 7f 7c 7b 63 2c 10 06 06 03 0c 06 07 05 00 06 05 03 00 06 05 03 00 06 05 07 02 0a 0c 09 06 06 0c 10 1d 46 96 ba c0 c8 c6 b7 bf bc c0 ba c0 b4 a8 a7 a4 96 9c 95 94 8f 90 85 80 8b 85 85 85 81 86 88 83 8b 83 8a 86 87 8e 8c 90 8b 84 89 82 8b 86 77 7b 86 84 83 7e 77 81 81 71 76 7d 79 7a 76 76 73 76 73 72 6e 60 67 63 60 64 65 62 62 61 65 62 65 6c 6f 63 65 6a 5b 61 58 4c 55 54 4c 4f 43 52 4c 5a 5a 4c 42 2c 1b 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 24 31 3b 4c 4e 51 59 56 4d 45 4d 49 53 4b 57 59 54 6a 6f 6d 71 65 74 66 65 61 67 69 67 70 74 70 7c 83 88 88 8a 90 88 8f 91 86 90 99 8e 8e 8f 90 91 8b 8f 92 92 91 8e 8a 96 8a 91 8f 90 95 90 93 8d 8c 8f 8e 91 95 93 97 91 93 97 85 90 8f 8a 8d 8e 89 94 92 95 8a 8b 89 88 85 87 7f 82 8a 90 9a 91 91 8d 97 96 94 8e 92 8f 89 86 81 87 7e 5b 27 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 09 03 00 06 05 0a 09 09 09 0e 19 3f 98 bb c1 c5 be b5 bc bd b5 b4 ba b0 b0 a6 a1 a4 98 8e 92 93 8d 88 8a 87 89 88 8b 88 8b 89 8f 8d 8c 91 8a 88 8e 8a 84 82 83 8c 7a 86 84 7c 7a 80 80 7c 7f 75 77 76 73 79 7a 6d 6f 75 7a 75 72 71 64 60 62 5f 5d 58 5e 5e 5b 62 54 5d 64 62 5f 61 5f 6a 5a 60 60 52 4f 4a 4f 43 4f 46 45 53 52 55 45 34 2e 17 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 1c 1b 2b 39 41 50 52 57 5b 58 4a 48 41 56 50 5c 52 5b 65 5e 6b 69 6c 6d 6f 6c 69 66 5f 61 6f 69 72 7c 7e 7e 8c 86 93 8e
 8f 91 8a 8c 95 99 8e 99 90 8b 90 91 91 90 8e 8f 8a 91 95 88 8e 95 92 8d 8d 8f 8f 92 95 94 92 94 90 98 91 8e 8b 8b 89 88 8d 94 8e 93 96 8e 7e 88 8b 84 85 88 80 8a 8b 88 90 86 96 94 95 93 91 91 93 8a 88 98 80 7c 7e 5a 2a 0a 07 05 03 03 06 05 03 00 06 05 04 00 06 05 03 09 06 05 03 09 0b 05 03 04 13 0e 0c 15 36 8e b2 bd c5 bb b8 c1 bc ba b3 b4 a6 a9 a0 a9 9d 9b 97 90 8e 91 8a 8b 85 89 8c 8e 8b 8b 8f 8e 96 8f 94 8a 85 86 86 84 87 80 89 7e 7b 87 82 7a 77 79 7f 74 83 7e 6e 70 73 7d 71 76 77 6f 70 73 6f 62 62 65 66 5d 5c 58 5d 64 5c 69 5d 65 60 5a 5e 56 64 5f 60 52 4e 4f 55 46 50 4c 55 4e 49 59 56 40 32 24 15 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0e 14 1c 29 42 4b 50 4e 58 51 4b 55 49 4f 4d 49 54 57 55 5e 54 5f 6c 66 69 66 64 6b 64 63 67 62 64 74 6d 7b 7b 78 80 8b 8d 8c 92 8e 92 94 8b 8a 91 9a 94 90 92 90 89 8d 90 8a 93 8d 98 8f 8e 8f 88 91 89 92 8e 8a 94 90 90 94 8b 8b 92 8b 90 8c 8e 98 90 8d 93 86 8b 86 82 7f 7e 82 8e 84 8a 8e 89 8a 8f 91 91 92 92 8d 96 8d 86 87 89 7b 78 76 65 30 05 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 09 05 11 06 0b 0c 15 41 8d b1 b9 c0 bb b5 bf b4 b5 b3 b7 ab ac a2 a1 a5 98 98 93 8f 94 87 8f 90 8b 86 90 8b 86 93 8f 96 8f 8c 8b 8b 89 8a 82 85 7c 82 7c 7e 7e 76 78 7e 7d 76 77 78 78 76 75 76 75 70 70 78 77 70 67 5d 64 5d 63 5d 5e 59 66 59 64 62 5d 61 62 5e 59 58 56 59 58 4b 52 50 4d 54 44 49 4b 48 4e 51 51 51 42 30 24 13 0f 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 17 23 3b 41 47 51 52 5b 59 4d 47 4d 46 4d 51 46 5a 55 50 5a 59 69 6a 65 65 62 6b 65 60 5e 67 71 62 71 71 76 6d 79 8b 88 8a 90 92 8c 8d 8f 90 87 96 92 8b 8a 8b 8f 8d 89 8c 89 91 8f 8e 91 85 8f 90 92 8e 91 84 80 88 88 8d 8a 85 91 87 86 94 91 93 97 8d 89 8c 7c 86 89 88 85 85 88 85 8a 88 89 88 90 92 92 96 90 8b 84 86 85 83 7c 73 74 72 5b 26 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0e 0a 10 29 85 ae b5 be b9 b1 ae b3 b8 b3 ae ae a7 9d 9f 96 96 96 8e 90 8c 8b 8f 89 90 86 8c 89 89 8a 97 89 8a 8b 84 7f 78 7c 78 77 82 73 7b 7a 7e 74 78 7d 71 72 74 6e 75 6f 6f 74 74 73 72 76 68 62 66 5f 63 66 5c 60 62 5d 64 5a 63 61 68 5e 5c 54 55 56 55 56 5b 54 4b 4b 50 4c 50 52 4f 4b 4e 4c 51 4e 3b 2b 20 1b 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 08 19 22 31 40 48 51 52 5e 5b 4a 4a 46 3a 46 47 4f 55 51 54 59 5c 61 61 62 62 61 67 60 5f 61 65 65 61 66 63 75 75 7b 89 7b
 84 89 89 84 94 86 91 8e 92 9f 8a 8c 99 90 8d 87 88 8e 8b 8e 8b 85 8d 86 8c 8e 92 98 8e 90 8a 83 8c 88 8c 8d 8b 8e 92 8e a1 99 94 90 8f 89 83 82 84 8b 88 87 85 81 83 8e 90 8d 9a 8c 8d 89 85 86 8e 85 7f 77 7f 78 7c 5d 2d 03 06 05 03 07 06 05 03 00 06 05 03 00 06 05 05 00 06 06 03 03 06 0b 0e 01 09 08 0d 10 2a 7b b2 b0 ba b8 b1 b4 bc a9 b2 b0 b0 a2 a3 95 96 9b 96 9b 92 92 94 86 85 8d 8f 87 90 92 92 92 8f 8d 8d 88 84 7f 81 7b 74 7b 75 75 7e 79 79 73 76 7f 77 70 73 72 72 74 7b 6e 7b 70 69 66 5e 60 5d 62 5f 60 5a 5c 58 5a 64 5e 67 65 62 6a 5b 5a 56 49 56 4f 55 4f 50 53 4e 51 4f 48 50 4d 4d 4e 47 36 2b 1e 14 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 18 1d 23 37 40 4c 50 58 59 55 4b 49 43 48 4c 4d 44 50 4d 5a 5e 5b 61 5f 59 5d 59 56 5f 65 5f 6b 67 6c 65 66 70 6e 6f 7b 7c 81 87 85 86 84 8a 84 8a 92 90 95 92 91 91 8c 87 8a 8e 8e 86 86 87 81 8a 89 8a 92 93 91 89 87 89 8a 8d 8d 8d 88 8e 94 97 9b 90 97 90 86 8a 87 84 89 7b 8c 85 95 8e 8a 8c 92 8f 8e 8b 8d 8d 89 8c 88 8a 82 7c 75 78 72 4d 20 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 09 06 11 10 2d 7e a8 b5 c0 b6 ab b4 b6 ad ad ae 9e a9 99 9a 9a 92 9a 9a 8b 93 8b 92 8c 8e 90 90 9c 9d 9b 98 90 8a 84 81 85 7b 83 7a 73 78 7a 74 76 7c 6d 6d 7a 74 73 77 70 74 78 75 74 7f 77 72 6f 67 66 5b 5e 61 5b 62 5d 56 60 6a 5e 64 61 68 5b 5f 55 57 58 51 51 50 5c 55 4c 4d 4e 4e 52 4b 4d 43 4b 4d 39 2f 2a 2d 14 11 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 0b 1e 30 37 45 56 4c 50 51 4d 48 3e 3a 48 48 4c 4f 4f 50 50 5f 57 4f 5a 54 52 5f 59 57 5a 5e 5d 5e 60 62 68 70 6f 67 72 7c 7b 7c 7f 84 80 87 7f 89 86 8a 91 91 8e 90 93 8d 8d 83 80 84 83 8b 85 7e 89 86 86 8a 89 8e 8a 8d 8a 85 89 8b 8d 8c 8b 91 97 86 8c 8b 83 8b 84 88 8d 86 85 8c 8a 87 8d 8d 8b 8b 8e 89 89 84 82 7e 7b 80 7e 7a 74 79 72 59 28 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 08 0e 0a 2e 6b ab a8 ad ad a3 af ad ab ab a7 a6 96 98 95 95 9a 92 8c 8a 86 8d 8e 8b 8f 8e 8f 95 98 94 8b 8b 88 80 76 81 80 77 77 7a 6d 74 6f 6c 78 71 77 78 75 74 71 74 78 6d 7e 74 71 72 68 69 61 56 5e 58 61 57 5b 5f 63 5f 63 5d 5b 5d 5e 61 5c 55 55 4c 47 49 4e 4f 54 49 4e 4c 4d 46 4b 4a 45 46 43 35 28 22 24 10 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 19 24 35 47 52 4d 4d 54 50 44 4d 44 47 4c 47 49 58 4f 54 52 51 4e 53 4d 60 5b 56 58 58 5f 5d 61 5b 5f 5d 66 65 72 75 70
 76 7e 80 81 86 79 85 7b 7f 8a 84 88 8f 8b 89 94 8c 87 8d 82 8c 86 84 84 8a 8c 89 93 8b 90 92 92 8d 8d 8b 8f 90 8f 92 94 92 8e 88 87 87 80 81 82 86 90 8b 88 88 90 87 8b 89 8a 92 86 81 88 7c 75 73 7a 76 71 81 6f 77 59 1f 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0d 08 09 0b 0f 24 71 9f a0 a9 b1 a4 b5 ac a9 a8 a0 9f a1 96 8d 92 8a 92 95 8e 91 8f 8b 87 8e 94 91 9b 9a 8c 8e 8d 7c 84 80 80 74 76 70 71 6e 71 6e 71 75 72 6f 72 74 73 74 6c 78 7b 7b 72 74 6c 70 66 5d 59 5e 57 53 59 5c 5a 5c 59 65 5e 5f 5b 59 56 59 52 50 4b 4d 4f 49 53 52 4e 4e 4d 48 4c 44 48 44 44 41 2f 29 25 1f 18 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 1f 20 2c 3e 50 4a 55 51 58 52 4e 42 42 3c 46 44 49 52 4d 51 56 55 49 49 54 54 54 50 55 51 57 66 5c 58 67 66 6e 6a 6f 74 74 6f 75 7d 79 82 80 7c 80 7d 80 86 83 8c 89 90 90 96 8f 8a 88 7b 87 87 89 8f 90 8d 94 90 85 88 8e 8c 83 91 94 8d 8c 8d 8a 8c 8b 84 88 84 8c 80 86 8c 8c 94 8e 8e 91 89 8e 95 85 8d 88 86 80 7b 7b 85 7b 6f 78 72 6e 6a 5a 1b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 08 03 00 06 05 03 0e 06 10 0d 0e 1d 63 a2 a9 ac a5 a3 ab a6 a1 a6 a9 a6 a4 99 90 91 97 91 8f 89 89 8d 90 98 8d 93 97 94 9b 87 8c 84 84 85 7d 7f 7a 71 71 70 74 70 6c 74 75 70 74 76 79 70 70 7e 75 77 72 74 6c 70 6e 62 61 5f 5d 61 59 55 5c 60 5a 60 64 5e 5f 5f 58 55 53 52 52 4f 4e 53 52 53 56 51 50 4d 48 48 48 4a 4d 3c 3a 31 21 20 19 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 15 0c 1d 2f 38 4b 55 57 5c 55 52 4c 3e 46 3f 4e 49 4f 52 4e 50 53 4b 47 4e 4c 52 55 55 4e 51 54 5a 60 5d 62 65 69 63 69 71 6c 6a 7a 74 72 7b 83 7a 82 84 81 76 77 80 86 86 8b 92 8a 87 8e 8c 8a 8a 92 8f 8e 8d 91 8e 8f 8d 8a 8e 92 8a 8e 8a 85 82 84 81 7d 79 81 88 80 8c 87 91 8e 8d 80 8a 91 88 8c 8d 83 87 84 78 80 83 83 72 75 76 6e 7d 6e 69 57 21 09 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 0c 07 12 09 06 1c 62 98 a2 aa ad a7 ac a6 a3 a3 a1 9a 99 97 9c 98 94 9c 94 8b 8d 8a 8e 92 93 98 99 96 93 96 8d 89 83 79 7e 73 75 71 6a 72 67 6b 63 69 75 6e 73 75 67 6d 72 75 7b 6c 6e 6d 6b 60 6d 59 5c 53 54 5e 58 56 55 5d 5e 60 64 59 5f 54 58 52 50 52 4f 52 4e 4c 4c 4e 51 4d 4d 46 48 49 4c 48 4e 3a 31 29 22 21 14 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0b 17 2a 31 3d 4f 49 53 59 5c 4b 49 47 44 46 47 49 4c 4e 4d 4b 44 4b 51 54 4f 53 4f 51 51 5a 58 5b 5c 5e 60 65 63 67 68 63 6e
 69 6a 70 73 72 79 79 80 7e 7d 7c 74 7b 81 84 8d 90 86 8d 99 8f 93 8d 80 90 7f 8e 84 8d 8c 88 89 91 8a 87 84 78 7c 86 7f 7c 87 84 8e 84 8a 86 7d 8f 8c 8f 93 93 93 91 8a 84 85 81 80 83 79 7f 7e 7a 76 78 73 74 6f 71 55 21 04 06 05 03 00 06 05 05 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 06 00 06 05 08 09 1a 58 9c a0 a1 a4 a1 a9 9b 9b 99 9c a2 9a 9c 90 9b 98 91 8c 93 99 91 94 87 97 92 99 93 91 96 81 80 7e 7b 7b 77 7a 70 6c 67 71 67 6a 6d 6b 6c 65 6d 70 73 7a 6e 77 71 71 6b 6e 64 5a 5f 59 55 59 5b 54 58 57 55 5d 58 65 65 61 5d 54 56 4a 57 42 48 52 4a 44 52 49 3f 4b 50 42 46 49 49 47 38 3a 2d 22 1a 16 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0c 12 2c 2d 49 54 55 52 57 5a 48 4b 3c 42 46 42 4e 4a 46 4a 4a 4e 44 4a 52 4d 4f 51 52 55 52 5a 5b 5a 5a 5d 62 63 61 67 6c 69 6c 6f 6f 6d 76 7b 83 7a 80 7d 7f 80 7c 80 77 7e 86 98 98 97 94 92 8c 94 87 8a 8c 84 85 8b 85 8c 82 86 88 84 81 84 84 82 84 83 8d 8a 8d 8f 85 87 90 89 8c 8d 91 94 87 87 87 89 82 82 7e 79 79 7b 74 75 74 71 6e 6d 74 57 28 08 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0b 11 10 4b 91 9f a4 a2 9d a5 a0 a0 9f 9a 99 a0 92 96 96 94 96 90 91 90 90 94 94 a0 99 95 95 89 8c 8c 85 79 77 76 6d 72 6d 6f 6d 6d 6f 69 6f 69 69 6f 72 6a 76 6f 7e 73 6e 71 66 67 5c 5e 61 5d 5b 53 5d 57 5c 61 60 64 53 63 61 62 55 54 4d 4e 4c 4b 4b 4e 4c 4e 4a 4c 4e 50 55 49 4d 46 4e 46 3e 2f 20 20 24 17 13 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 14 1d 29 33 41 50 55 61 5c 55 41 48 41 4b 3c 49 47 4b 4e 4b 49 47 48 49 4f 4f 51 4e 52 56 58 54 59 57 5b 62 5f 65 65 5f 65 66 67 66 6d 69 69 72 6d 75 7d 82 81 7b 7e 7f 82 7f 84 85 8e 92 92 96 92 91 85 7b 85 83 80 7a 82 85 88 84 7d 84 82 8c 79 88 87 80 85 89 8a 8e 8e 8f 95 91 94 89 8a 88 87 88 81 7d 82 7c 7a 82 78 73 73 74 78 71 70 71 68 5a 22 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 03 00 06 05 03 06 07 05 03 00 19 4d 8e 98 a3 a2 98 9c 9a 9c 9c 9c 9c 98 99 92 95 98 96 94 96 9b 9a 9c 95 a1 95 9e 96 82 8a 81 80 80 7b 73 70 72 6b 6a 6b 60 6c 68 70 67 6a 6d 6f 72 79 70 71 64 66 6a 64 62 5a 5d 5a 56 50 50 54 5a 54 53 5c 5d 61 59 64 5b 5b 54 52 59 4c 53 52 49 4a 4b 4a 48 4e 4a 4d 48 4a 47 48 49 40 30 25 21 1f 14 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0b 1a 19 26 34 42 4e 52 64 5a 54 48 42 47 40 47 4f 3d 43 47 46 43 4b 4c 4c 41 4b 48 43 5a 4c 53 4f 51 58 59 60 5e 63 68 63 5f 65
 63 70 6c 6c 61 6b 69 67 72 71 76 7f 80 75 86 84 7e 87 88 95 8f 92 94 89 87 8d 81 7c 84 80 7b 7e 80 7a 84 84 7f 85 84 7e 86 83 88 91 84 91 8d 94 8b 88 8f 93 85 8b 8b 7e 83 81 84 82 78 7b 75 75 75 71 73 73 69 70 72 5f 26 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 0a 03 06 15 49 92 9d a5 a3 a0 92 96 9d 9b a0 9d 99 9a a1 99 9d 94 9f 95 9e 91 9f 95 9d 97 9e 9a 8a 8f 85 7e 82 6d 74 74 6a 73 64 6e 69 68 69 70 68 6a 6b 70 75 73 70 66 6a 62 63 5f 67 59 50 50 54 53 58 4e 4d 57 58 5e 5d 5d 61 5e 58 5e 5e 51 51 4a 4d 4a 4a 49 50 47 45 4a 49 46 48 48 49 3d 46 32 32 20 1b 1a 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 17 1c 29 32 45 58 59 67 61 59 4e 4c 3f 40 44 40 44 4a 47 44 4b 43 50 45 44 43 47 50 51 4e 53 54 49 5d 55 52 62 61 60 5f 65 6d 63 6f 67 65 69 6a 6f 6b 68 69 70 73 79 8a 83 86 80 87 86 85 87 86 8b 82 89 84 7d 85 80 7c 80 82 81 88 7d 7c 79 82 82 84 8b 86 8c 94 83 8b 8d 83 8e 90 8f 86 87 81 82 84 87 7b 82 75 84 76 7b 76 76 7a 77 7a 75 72 6e 5a 22 03 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 05 0b 4a 8d 9f a2 a3 9f 9e 9d 94 9b 98 9b 9e 97 99 95 98 a0 9d 9a a5 97 a3 99 97 9c 9c 95 90 86 89 7f 7d 6f 71 74 6b 68 6f 63 70 73 69 68 6d 6b 6f 74 6c 6d 71 6a 67 67 60 58 57 56 5c 53 59 4e 4f 51 57 5a 58 5f 5c 5d 5f 62 5f 5b 62 4f 5b 51 4d 51 48 4f 4e 44 4e 4a 52 4a 4f 50 47 47 43 38 2b 20 1f 17 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 18 33 39 4a 5a 58 66 61 61 53 4c 41 4a 47 47 4b 4b 4b 50 50 42 46 46 42 4e 4e 4e 4c 4a 4f 51 4f 56 5b 4f 54 58 63 60 69 63 62 65 67 6a 65 61 66 6a 69 6e 67 6a 75 75 80 82 83 8e 88 88 85 82 8d 7d 84 81 7c 81 7c 74 81 82 7d 82 83 81 7a 7f 83 80 82 7e 88 8b 93 8e 8d 8e 8b 87 88 93 89 8a 85 89 81 78 85 76 74 7c 81 7d 76 71 75 6d 6e 73 72 5e 25 0a 06 05 03 01 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 04 00 06 05 03 08 11 44 89 a0 a1 a1 97 99 a0 99 9d 94 9e 98 a1 a1 a2 a1 97 9b 99 9b 9c 90 92 93 92 91 8c 84 88 7f 78 77 82 75 75 6d 6a 64 66 5e 6b 69 64 75 61 70 6d 69 6d 66 61 5d 59 54 5a 58 57 59 5a 52 4e 51 56 53 50 54 5a 54 56 62 5a 55 58 5f 58 51 4e 4e 50 44 4c 4c 47 4a 46 4b 47 4a 50 46 49 40 2b 2f 20 25 13 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0c 0b 20 20 2e 43 53 53 60 69 64 4f 44 49 3f 3c 49 42 43 3f 4d 48 42 4a 44 46 4a 44 4d 44 48 4a 44 4f 50 55 59 57 59 62 60 63 63
 68 62 61 60 5f 62 65 66 61 66 61 6f 6a 6a 72 7e 7c 81 89 88 87 83 87 87 8b 82 77 7c 7c 7c 7d 7d 7a 76 71 83 7e 78 78 7e 89 73 8e 84 80 8b 85 8f 87 83 8a 87 7e 83 80 7b 82 78 7c 78 77 74 6e 75 76 75 70 71 6a 70 69 5f 2d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 3b 84 94 98 99 94 9c 9b 9e 9d 9e 9b 9b 99 a1 9a a0 9e a3 95 9b 9b 98 89 85 8a 87 81 7e 7d 81 80 7a 72 6a 6c 68 63 67 65 67 64 60 68 69 68 6a 6d 69 60 5f 5f 56 50 57 56 51 55 4d 4d 58 47 47 52 51 57 51 49 54 50 57 4f 56 53 5a 50 5c 43 4b 48 46 48 4e 45 4d 43 49 4c 4a 45 41 47 46 29 22 1a 1c 13 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 13 20 23 32 41 52 59 6a 68 68 5a 50 42 46 3f 4a 40 49 41 46 4b 4b 3f 49 49 4a 4c 45 43 40 49 4b 4d 56 51 52 53 5b 5c 61 65 64 61 67 57 64 66 5c 68 62 66 60 61 66 64 65 72 73 72 80 83 86 86 84 83 84 80 7f 87 7e 7c 77 70 78 7b 7b 7f 7e 7b 79 7b 77 81 83 83 84 82 8d 8e 8a 8c 8b 82 8b 88 7a 81 83 76 77 77 76 6c 75 75 7d 72 6f 75 71 6f 74 70 61 26 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 10 39 86 96 9b 9b 99 99 9a 92 91 98 97 9f 9e 9a 9b 9b 9b 94 94 96 97 96 8b 8c 7c 82 76 7f 77 73 6d 73 71 6b 69 5c 63 6f 67 67 6c 69 6d 6c 61 60 5e 60 60 5c 51 54 56 55 55 56 52 4f 50 50 56 4f 57 53 52 51 56 5a 53 4d 53 51 4f 4f 5b 53 46 48 48 4d 4e 47 4d 4b 41 44 48 43 44 42 48 3d 34 29 21 14 11 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 08 14 21 1a 2c 41 4a 52 66 64 6c 5a 53 4c 45 48 46 43 41 47 3d 43 44 3e 46 42 44 48 48 48 47 42 4b 4e 51 57 56 55 56 5c 56 5e 5d 61 62 65 5c 58 5f 60 59 59 62 5e 60 63 6a 66 63 6f 77 7f 84 87 86 89 84 80 80 7f 7a 73 74 7d 79 7d 77 7c 79 79 7a 7e 7f 80 80 84 84 82 87 82 82 8a 87 85 81 7c 80 7f 7e 77 76 77 73 70 7a 75 73 6d 70 73 6b 6a 6f 6a 5a 23 07 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 03 01 12 30 79 98 93 97 8f 90 94 9a 97 9a 97 9a 92 93 9b 9b 94 9b 95 96 8d 8c 86 84 77 7a 71 78 79 71 6a 70 71 6b 6a 65 63 62 69 68 6d 69 6f 62 6a 60 5a 5b 56 54 54 4b 53 56 55 52 50 4f 50 4f 4d 56 58 4b 4a 53 54 5f 4f 51 46 47 45 54 54 58 52 44 46 42 47 49 46 4f 49 4c 4b 48 4e 43 42 3e 2e 22 17 16 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 1d 1c 2e 40 45 56 5d 72 65 66 59 45 3d 3a 3f 45 45 48 42 4a 3d 44 3b 43 3f 43 4c 46 48 46 46 4f 50 4d 52 5e 60 5e 5d 64 5e
 5b 59 59 58 5b 52 5b 5c 5b 5c 5c 5a 58 61 5d 65 6a 6a 6a 7d 7b 81 86 86 8a 81 7e 73 75 77 77 73 75 71 70 76 76 7b 6e 79 7b 79 7a 81 7b 82 7b 82 85 82 81 7f 75 80 78 78 71 6d 78 73 7b 6f 75 76 6b 6e 79 73 69 6f 70 69 26 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 35 76 8a 96 95 8f 90 94 91 93 94 97 96 99 8d 92 8f 95 9b 95 8f 8f 7e 80 80 6f 7c 74 76 73 6e 70 70 68 67 67 69 61 66 63 68 6b 65 68 5f 5d 57 58 54 52 51 4a 4e 53 50 49 52 50 4e 56 50 4f 4d 4b 4b 50 51 4a 4b 48 44 3b 45 4b 46 48 46 44 46 4e 3f 45 45 4d 3e 4f 50 46 49 46 45 46 35 25 18 19 12 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0b 11 1a 21 29 39 3f 4f 5e 6b 75 6f 5c 4e 3f 44 41 41 45 41 4b 3f 41 41 46 4e 43 48 48 43 4b 45 46 51 4e 51 53 55 58 5e 5e 59 5d 61 5f 63 5c 5e 59 5c 63 55 5d 59 59 61 61 56 60 66 5f 72 6e 6e 77 7d 80 87 8b 7c 85 79 78 7c 7a 7c 80 7c 79 6e 71 75 76 75 79 79 7e 78 7a 7d 83 85 80 7f 81 7a 79 73 6e 76 70 67 73 71 6e 72 6e 71 6b 77 7f 73 6e 76 5f 2a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 25 71 82 8c 8c 83 90 8e 8c 93 96 92 99 8e 93 95 8b 93 84 85 82 81 81 78 7a 73 70 6e 6e 69 69 63 63 61 61 6d 6d 6f 72 6d 73 68 67 67 53 50 4f 4c 47 53 4d 51 4d 52 4f 4e 4d 4f 4e 54 48 48 4c 4e 49 52 4f 4e 4d 42 44 45 46 4e 49 45 46 46 42 4a 46 4b 4b 48 42 46 46 48 51 49 4b 45 3c 23 20 14 0b 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 07 12 10 20 20 39 40 4b 58 5d 68 74 60 4d 45 44 47 49 49 4e 49 47 3c 4b 3f 4a 3d 42 49 4d 41 43 48 44 4e 52 53 55 52 54 57 55 5d 58 60 5f 5a 5c 54 58 51 60 59 50 59 59 5e 57 62 60 64 61 6b 6b 76 78 7a 76 7f 88 87 85 7a 7e 80 77 76 7c 76 79 7b 71 74 7e 75 7d 79 79 78 7f 82 7a 7b 74 79 7d 7e 77 76 7a 78 81 74 71 75 70 71 75 73 79 7e 75 6f 7b 69 2c 04 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 08 26 67 87 86 92 81 8c 8e 8d 85 8e 90 88 89 89 8e 8a 7f 84 83 81 76 7d 75 76 6e 6f 6c 6f 66 68 6f 64 62 69 6a 64 6d 6d 6a 67 67 5e 54 5f 57 4e 51 51 4c 4f 57 47 4d 51 51 55 53 56 4e 45 47 4d 52 4b 4b 4d 49 3f 42 43 44 40 3e 4c 49 50 47 4e 46 4c 4d 49 44 47 45 4a 4c 4d 4c 4a 3a 39 2e 1f 16 08 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 11 16 1a 28 2a 41 3c 42 5a 68 71 6a 5b 45 40 45 46 48 49 41 48 37 35 3c 3e 43 45 39 44 44 43 41 45 4b 50 4f 54 5e 4b 4b 52 58
 53 5f 56 59 5b 5d 55 5a 58 58 4e 5d 58 50 5e 5e 5d 5f 61 64 67 5f 6f 71 7b 76 7d 81 7b 81 85 7f 7c 7b 76 7b 70 75 72 71 7f 6d 74 76 7d 7e 7a 7f 7c 73 78 77 76 7c 78 74 77 68 71 70 6d 71 77 73 7b 80 8a 89 85 7e 85 6f 30 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 1b 62 7b 8a 86 79 7f 83 84 8b 8a 7c 89 89 80 80 79 83 7d 78 7b 79 6f 6e 6e 63 6f 67 6a 69 65 66 68 65 6e 68 6a 69 69 60 61 54 59 55 4e 4e 4b 52 56 4f 50 4b 4d 3f 4e 4b 49 4a 47 48 55 47 48 52 44 4a 49 47 42 45 3e 4b 42 41 4b 45 44 49 43 42 46 4f 46 4b 41 49 4b 47 4d 4a 41 44 30 2a 1a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 17 16 21 2a 2e 3c 35 4b 60 6e 69 58 49 49 3c 4a 45 47 3f 43 44 42 43 3e 44 4a 44 3a 42 50 46 46 4e 47 52 51 55 57 55 5a 57 59 55 56 59 4e 55 50 54 57 56 55 57 56 5d 4d 5b 5f 53 5e 5c 5c 66 5d 6a 6b 77 79 7f 7b 84 82 80 79 7e 77 7b 71 6f 75 77 72 77 7f 74 72 75 71 75 7a 73 77 76 75 70 70 70 76 77 78 72 70 74 6f 7e 7d 80 83 77 7e 7e 7c 70 2c 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 5e 77 7a 89 79 84 84 7d 85 82 82 83 7a 7c 7c 79 7d 76 6f 70 6a 71 62 68 6c 6e 63 6c 61 68 63 63 5f 6b 65 69 67 66 5d 5a 57 4d 4f 47 44 45 4b 47 4f 4f 4a 48 4d 4e 4b 4f 49 45 4d 47 47 4b 4b 47 4c 49 41 3a 41 39 3c 4a 3f 45 47 40 4e 47 42 43 45 47 43 44 40 46 4e 4a 50 3f 3a 33 22 15 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0d 14 19 1c 27 32 35 33 42 52 60 75 65 52 48 47 41 4a 44 4b 43 4a 48 48 44 40 3e 4c 4a 40 47 3d 45 4c 4e 50 55 57 4e 51 53 55 58 60 60 58 56 52 5c 5a 54 60 5c 58 55 59 56 53 56 60 5a 64 5b 60 67 64 6e 60 69 71 7f 78 81 84 7f 86 7a 84 80 7c 74 7a 73 7a 74 7a 79 70 76 79 6e 7b 7a 6e 6f 70 73 72 6d 70 78 77 73 7b 79 77 75 74 76 7c 77 7b 74 65 31 08 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 06 15 5b 72 76 81 73 7d 81 84 76 80 82 80 78 7c 82 75 76 79 70 6b 71 6b 66 6a 67 5f 6f 6a 64 67 6b 6b 64 68 68 63 5c 5a 52 51 52 51 50 56 4e 47 53 4a 50 50 4a 45 40 4a 49 4a 4e 48 47 4d 45 48 4c 4a 4b 46 47 44 47 46 50 4e 40 44 3c 4d 4a 49 4b 4f 40 4b 4c 49 51 43 4d 4c 48 45 34 2b 1f 0f 10 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 17 15 19 28 28 2b 38 3a 41 56 62 6a 56 48 4a 3e 41 49 47 3e 4b 44 48 44 45 46 44 42 44 42 42 46 42 45 48 4d 58 4a 4c 49 52
 5c 61 5a 59 5e 56 5b 60 5a 5b 4e 5c 5d 58 59 59 51 60 57 61 55 60 5d 5d 5d 59 62 6b 62 6b 75 7e 7a 7e 79 78 81 81 73 7d 74 7a 7a 74 77 74 71 63 79 6e 72 79 73 70 71 74 74 72 66 69 71 74 76 78 7b 70 72 6d 6f 74 6e 68 36 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 1b 4b 7d 7e 7d 78 7c 79 72 7c 77 78 7a 74 6d 72 64 6f 70 71 6e 6b 64 5e 68 5e 67 64 66 69 66 66 65 64 5d 61 5b 5f 58 4f 4b 4d 48 4f 4c 48 4b 4d 4c 49 48 44 43 45 3d 48 48 4a 47 48 4b 48 40 3d 43 4c 47 49 3f 42 3c 40 46 46 46 47 48 41 43 4e 3c 44 48 4c 4c 4f 46 4d 51 55 41 34 24 18 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 0a 17 1d 25 29 2a 32 3d 53 61 67 5e 46 4a 44 44 46 3e 48 42 46 4b 44 4c 48 47 45 4e 42 46 48 47 3f 4d 44 4e 50 53 5a 51 4f 5a 53 5e 60 5f 5f 62 63 63 5c 59 5a 5b 60 60 60 5a 5f 5b 5b 53 57 55 5d 56 5d 60 62 62 66 69 73 7d 7d 89 85 81 7d 84 7d 7e 7c 69 70 71 6d 76 70 69 6d 75 70 73 6e 70 6b 75 75 71 72 76 7d 71 6f 71 77 6c 6a 66 6e 65 31 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 52 73 74 78 70 6c 73 79 72 6f 71 6f 74 6c 6d 6d 6b 6c 6c 68 6d 61 64 64 5f 60 6c 64 64 69 68 68 61 5d 66 5b 54 50 52 4f 4b 4a 52 45 45 48 50 4a 4d 46 48 4d 48 4a 49 47 46 44 4c 44 44 45 4c 3e 3c 3d 45 3c 3e 48 41 3f 44 43 44 4a 45 4b 43 45 4c 3f 48 44 4a 4c 4e 52 49 44 2a 20 0c 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 11 20 29 2d 2e 36 3a 4a 5d 5d 5f 4b 49 3e 4a 41 4b 40 46 43 44 4a 44 43 4b 45 41 40 45 49 49 54 4f 49 4f 45 51 5a 4e 55 5d 5c 5b 58 58 59 64 5a 6a 5e 60 68 60 66 5c 5c 60 64 5f 59 59 56 5c 58 5a 62 5c 65 64 59 66 69 69 73 7c 7a 81 86 83 84 78 77 77 77 6d 74 73 74 72 74 66 71 77 7a 6e 76 79 74 7b 7b 7b 74 79 68 6f 73 6a 66 73 67 5f 38 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 4d 6c 78 71 69 6f 73 75 73 76 6a 68 6b 70 6f 6d 71 6d 67 6c 61 62 5f 67 66 65 5e 66 63 60 6c 5d 5b 5b 52 4e 4d 50 4f 45 48 48 4c 45 46 50 48 54 4d 4f 48 45 3f 44 46 48 50 46 43 43 40 41 45 40 42 4c 47 49 3d 44 42 41 49 52 47 4c 42 48 40 4b 47 4d 4a 48 4a 48 5a 56 4f 34 33 21 05 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 19 16 1c 24 26 35 38 43 56 5e 5a 4f 4c 3e 49 44 4c 48 3f 41 4a 43 4c 4a 4d 4c 47 47 4a 4b 4a 4d 44 44 47 48 4c 4e 52
 4f 59 55 54 5e 5e 61 62 6b 5d 63 5c 65 68 5f 5d 68 5b 5a 55 5a 59 55 5c 5e 57 52 51 5d 5a 58 64 67 66 63 6d 65 77 7f 7b 85 78 7e 7b 80 6f 6e 72 75 74 6e 76 6e 6d 74 68 76 75 71 6f 71 7e 73 72 72 78 6d 6e 63 68 67 61 33 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 3e 6e 77 74 65 74 76 64 75 6c 77 6e 69 6a 62 67 62 5c 61 5a 5d 5d 5d 61 59 62 5f 68 63 61 5d 52 53 54 4d 51 4b 4b 49 47 4a 4a 46 45 44 42 4a 4c 48 4a 43 44 48 45 49 44 46 42 40 4a 3f 45 43 48 40 46 44 3b 3a 3d 41 3a 41 4a 44 44 40 47 42 44 47 46 47 46 44 55 53 59 47 36 27 1a 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0e 13 20 1d 23 2c 37 3a 50 5a 60 4a 43 49 49 47 4f 4c 46 4b 4a 49 48 48 4d 4a 4d 46 50 49 43 4c 42 49 4c 4d 53 50 44 4b 52 4f 4a 54 57 5d 5d 62 65 6a 5b 60 5f 5a 64 60 5b 55 52 57 52 5f 4d 58 53 56 55 59 5a 58 63 61 5e 65 5b 6b 6c 72 71 7c 75 7f 7f 72 73 76 7a 76 76 6a 64 6d 6b 70 71 70 76 71 74 69 74 76 78 72 6d 67 65 65 67 61 5b 34 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 40 64 73 71 6b 72 68 6c 64 6e 65 68 65 68 66 62 65 6b 63 67 61 67 5e 60 5c 5b 5f 5c 55 5a 5b 58 52 50 4d 47 40 4e 43 4e 45 44 4a 4b 45 44 49 4d 45 3f 3e 3f 46 48 43 4a 40 44 3b 43 3f 45 39 39 41 3e 3b 42 3d 45 49 47 4c 44 47 41 47 49 4b 46 48 49 43 4a 4d 4b 58 4b 3a 25 1d 14 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 15 17 24 1f 25 37 41 4e 58 61 58 46 3c 43 49 49 47 45 42 47 4d 4a 4a 51 4c 49 43 3e 4d 48 49 49 43 46 4c 50 4c 4a 51 50 4d 4f 52 5c 5c 6a 65 6a 64 64 64 62 5d 5c 62 58 5a 51 52 5a 55 5d 54 56 58 4d 4f 5f 55 5b 5b 53 55 62 62 66 6a 5d 6d 73 76 7b 75 7c 6f 78 75 6e 72 79 6e 6e 76 6e 72 6e 78 76 6c 72 6e 6d 6c 71 6e 71 6d 67 6b 63 39 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 3f 64 77 77 73 6d 6a 6c 63 6e 68 67 68 5e 63 65 62 67 5f 5a 65 5e 5a 64 59 5c 55 63 50 5f 5a 52 55 50 4d 4d 42 47 44 4c 47 4b 49 44 42 4b 4d 4a 43 47 45 4d 4a 47 41 42 40 3b 3b 43 3b 45 3d 42 41 45 3c 40 43 41 42 3f 49 48 40 4b 45 49 49 48 4d 45 4a 4d 44 59 4c 4d 39 24 1b 10 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 01 10 14 1c 2a 2b 2a 34 47 59 67 59 4a 4b 43 4a 51 47 48 4c 49 47 4e 50 4e 4a 41 4a 46 4c 51 4f 49 4e 4b 48 46 47 4b
 4a 4d 51 4f 53 59 60 64 63 69 65 66 66 60 5d 52 5e 54 52 59 51 54 4a 52 51 54 53 58 50 53 53 55 59 57 52 58 59 56 56 5b 67 60 67 74 71 65 75 75 73 75 73 79 6f 73 7e 75 6e 79 78 78 70 74 71 72 71 78 75 67 6d 69 71 65 3d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 35 67 73 70 65 68 6b 6d 69 69 60 63 61 5d 66 63 64 66 66 64 5d 5a 5e 5e 4e 58 61 53 56 4e 4b 53 45 47 4d 44 4f 4f 4e 4d 4d 4b 4e 4d 48 41 50 4c 45 49 43 4e 4c 46 3a 47 44 3c 44 3e 3c 3d 3b 3d 41 44 3d 44 43 4a 42 45 46 4b 46 45 51 45 41 42 4c 4f 4b 4f 47 4f 50 43 38 25 15 0e 03 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 08 10 11 1c 25 2c 39 4d 5b 5f 52 4f 3f 46 41 48 41 4d 44 4d 53 4e 4d 4d 46 42 48 42 4e 4c 48 39 3e 4a 4d 47 45 4f 4c 4e 49 49 51 5b 56 55 5e 61 63 55 60 58 63 56 50 52 63 58 5c 59 52 5a 5c 5b 4c 55 4a 4f 53 50 4e 51 54 56 58 5d 5f 55 5f 5c 65 60 5f 68 6d 64 66 70 74 69 70 73 7a 78 71 72 75 78 6e 71 70 70 71 69 71 72 73 69 6c 63 3e 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 2b 68 67 67 66 66 6d 69 6a 68 61 62 68 5d 65 64 59 65 65 61 5e 5b 57 59 5b 51 55 4a 4e 4c 51 4f 4b 4d 4c 41 45 47 46 47 45 49 46 48 4a 4c 47 4a 45 43 48 4a 47 3d 36 3f 3e 41 3e 39 3a 3d 3a 40 42 43 39 3c 3f 45 43 42 3e 47 48 49 48 41 3d 44 4b 42 45 4a 46 50 4b 35 26 1a 09 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 09 0b 19 22 25 22 40 48 59 64 5a 4c 45 49 47 44 49 47 4a 46 4b 4a 49 4b 4b 4d 44 46 4a 4b 4e 48 4d 50 41 4a 46 4b 56 4d 4a 4d 51 5a 56 52 5d 61 57 5e 4c 60 56 54 5d 5c 5d 67 59 50 5b 51 54 52 59 54 50 55 52 52 53 55 55 54 51 50 56 5b 61 5f 5d 5d 5e 60 63 5b 66 5f 67 67 6c 65 6c 6b 6a 78 78 75 77 79 77 72 70 72 75 6b 6d 70 6e 66 44 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 36 5f 72 6c 68 6c 66 66 6c 68 66 64 67 60 66 5e 67 60 59 5e 60 5a 58 56 54 58 52 56 59 4d 4d 46 46 44 41 41 49 45 45 4a 51 4e 51 48 52 57 4f 4c 4a 47 42 4a 45 38 42 3f 3b 37 39 3f 37 3b 3a 3f 41 41 4a 40 40 41 3e 3c 42 55 43 46 45 4f 4a 46 4b 49 4d 47 46 45 41 2c 2c 12 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 11 1d 1d 27 2a 32 49 52 67 5b 53 47 45 4c 4c 4a 4a 3e 46 49 57 48 54 51 4d 48 44 4f 4b 4a 49 4c 49 4c 46 40 4d
 4e 41 48 4a 4f 53 47 4b 55 58 5c 5c 53 4f 54 4e 5c 5f 5e 65 59 51 56 46 53 51 4d 50 4e 58 5c 55 59 56 59 57 53 5a 56 5a 59 58 57 5b 5e 56 5f 5e 60 61 64 5e 66 6c 64 6f 6b 79 78 7c 72 79 74 74 7b 7c 77 6d 74 75 74 70 3e 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 2c 6c 68 6f 5a 5f 64 64 64 65 6a 65 62 65 65 60 5f 63 63 59 5b 55 55 5a 52 4e 49 49 4e 4b 4f 4a 43 47 4e 48 4b 42 49 47 4e 48 4b 4d 44 54 50 58 4b 4b 4d 42 46 3b 42 41 3c 39 38 37 3b 3e 3c 3d 42 47 40 48 43 44 3a 3d 4a 4c 50 4d 4a 4f 43 47 44 42 46 53 48 42 3f 2c 1d 10 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 0d 10 1a 20 29 30 39 4a 5d 5b 51 4d 46 48 4e 4e 4d 4b 49 48 47 42 4f 4a 48 47 40 3f 4e 40 42 47 44 42 43 47 49 45 4c 47 48 47 47 45 4b 4a 50 44 52 4d 46 47 50 50 5a 53 55 47 4a 4e 56 52 4f 53 4f 4b 47 55 53 52 59 4d 4d 53 4e 4c 4f 54 52 54 56 54 60 63 5c 5d 5a 5e 61 61 5e 66 61 66 6a 71 78 74 75 6e 75 75 78 7b 75 78 72 7f 71 46 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 25 58 6c 71 6a 63 6b 5f 67 69 64 63 60 61 5e 5a 60 59 5a 54 51 59 50 54 50 49 47 50 45 51 46 41 48 44 47 46 41 48 49 48 49 3f 41 50 49 4d 4a 51 4b 43 4f 49 3b 42 3a 3b 38 3a 36 33 3c 3d 40 42 42 38 39 43 3c 41 43 44 44 45 3e 4c 47 4f 4f 4a 4f 4b 4f 52 48 46 38 21 15 0a 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 13 20 1b 1c 36 36 42 56 56 50 4e 4e 4c 4a 40 48 46 46 49 47 4a 45 52 44 48 4d 48 43 41 4d 4a 49 4d 3c 4b 49 4a 4a 4b 49 46 47 44 49 50 4b 4f 43 43 46 4c 46 45 4f 4f 4f 47 4a 4d 4c 4a 49 4d 4c 52 51 57 58 58 58 4c 4f 4b 50 56 53 59 4e 55 51 51 58 5a 5a 53 54 5a 5e 56 68 60 5e 68 62 67 64 73 69 74 70 6c 6e 72 79 74 7d 76 72 4f 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 27 53 67 6c 5d 64 68 64 5a 5e 61 64 62 5e 5d 51 57 5c 55 55 4a 59 4f 4d 4e 4c 46 49 4a 4a 46 41 44 46 4e 47 39 4f 4b 46 4a 46 43 56 4e 4b 4d 4c 43 42 49 40 3a 3d 34 3b 3d 3a 39 37 40 3a 3e 3c 39 3e 39 34 45 49 43 44 46 4c 49 49 4a 4a 4a 49 50 45 51 45 49 3b 36 20 15 0a 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 08 10 19 28 26 40 43 47 5a 54 4b 44 49 48 49 47 43 45 42 41 50 4d 4c 49 3e 42 48 45 4f 49 4c 49 43 4c 4f 4f
 51 4e 4c 4d 51 4a 46 4f 50 50 44 40 48 4b 49 54 4a 4b 48 4b 4f 49 45 4a 52 52 4c 52 53 57 59 4e 53 4d 48 57 4a 53 4b 4f 54 51 54 56 54 55 58 54 60 5b 5a 5a 60 60 58 5d 62 60 6a 6c 5e 6b 68 69 72 6f 75 71 70 72 74 71 48 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 22 5d 68 6d 5f 62 62 60 63 61 5d 63 64 5a 59 57 54 55 4f 51 52 59 44 58 45 52 48 4e 4a 4c 4b 4b 48 3f 47 4a 45 45 46 46 48 4d 4b 4d 51 50 54 45 4b 45 40 44 3d 3e 2e 35 46 39 3b 33 3f 3f 3d 36 3d 3c 42 41 3b 41 47 3d 49 52 41 4c 50 4a 4f 42 4a 4d 51 46 45 36 32 23 10 05 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 11 17 21 2b 32 35 42 4d 4b 46 44 4b 48 44 3f 4a 4b 44 3d 40 47 49 49 46 42 48 4a 45 45 4a 3d 42 41 40 48 49 50 4a 4c 43 41 42 4f 52 40 4b 43 41 4c 44 49 4c 47 4f 4c 40 50 4b 4d 48 4d 52 4d 4a 4b 4b 47 52 4f 52 50 49 51 4e 47 53 4e 51 59 5b 56 57 55 5a 53 62 59 57 5f 65 60 64 5e 64 62 6a 5f 68 6d 6b 62 5f 6e 70 6f 6e 61 3c 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 21 51 68 72 60 65 60 64 5b 62 62 66 5b 57 56 4f 55 59 56 5a 4b 51 4b 52 50 4c 4a 44 47 46 47 46 3c 47 40 44 49 46 45 4a 59 4e 52 55 4b 4e 49 40 3d 41 47 46 3d 36 36 36 3a 3a 33 3c 36 3a 39 3a 3f 3a 44 41 3a 3e 45 4b 4b 40 4e 47 42 50 50 49 4f 4a 4d 44 3d 36 29 13 19 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 1c 24 2c 2c 3f 42 45 41 4a 45 4c 4d 42 47 3f 4b 44 40 43 4f 47 48 46 46 4b 46 42 44 45 45 42 45 45 4b 48 50 48 42 43 45 4e 4d 43 49 36 42 42 41 4e 49 49 45 4a 45 3e 43 49 46 47 4b 4c 4a 45 48 4e 52 55 55 4c 4b 49 4a 51 4e 4c 50 50 54 57 55 4c 58 5c 50 5b 5a 5c 55 57 5c 61 65 65 6a 64 6e 5d 67 5d 65 66 64 65 69 6b 5e 43 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1d 4f 64 5f 5b 65 64 5b 5a 53 60 5c 55 59 4d 50 4f 54 55 54 4e 4d 4a 59 48 4d 44 4c 44 44 43 52 4a 48 4d 3c 49 4a 4c 54 52 52 4c 50 4f 4a 4a 47 3b 3f 39 3f 3b 3d 3d 3a 3a 35 39 3e 37 3c 38 38 40 35 3f 38 40 3f 4d 46 47 48 4e 44 53 55 50 4f 42 48 41 43 3d 2f 23 16 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 0d 15 1a 27 2e 3d 3d 48 48 44 45 4a 48 3e 45 4d 47 46 4b 41 3f 45 45 47 43 49 41 46 47 46 42 46 44 4a 4a
 4f 45 48 44 4c 43 3d 49 40 45 48 45 41 4a 41 3b 47 45 45 45 47 42 49 3f 4b 4b 50 45 46 4a 46 51 48 4b 4a 4e 47 4f 4e 49 4a 4a 50 52 56 54 58 55 56 58 5b 54 60 56 5c 5f 5d 60 65 5f 5f 65 66 66 5e 63 5b 67 5c 6d 5f 59 47 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1c 58 5e 5f 5d 5d 5c 55 59 59 5f 5c 5b 58 58 55 55 54 4d 53 51 4b 4d 4c 4d 50 4b 43 4b 4a 47 4a 4c 43 3f 4b 49 4f 4d 48 49 49 48 48 4a 4e 4c 42 3a 3d 42 40 41 44 38 3b 46 43 3e 33 34 39 3a 3a 3d 39 40 3e 44 54 45 43 43 4d 4d 54 47 56 4e 44 50 43 4b 3c 39 21 1e 11 05 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 10 17 24 2a 38 3e 3d 4e 48 40 4c 48 45 44 40 4b 42 42 45 4b 46 44 42 43 47 45 44 45 41 45 3b 40 3f 4d 45 45 47 40 43 46 40 4f 45 46 49 45 40 35 48 3f 3f 3d 3f 46 46 3b 42 43 42 47 41 43 3d 4b 55 52 52 50 46 46 59 51 52 47 4d 52 59 55 52 4f 55 54 58 58 56 5a 58 53 5b 5c 5a 5b 60 5b 5f 61 67 66 64 56 5d 58 58 56 5e 58 37 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 4d 5d 5d 5c 5e 5e 53 5c 56 55 5b 55 54 56 4b 48 53 4e 4f 40 56 43 50 45 48 42 43 3d 46 4a 45 47 49 49 46 42 4f 41 41 50 42 40 49 45 46 45 46 4a 3b 3f 39 3f 42 41 3b 39 40 3e 3b 37 37 38 3c 3d 41 3e 40 43 39 49 43 46 4f 4c 49 50 4f 56 4a 48 4b 44 41 32 25 21 0a 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0b 0f 1f 27 40 41 42 4c 3a 48 43 45 41 40 44 40 47 4e 3c 45 41 41 47 3e 45 43 3d 42 46 42 46 48 4a 44 4b 43 3c 41 3d 40 47 3f 49 40 3f 42 3c 40 41 42 47 45 46 38 47 39 3e 45 44 44 45 42 4d 49 50 4f 46 54 53 4d 4d 52 47 46 4a 4d 51 5a 49 50 4f 52 4d 50 53 51 53 52 5c 58 50 5e 5e 5e 63 60 60 5c 58 5e 50 50 58 58 4e 3f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 44 54 5a 5e 5d 56 56 51 5b 52 54 4e 51 4f 4c 4e 4f 52 4b 4c 4c 48 45 47 46 40 45 3c 4e 42 45 47 42 45 46 49 3e 3f 45 43 46 3c 41 3f 44 43 3e 4b 38 41 45 38 41 39 3f 3a 3d 39 38 3a 41 37 39 3c 42 40 45 40 3e 41 46 49 4e 4d 50 44 4d 48 48 4d 44 47 36 2c 20 14 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 07 09 16 1f 29 3a 41 42 47 44 45 40 45 45 42 46 4c 47 3d 46 45 3e 45 46 48 4f 44 46 47 46 3d 42 43 44
 3e 45 45 49 47 46 43 46 44 43 3f 43 45 3b 3d 40 46 47 41 44 3f 42 48 3c 4a 42 46 46 40 47 4d 56 57 4f 51 52 4e 52 49 4b 52 4f 4b 55 53 4a 4c 50 52 4f 53 4f 51 4f 5c 55 55 58 5e 60 61 5e 5e 53 5f 5a 58 5a 52 55 53 53 3f 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 39 56 5c 5a 58 55 48 58 50 5b 56 4e 54 54 4d 51 51 48 51 4a 47 4c 46 47 43 43 44 3f 41 43 45 45 4b 4a 4c 45 39 47 3c 41 47 42 41 3f 48 44 49 41 44 42 3a 40 42 37 44 3c 39 3f 3e 42 3b 3d 44 3f 44 40 42 40 48 40 4c 4e 47 52 49 46 50 55 56 52 46 49 38 24 22 0e 0b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 1f 2a 30 38 42 47 45 47 44 41 3c 3f 4a 42 3c 41 41 43 48 44 41 40 44 41 45 44 48 42 47 46 43 42 46 39 44 41 42 40 42 41 3d 3a 38 3b 46 3e 44 3f 3e 41 40 42 3f 3f 41 40 44 4c 46 3e 41 51 55 51 54 55 4f 50 4c 55 4d 51 50 4c 4f 4a 4f 52 4f 51 4b 4b 4f 4d 51 51 50 4f 5a 5e 5b 57 64 59 5a 56 55 4d 4f 4c 4f 4b 4e 3e 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 37 57 60 56 59 56 55 54 50 4d 4c 4c 54 48 4a 54 50 4d 47 44 4e 43 49 46 3e 44 3f 3d 43 44 43 43 44 44 49 48 46 3d 3e 43 42 3e 3f 42 42 44 47 3e 44 37 3a 3a 3f 39 45 36 3d 3e 39 3c 3d 43 45 43 3e 41 45 44 42 49 4f 49 4b 4c 4f 4c 4c 52 50 56 4a 3b 31 1d 12 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 11 28 2a 36 38 3d 41 47 47 42 47 3d 40 4b 3d 3d 46 45 44 3f 41 3a 3a 48 47 3d 4a 42 43 41 45 44 40 3a 3e 41 42 34 44 3d 51 3a 38 42 4a 3e 3b 38 3f 3a 43 43 3a 3e 3c 41 41 49 33 45 46 52 55 4b 4c 4b 57 49 4a 4b 4f 56 4f 4b 52 4c 54 47 51 52 4b 49 4f 45 51 4c 51 56 52 55 59 5b 55 59 57 53 51 4c 4d 49 46 52 4b 35 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 35 54 56 46 57 4b 49 51 51 4e 4e 44 49 4d 4c 50 49 4d 50 49 42 3d 48 3f 47 4c 46 4a 48 4d 46 55 43 47 4c 45 43 41 40 40 3f 47 46 36 38 3e 38 42 36 43 40 3c 41 45 42 3a 37 34 3e 3a 3e 43 3f 42 42 42 45 3d 42 44 44 4b 4a 49 50 43 50 52 52 4f 3e 3e 33 17 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 1c 1a 26 30 3d 3e 44 47 46 47 43 3f 4a 4a 46 42 47 41 45 48 40 44 41 43 42 42 47 39 3a 3c 44
 3f 44 42 41 41 44 40 4e 40 3e 49 44 3a 3d 40 45 40 43 3a 49 40 47 3e 35 40 3e 3e 43 43 48 4e 4f 4d 4a 43 4c 42 4c 52 4d 4f 4a 4d 4e 48 4f 49 4d 4c 4d 50 53 48 56 4c 4b 4d 4d 58 52 59 4f 53 4f 4e 4c 54 4c 55 4f 47 4b 3d 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 3f 4b 50 4c 52 4f 48 4c 4a 4b 51 47 46 47 4c 4d 49 40 4c 47 50 42 45 47 46 47 4f 4c 49 4d 4a 49 46 44 45 3f 3e 3e 46 3e 3f 44 45 3f 41 45 3d 3f 34 43 3c 37 38 3a 43 42 3e 42 42 3e 3e 44 3e 40 48 48 48 40 44 44 4a 40 46 49 47 49 50 4c 4d 4e 3b 30 27 18 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 12 10 23 30 36 34 42 4d 47 42 45 42 40 40 49 4a 40 48 48 3d 3f 3c 45 42 4b 3f 42 3f 3d 44 3d 40 46 42 40 3f 39 3a 48 40 47 3f 43 3c 40 43 3c 45 3e 3a 3e 3a 41 40 3f 40 39 38 46 48 46 4d 46 4a 4d 4a 4e 4d 44 47 4b 53 4c 4e 4f 42 4b 48 46 51 4b 4b 4c 3f 4e 50 51 41 4f 55 4f 54 4e 4d 4f 46 50 4e 4a 48 4b 4f 4b 38 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 2b 44 50 4b 50 4b 47 45 4e 42 4d 4a 4e 4a 4a 51 4a 47 4c 49 45 41 49 4d 52 53 51 4e 50 4c 47 43 46 45 45 41 3e 3d 3d 3e 41 40 41 3d 3b 46 43 41 3e 43 3b 3b 40 3d 3c 46 3c 3e 3c 41 44 3a 44 45 41 45 41 45 42 47 45 45 4f 4a 4d 40 44 4f 4d 41 3f 31 25 0a 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0b 18 1b 29 35 37 45 41 3d 44 40 3f 4a 3f 47 37 39 45 3d 4d 45 43 3c 3f 3d 3c 41 39 3e 3d 44 39 48 39 44 3a 36 3b 3d 3c 3e 43 39 3f 3a 34 47 3d 40 41 44 38 40 3d 40 3d 3e 34 47 3a 3e 43 46 42 42 4c 49 53 42 47 4e 4b 4c 44 42 41 45 4a 44 4f 45 4c 48 45 4d 45 46 49 4b 53 50 4d 46 4a 4e 4d 4e 4c 4a 49 48 53 3d 3a 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 2f 3e 56 45 4b 44 42 49 45 47 4b 4a 43 4a 43 45 44 41 4f 49 49 4b 49 57 50 55 54 50 4d 4b 44 43 40 41 4c 44 3e 44 49 3a 3d 44 45 40 41 42 3d 3e 3c 47 40 3c 3c 3a 42 3f 42 49 46 3e 41 4e 43 48 45 44 45 38 41 42 40 47 43 3b 4a 3b 43 4e 48 43 35 27 22 11 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 13 1c 27 33 33 3f 45 3c 45 40 3f 47 42 4c 38 42 41 40 47 46 3d 39 48 3e 3a 3e 3b 4a 42 49
 37 3d 3c 41 44 41 38 40 45 3f 47 40 3d 41 43 41 41 3a 3a 40 42 3e 3b 46 43 3b 3c 37 3c 3e 44 39 43 46 41 4a 40 46 4a 50 51 46 47 3f 48 45 44 48 4f 4b 4d 4c 47 51 4e 46 4a 51 4d 49 49 50 54 51 45 49 4a 4b 4d 4a 4a 4a 3d 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 2d 43 49 47 4c 4a 49 49 46 4e 4a 4f 49 43 4b 43 46 44 46 44 49 4c 59 57 59 54 4f 55 4f 41 46 43 3c 44 46 41 3b 42 44 4e 49 44 42 41 3e 49 4c 44 3f 39 42 41 3e 3d 45 42 40 46 3d 3e 46 47 3c 42 4b 3b 47 45 4c 44 46 47 4c 42 4a 44 47 4d 44 3f 34 26 1f 0c 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 1a 21 31 3b 39 41 3f 41 44 45 40 34 38 40 44 40 43 38 40 3e 45 3c 4a 3f 44 44 44 42 3a 41 43 3c 40 45 3d 37 42 3a 39 3c 40 41 37 3f 40 3e 3b 44 38 3b 40 42 40 3f 3d 3a 37 32 2f 3d 3f 49 44 3e 41 44 49 52 4b 4c 47 4b 4a 46 46 47 47 4e 44 4c 52 4a 4b 4a 4b 47 49 4d 54 4a 4d 4c 47 4c 44 41 44 47 42 40 4a 33 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 24 41 47 49 49 4f 40 45 46 3f 51 49 44 42 4c 46 46 44 45 49 4d 4c 52 58 5d 53 4b 51 4c 44 48 40 44 42 4a 42 45 3b 48 47 3b 3f 45 43 37 3f 42 3c 3d 48 46 42 3c 3f 45 3e 3e 49 40 38 39 47 44 45 3e 43 49 3a 47 42 43 46 4f 48 4f 40 46 39 38 3e 25 19 0e 08 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0d 12 10 25 30 3e 3d 3a 3e 45 45 3b 45 43 42 3a 47 44 3c 3d 44 47 40 3e 46 49 3d 3f 3e 38 3d 3b 3e 40 3a 3b 42 3a 45 41 3e 3d 40 40 3a 41 41 41 41 3d 34 43 43 3f 4a 45 37 34 35 39 3f 48 47 36 3f 46 47 3d 44 46 44 4c 4b 46 48 47 3c 4a 4e 49 4a 49 4d 4b 48 4e 42 4d 43 48 49 4b 46 49 44 49 45 45 47 46 44 44 2f 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 20 3d 3d 46 47 44 45 45 43 4b 40 49 4a 46 44 45 43 46 43 4f 4b 51 5c 5b 5d 51 50 4b 3b 49 43 39 3f 40 3e 3b 42 40 3f 40 3f 41 41 43 46 45 38 43 44 45 3b 42 4a 3a 4d 48 45 44 4c 45 41 43 3f 46 40 43 44 3e 46 48 49 44 44 43 44 4a 3d 42 35 2e 21 17 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 12 28 2d 37 40 37 3b 42 3c 44 40 40 46 3d 3e 36 3d 3d 40 45 48 42 43 43 48 3e 44 44
 3c 42 48 35 3d 39 3e 43 41 3a 44 43 45 40 3c 3f 3d 3f 40 42 39 3c 41 3b 42 3b 3b 35 3a 38 48 32 20 2f 49 47 41 3f 3d 44 46 4c 48 42 3e 41 40 46 4f 49 50 48 43 43 48 43 4e 46 45 46 4b 50 41 44 4c 45 45 45 40 48 3a 46 37 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 1c 42 49 47 40 49 43 42 44 41 48 41 47 4c 47 3b 4c 51 47 4c 55 54 55 4e 53 55 47 44 45 3c 3c 45 3d 48 40 3b 34 37 43 48 3d 3d 48 41 43 49 44 46 47 45 43 42 41 42 4d 40 44 47 47 49 42 42 3f 3d 3e 4b 45 47 46 4a 51 45 3e 49 48 45 43 3e 33 2a 1c 15 0e 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 0f 1e 27 33 3b 42 3d 44 3b 3e 43 42 42 45 3d 43 41 44 43 42 43 45 40 41 45 41 42 3e 3d 40 3f 40 40 40 40 41 3f 41 47 3d 48 3e 35 3f 41 36 42 3b 42 41 3d 36 44 3a 39 43 39 42 3d 3c 41 43 47 40 3c 41 42 42 4a 44 45 49 42 44 45 40 44 44 44 4b 50 4f 4a 51 47 4d 4b 49 42 49 44 48 44 44 48 46 3e 40 43 3c 3b 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 39 44 3f 47 47 39 44 43 40 47 44 4d 4b 42 46 41 46 45 4d 55 5c 51 53 52 4b 43 40 47 4c 45 3b 41 46 43 40 42 48 4b 45 44 46 3e 3a 49 48 44 3f 45 3b 4f 3f 41 48 51 3e 47 48 45 4a 43 49 45 3e 43 3e 4f 3e 4a 3a 4d 45 49 53 4e 48 45 3f 28 23 1b 13 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 19 21 2c 3f 44 3d 45 41 37 40 3d 41 41 43 44 42 3c 42 3e 42 35 42 43 3f 46 3b 40 3d 3a 3d 39 3d 47 3b 3e 3f 3b 39 37 41 47 3a 3b 40 3e 3f 3b 3d 42 3a 3f 42 45 3a 41 3e 39 48 42 3d 36 3b 42 35 3c 40 39 47 49 48 49 41 47 44 49 51 4d 49 44 4a 4a 43 4d 41 44 44 41 48 4c 3c 47 46 44 47 3e 37 41 38 3b 30 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 13 3a 4d 3d 45 3e 42 3e 45 3f 49 3d 48 42 43 47 49 4e 50 4f 5a 4d 54 50 4b 45 43 38 3f 3e 44 41 3d 45 3c 40 3e 40 3e 46 4c 3e 44 37 45 49 48 44 45 44 46 42 3f 42 4b 3d 43 3f 43 3e 48 3c 4a 3b 45 45 40 41 46 44 45 45 4b 4e 50 41 3c 32 27 1e 0d 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 06 05 03 12 16 29 38 3c 45 40 3c 37 41 3b 41 3b 40 39 35 40 41 47 41 46 41 3f 41 39 46 44
 3a 3f 48 3a 42 3c 40 3d 3c 40 3e 3d 37 43 41 41 3a 3c 3d 45 35 3c 35 38 3f 45 39 35 3f 36 3f 41 41 3a 3b 42 3b 39 3b 3d 3a 44 4e 4c 46 44 3e 44 4b 50 4a 4b 46 4b 43 48 4a 44 47 4c 48 45 4a 40 40 3d 35 44 40 37 4d 39 35 26 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 39 42 3d 45 43 45 41 42 3b 3f 47 48 46 44 4a 4f 52 4e 4f 51 4d 4b 4a 45 3d 43 42 46 43 42 41 42 42 3f 3b 3f 42 43 3e 4a 4a 45 41 46 40 42 45 4d 43 46 4f 49 4d 43 46 49 45 45 3d 38 45 48 44 44 48 45 3a 46 42 45 49 4f 51 52 48 34 2d 1e 1c 0f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 10 17 20 35 3b 45 3e 40 43 3a 37 3f 3b 3c 3c 39 43 3e 46 3c 47 45 43 46 3f 45 45 42 3c 45 3e 3e 3c 40 46 40 3c 3f 45 3e 40 3c 42 3e 43 3a 40 3e 3b 3d 40 3e 32 3e 43 3d 3e 40 3f 41 3e 4a 42 39 45 3f 49 4d 40 46 46 44 44 4e 44 40 41 4b 4e 50 4e 4c 47 49 45 46 49 3d 43 46 43 41 45 3a 41 41 3d 3e 42 35 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 16 2f 42 41 49 3b 4b 40 42 42 54 42 43 49 4b 44 4d 4d 4f 51 57 55 54 44 49 4a 41 45 40 3f 41 42 45 3f 41 43 3a 47 46 49 55 4b 47 47 4b 40 49 4d 4a 59 4f 49 4c 47 48 3e 47 47 44 41 42 47 43 4d 4a 4e 4b 41 49 3f 48 45 4d 47 44 3d 39 2c 24 18 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 10 1c 2b 34 36 42 35 3e 44 3e 42 3d 43 39 42 3c 43 3f 45 45 4a 48 45 48 41 4b 48 3e 3d 40 3e 43 43 44 39 42 44 41 3f 3e 3b 3b 40 39 47 41 3e 41 3e 3d 3d 42 43 4b 39 33 3b 3b 41 41 3f 40 3c 3c 3e 40 4d 3e 3b 41 43 4b 48 4c 45 4a 4b 45 41 41 41 3c 40 45 4d 51 48 48 3c 45 42 41 35 44 42 42 47 41 34 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 2c 40 42 4d 40 40 41 3f 42 46 46 47 42 50 46 4a 4f 52 4e 55 4f 49 3f 46 38 44 4a 45 48 44 3b 49 41 3e 48 4a 52 59 5e 5a 52 57 54 4e 57 52 4a 51 55 5a 49 48 43 4d 47 49 4a 45 3e 41 3d 42 44 44 45 50 44 46 48 41 4e 49 40 46 33 2f 24 1f 15 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 09 18 22 2d 40 4b 3e 44 38 3b 3d 3b 3e 40 41 38 47 41 50 41 44 46 44 43 40 41
 42 44 46 39 44 40 3e 3f 42 3e 41 41 39 3d 3b 3d 4c 3f 39 45 3f 3e 45 3f 4a 3a 38 3d 3c 3a 39 3a 46 3a 3e 42 45 3a 3e 46 44 39 49 3c 3c 46 3e 4b 45 3e 44 49 4c 44 44 42 4a 40 40 46 48 46 3d 45 42 47 44 3e 38 31 37 39 36 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 32 47 3e 4f 4d 47 40 45 45 45 50 49 4a 47 48 55 49 4e 4b 4b 49 48 46 44 46 3d 47 40 39 41 3f 49 4c 4b 40 50 65 5c 64 60 56 64 60 56 61 55 62 62 64 64 55 5d 55 55 56 58 5a 4a 41 41 39 3c 42 4c 3c 46 44 45 43 41 3e 42 4c 3f 35 26 25 14 0c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 0a 1c 2f 30 3e 42 48 39 40 3c 48 37 38 41 3e 4b 49 50 4b 47 45 42 42 42 3e 48 4b 44 49 46 46 43 42 3d 3e 43 3d 3c 44 3d 40 3c 39 43 46 3e 47 4a 42 42 3c 3f 3d 42 39 3b 3b 3f 3a 3b 3f 3f 3e 3f 43 41 3b 42 46 42 42 43 4d 44 48 41 46 40 50 42 40 3d 45 44 49 4b 48 45 46 3e 39 3c 42 45 3b 3d 3b 2d 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 14 32 44 40 42 41 43 49 4a 4a 42 46 4f 49 4d 44 54 50 59 44 45 4b 48 42 49 48 4a 46 3e 45 44 45 4c 47 55 52 67 62 6c 73 6f 72 71 7a 70 6f 72 7a 73 79 6f 69 70 62 6c 65 5f 66 52 3f 3d 3d 49 47 46 43 42 3c 48 44 46 48 41 3f 3c 2f 25 25 14 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 17 1e 29 3e 42 42 3f 37 43 41 3d 3f 3c 49 4a 4e 4d 43 49 41 40 40 48 3d 3d 50 47 47 4c 4a 45 44 47 43 40 47 45 42 3c 43 3e 38 3b 3b 38 42 3e 45 3e 3b 44 3f 3d 3e 37 3c 44 43 45 44 49 3a 3a 3d 3c 3b 46 3d 42 3c 41 41 3f 43 45 43 41 46 3a 43 3f 3e 42 44 45 43 46 47 43 41 3f 38 3a 3e 45 41 37 25 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 33 4a 45 46 44 43 49 3f 45 48 46 4f 4c 4e 44 50 4b 50 4a 41 4a 44 42 42 41 48 3d 4e 44 4e 4a 50 55 57 65 6b 6a 76 7a 7c 7e 83 7a 77 85 83 84 86 80 7b 7c 7c 79 75 73 69 60 63 53 58 3f 41 3e 3e 39 47 40 3c 41 44 52 40 3d 3e 2a 1b 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 11 1a 1d 34 3b 42 43 42 38 45 38 3d 3e 4c 4c 49 51 44 47 44 42 41 3d 45
 4f 4b 44 47 45 50 48 45 3d 3b 44 46 38 3a 40 48 3b 42 3f 45 38 42 40 3f 42 3b 3f 44 3f 3b 3a 3e 3d 42 3d 40 3c 3a 3f 40 3c 3c 42 3d 3b 39 3d 44 42 3c 41 40 3e 41 4a 3f 3f 3f 45 48 44 4c 3a 45 3e 43 44 3e 37 3d 37 3c 3a 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 31 43 44 40 3f 42 40 4c 40 54 3f 4b 4b 46 49 47 47 45 44 4b 44 41 45 48 42 40 3f 42 4f 48 4e 54 5e 64 76 76 7d 87 83 80 81 83 85 80 85 84 85 80 7b 7c 79 86 80 80 85 7e 79 76 61 52 41 3d 3c 3f 3c 41 44 46 44 51 4c 3f 3a 28 24 1d 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 12 1d 2b 3f 43 44 44 41 43 3a 3d 42 49 4b 4d 47 42 44 42 3f 41 44 4f 48 49 49 43 41 4b 45 43 44 46 42 39 36 43 44 45 44 38 3f 4a 40 3b 45 3d 3e 43 41 46 40 40 3c 47 42 42 3a 3a 40 3e 3f 42 40 3b 41 3d 3b 45 35 45 42 3a 3a 44 44 45 46 3e 36 42 3c 47 43 49 48 45 47 4a 41 43 3c 42 40 3b 34 27 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 33 49 40 3d 42 3f 44 4a 48 4a 46 4c 44 49 49 4a 50 42 44 4a 49 4c 47 57 41 46 4b 4f 59 5e 60 67 78 78 80 87 8c 8b 8d 8d 80 89 85 87 8c 87 86 8a 87 8b 84 81 81 89 88 7a 7d 79 6e 6c 53 4a 44 42 3b 4b 43 45 51 48 3e 44 35 32 1c 1a 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0c 0c 12 26 2c 41 41 46 3d 3b 41 41 3b 3e 47 4c 3f 46 43 3f 42 3d 3c 4b 53 5a 48 47 48 4a 44 41 41 45 3b 44 44 42 45 44 45 42 42 45 3b 44 44 3d 41 3e 3e 45 43 4a 48 43 41 41 43 3b 3c 3b 3d 43 40 39 40 44 3e 47 38 43 41 3c 3c 3e 34 48 3c 43 3a 42 42 44 4d 44 3d 38 40 3d 43 41 40 43 3b 43 3d 2e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 2d 3f 40 41 47 45 3e 44 40 4a 46 4b 4d 47 48 45 4a 4d 44 44 4e 49 49 54 50 54 54 62 65 77 72 84 88 83 87 87 85 8b 88 8b 8d 84 85 84 8a 87 7e 83 84 84 85 84 82 7f 87 82 82 7c 73 78 66 4e 49 40 35 43 42 4b 4b 52 46 37 35 2a 16 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 13 20 2c 38 48 45 41 41 3a 3f 33 39 3a 42 3f 3a 3e 44 46 41 41 3f
 3e 4e 46 46 41 46 43 44 43 48 41 3f 41 41 40 3d 3c 3b 47 46 3f 42 41 3c 39 3c 35 3e 3b 41 3b 3f 3f 3d 3c 3f 3b 44 3f 45 3d 3a 3c 3e 39 3e 3c 3f 3c 37 3d 39 3d 3a 36 39 3b 3d 47 40 45 49 49 3d 42 3b 4b 38 3c 3f 3f 36 32 2b 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 21 41 38 43 3f 45 43 41 47 49 50 4c 46 4c 4c 48 45 45 41 45 48 48 52 58 50 69 6b 72 79 84 85 88 8a 89 84 85 8b 82 86 82 87 84 83 80 7a 8e 7d 7a 81 84 7c 7f 80 85 8a 84 80 77 77 6c 69 58 46 41 39 3c 38 42 47 45 3d 2f 27 26 12 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0b 0d 24 2f 47 40 40 43 41 3d 44 38 3b 40 3f 3d 45 46 3d 3e 3e 36 42 48 40 41 3f 46 4b 41 44 38 3e 3c 3b 3f 40 3d 3f 3d 46 41 43 3f 41 3c 3f 3d 44 3f 3e 40 44 39 43 44 42 45 36 3f 41 43 41 41 45 41 37 3d 45 40 49 3b 41 42 40 3a 38 33 3a 48 45 45 4a 46 42 44 3e 3b 47 42 45 49 41 3f 32 2e 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 30 3f 3d 3f 4f 44 46 4c 4e 4a 4b 45 46 4e 45 45 46 46 46 4c 48 51 56 62 73 70 83 83 8f 90 84 89 84 8c 7e 80 85 83 85 7f 85 85 89 84 7e 7f 7d 79 7b 7d 7c 87 83 85 80 78 82 7a 73 75 69 58 52 4c 40 42 3b 41 47 41 38 34 22 20 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 1b 29 39 54 4a 49 44 39 36 3d 3b 45 3b 3a 46 3e 45 46 3b 3f 3f 49 3f 4a 42 46 45 46 46 4b 37 3c 3b 40 45 48 45 41 42 3e 3c 45 3c 3d 43 3e 47 3f 3d 39 3e 46 40 41 4a 3e 45 3d 3b 3d 40 4a 40 44 3a 3b 43 3d 40 46 3c 40 3f 46 3d 3e 3b 35 44 3d 41 47 43 4b 46 47 44 42 3f 45 3c 41 30 2d 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 2f 3d 3e 48 3e 44 46 4b 48 43 3b 4c 42 4a 49 4f 4e 52 4f 58 5b 6a 6d 80 84 86 8f 8c 8e 88 8d 8e 83 84 85 86 8b 81 7c 82 7d 7d 7b 76 7c 7c 7b 76 76 7d 74 7a 81 7e 7b 79 7f 7c 7b 7c 6c 5e 4e 54 48 43 3d 40 3b 38 31 27 19 11 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 11 1b 2d 32 38 40 3f 43 36 3b 33 38 40 39 3d 37 3e 36 35 3d 3e
 47 41 48 41 44 47 3e 43 3c 37 42 44 3d 3c 3d 40 4d 3b 49 42 44 3a 3d 45 3f 44 44 3d 3a 3b 3b 3c 41 39 3e 41 3d 3d 3e 3d 40 49 49 42 3e 39 39 3c 39 36 3d 3c 3d 44 37 36 36 39 34 49 45 43 3d 44 47 48 47 44 4a 40 38 40 3f 2f 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 2d 44 49 4a 41 46 45 46 3e 49 49 41 4a 48 4e 50 4b 53 56 6c 7b 7c 8a 8d 8a 87 8a 8d 89 8f 80 7c 85 84 80 7b 83 81 82 73 7d 7a 73 78 78 74 75 7d 74 76 78 77 73 80 77 82 80 78 7d 78 69 62 4a 49 45 3d 3c 42 40 3b 2c 24 0d 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0f 19 27 2d 41 4b 42 40 35 3c 3f 40 37 3b 43 3d 45 42 3b 3a 43 3d 46 42 3d 41 43 3e 3b 47 3f 37 3f 42 40 41 43 45 48 41 3b 47 43 44 45 3b 44 46 3a 3d 47 40 44 41 43 41 41 3e 4a 46 3f 40 43 3b 43 42 3e 44 3d 42 42 3c 41 45 3c 3f 40 3e 3f 46 42 44 4c 45 4c 4a 45 41 3d 44 49 3d 3a 2a 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 25 38 3b 4a 43 40 43 42 44 48 4d 52 48 54 56 56 62 69 76 84 86 8f 8f 94 8d 8c 8b 90 8b 85 7b 84 80 7b 80 7a 85 80 7e 7e 70 74 75 6f 75 79 76 73 76 71 78 7e 7b 80 78 73 84 82 7c 71 67 5f 63 4f 44 3b 3f 3f 3d 35 24 1d 12 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0d 13 1d 24 32 3f 39 38 36 3a 39 39 40 41 39 3c 3b 3e 3e 3e 41 43 3c 43 3c 45 3d 42 3b 46 44 3b 3f 43 3b 4a 3c 3c 40 50 39 3a 4a 42 46 4e 3b 4a 42 41 3a 41 4a 3d 4a 44 3d 3f 3e 43 46 42 45 3f 3b 3e 3d 47 3c 40 44 37 40 42 3d 38 3d 3d 3f 4a 3f 50 49 45 48 47 45 3e 3e 36 42 39 3c 29 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 24 3d 40 44 4c 44 45 44 47 49 4c 52 5c 64 65 6c 73 83 82 92 8d 92 92 8f 90 8a 91 8f 87 8b 7e 7d 82 7d 75 6f 78 74 73 73 71 6c 7b 75 74 75 71 6c 75 76 65 7e 78 7b 7f 73 78 7d 73 70 6c 65 5e 4f 49 3d 41 38 32 26 1d 16 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 10 24 35 2f 44 3e 43 3b 36 40 39 3c 36 35 35 3d 41 3f
 43 39 38 38 41 42 3f 39 41 41 41 40 3e 41 45 44 41 41 3f 44 39 4c 42 43 3f 45 46 42 42 3e 47 42 3a 43 40 41 4a 41 3e 44 41 43 42 49 40 3c 43 44 42 39 3d 40 3b 3c 3d 3e 3e 38 3d 41 3f 47 42 46 49 45 44 44 46 3e 42 3a 34 2f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 24 42 41 45 52 43 46 50 49 54 5f 62 79 77 7b 84 89 8f 83 8d 93 95 86 90 87 83 86 7f 7f 7e 78 77 76 77 79 72 73 78 71 79 75 72 6c 75 78 73 77 6e 6e 75 70 72 79 7b 7a 74 7d 74 70 75 6c 62 57 4d 4d 40 39 35 2d 1c 19 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 0b 1c 28 37 3a 44 3c 42 3e 3e 3e 41 41 43 3f 3b 37 3c 3f 41 3c 31 37 3b 3b 3f 3f 3e 41 38 3f 3b 43 44 3e 41 38 48 3e 4b 41 3d 3d 3e 3a 42 3d 43 39 43 41 3d 43 40 45 44 44 45 44 39 4a 3c 45 49 44 43 42 3f 3a 40 3e 35 3d 3a 43 41 3f 40 3e 40 44 42 45 43 52 4c 45 3d 3e 3a 3a 27 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 24 44 3b 44 49 52 58 59 5e 71 70 79 7b 84 8b 8f 87 90 8e 90 88 8e 87 88 83 84 82 81 7d 82 75 73 7c 75 74 6d 75 6d 6d 6e 6d 71 6a 6a 71 70 75 6b 6f 74 70 6d 71 75 76 71 7a 72 6f 70 68 5e 61 53 47 3f 3a 31 2a 14 09 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0e 18 20 28 37 41 43 45 46 41 41 44 48 40 3b 3b 41 3c 3b 39 41 3f 36 36 3a 3c 3f 40 3d 3f 45 3a 3b 42 46 3d 42 41 44 42 44 42 3f 46 3e 46 3f 3f 42 43 48 3e 3f 45 47 3e 41 43 47 48 43 3f 4a 3e 38 45 44 45 3c 41 42 3e 37 3c 43 3f 40 42 3b 44 40 3e 46 48 43 41 3a 41 37 3b 3d 2f 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 1d 49 44 4f 51 5b 69 74 73 80 7d 80 8e 91 99 8a 94 92 88 88 84 8d 8a 88 82 7c 7a 79 7b 7c 73 6f 79 74 69 70 69 6f 72 6e 72 6b 66 70 6a 78 6f 70 69 6e 6b 71 76 77 79 7d 72 74 6c 70 68 64 4f 4d 40 3d 33 32 1d 15 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 09 11 20 1b 2a 3b 3f 4b 49 45 43 4e 46 3e 47 3a 38 3f
 42 38 3c 40 37 3a 3f 3b 43 43 43 40 41 3a 39 43 47 43 3f 47 42 46 3e 3c 4d 46 48 42 3c 46 42 3f 44 45 3e 44 3d 44 3e 44 4a 39 3a 3c 3b 3c 3c 44 39 44 3f 3c 47 39 42 4a 41 43 3c 3f 45 44 42 41 44 4b 47 45 44 37 42 3c 34 30 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 23 4b 5d 65 75 76 77 84 82 89 83 88 8a 8e 91 8a 91 85 89 8c 84 82 7f 84 7f 75 7b 73 74 72 6b 69 67 69 72 71 68 70 6c 65 6b 67 6d 6f 6e 73 69 71 6b 69 69 70 6a 74 70 6d 73 69 6c 67 63 56 4e 43 39 2f 25 18 1a 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0e 1e 2a 2c 36 40 49 4f 4f 46 3c 46 34 34 3e 30 3b 38 36 37 3d 32 3d 3e 38 40 3e 45 39 44 42 44 3c 43 48 41 41 44 48 42 47 45 3d 44 3f 43 42 44 42 3f 42 43 41 40 40 41 42 3d 48 41 41 4a 40 43 3b 3e 39 3d 40 42 3f 40 43 3c 43 45 3d 3f 44 40 49 3e 43 39 3e 3b 39 39 2d 34 1c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 21 52 69 74 83 84 81 83 8a 84 8b 8c 93 89 86 87 81 84 88 87 7b 79 7a 7a 75 73 73 79 71 6a 6d 69 73 6b 69 64 6a 6f 6b 69 72 70 6c 60 69 65 64 6f 70 70 6f 6f 6d 77 6d 70 6c 67 66 67 5b 51 4a 44 35 2d 15 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 11 22 27 30 36 4a 4c 49 4c 42 44 3f 3d 35 38 37 3e 3c 3d 3c 3c 3e 3d 3c 40 44 47 3e 4f 43 48 43 3c 4a 45 3c 46 43 42 4d 42 47 4f 3a 43 48 42 48 48 43 3d 40 38 47 42 41 41 42 3d 38 48 46 40 48 44 3e 45 36 41 43 39 3e 45 4b 40 41 4a 49 46 49 4b 4a 46 44 3a 3e 3f 38 38 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 31 6b 72 84 87 82 87 82 92 90 8c 86 7d 7e 88 7d 85 84 7a 7b 72 75 78 7a 7b 73 71 6f 6e 6d 6d 67 69 64 65 67 73 6b 71 66 66 68 66 69 6e 69 67 6d 6e 65 6d 67 6b 6b 6b 69 6c 6e 63 65 57 49 42 41 34 28 13 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 12 1c 22 27 2c 39 3e 53 44 40 40 37 2f 33 3e
 35 3f 30 36 36 3d 34 40 3f 3b 40 41 46 49 47 3c 3d 42 3b 3f 44 42 46 41 43 40 3e 46 44 47 49 47 3c 47 45 44 3c 42 44 3f 41 3a 44 3c 40 44 40 3d 42 3e 3e 44 41 43 40 3b 42 3b 44 3c 3c 46 48 49 4b 45 3e 45 40 3b 40 39 37 2f 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 2a 75 7c 87 88 84 88 83 85 7e 86 82 7d 7e 7d 82 77 74 72 76 73 78 7d 69 71 6d 76 6d 68 6e 62 6b 69 60 64 6f 68 70 69 63 68 6f 66 66 69 6c 69 6d 65 6d 65 60 6a 67 70 69 6a 5e 5e 5d 4e 3f 40 2e 26 18 15 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 12 1b 1f 2b 29 37 48 43 3f 40 37 3e 36 2f 3a 39 3b 3a 37 43 36 3b 3e 3b 3a 3d 41 45 3c 35 39 38 37 43 41 42 47 35 42 41 44 44 43 43 42 48 46 43 4a 44 3e 42 47 40 42 45 4b 43 3f 3e 43 43 3b 3f 40 44 45 47 44 3b 41 3b 41 45 4a 41 48 47 49 46 43 37 40 33 3a 3d 3d 33 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 28 6f 7e 8a 8a 81 79 80 87 7f 82 79 75 7d 73 7e 72 77 71 6f 76 73 72 74 65 6b 68 64 61 6b 6b 67 64 64 6a 68 68 64 66 66 62 69 65 61 66 63 68 66 69 6c 63 62 61 68 6a 6a 67 60 54 4a 4b 39 32 30 1b 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0f 14 12 21 2e 2d 39 45 40 45 3a 38 3b 35 41 3d 39 38 38 42 41 3f 3a 3c 39 3e 3e 47 3f 39 41 38 41 41 3d 42 41 40 44 4c 3b 45 48 41 48 46 43 42 42 49 40 3d 40 41 42 40 39 3b 4b 3f 45 48 4a 42 41 3f 44 44 43 3a 40 38 4c 47 49 45 44 48 42 47 43 3e 35 39 3b 33 32 2f 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 25 69 76 7e 80 73 78 7a 78 7c 78 78 7f 73 74 75 6d 73 70 6c 77 6b 74 6f 68 6b 71 6d 73 6f 6c 62 6d 6c 69 61 66 63 68 67 63 65 67 62 6d 64 66 62 6a 64 65 5f 61 66 6a 5f 63 59 52 4e 3f 35 33 2a 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 12 15 20 2b 30 37 3c 41 3e 43 42 35 43
 3a 43 32 34 35 46 3d 44 3d 43 33 3b 37 41 42 37 3f 41 3b 49 44 3b 40 40 44 3c 43 44 3f 48 45 50 54 4a 4f 4c 41 4f 45 48 45 43 3c 45 4c 45 3a 3d 46 41 45 45 40 42 41 35 42 36 3e 42 44 4c 49 44 3c 44 41 3f 3b 35 31 30 36 32 18 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 21 69 71 7c 7e 7b 7a 73 78 7a 73 72 70 70 72 75 72 7c 6b 74 6b 67 63 6f 63 61 67 65 6a 64 68 67 6f 6a 68 65 65 68 5d 61 67 46 6e 67 5d 6a 60 60 5f 6a 62 64 64 64 5f 5e 5d 54 42 3f 35 30 2a 1f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 06 0f 17 1e 25 23 32 3a 44 41 3a 37 37 3c 32 30 38 36 3d 38 35 3d 3c 3b 44 3b 38 3e 39 44 43 3c 42 47 3f 40 35 3e 3e 44 46 40 42 46 43 4a 4a 4d 53 4d 44 3d 42 43 45 3d 40 43 3e 41 49 4a 47 3a 45 3d 3f 3e 34 3a 45 43 47 42 3d 40 3e 3e 39 3d 3b 3a 30 2f 2e 2e 30 1b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 22 57 67 71 78 68 6e 6d 73 74 6e 70 70 74 73 6e 6d 65 68 6b 6a 65 69 67 68 6b 5c 67 65 68 62 63 6a 60 65 6e 61 62 69 60 66 6a 5b 5e 61 5f 57 60 59 61 65 61 5d 64 5e 57 56 53 40 3a 30 25 17 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 09 1b 1f 31 32 32 37 41 3d 3f 3a 35 36 3a 35 35 44 3a 40 38 41 3d 3d 36 3e 39 3e 42 45 3d 3c 3f 45 42 3f 39 3f 41 3b 43 46 4a 44 47 4e 51 55 4e 4c 4c 44 41 42 36 47 46 40 42 45 4a 42 43 46 47 44 3d 41 37 3b 3b 3c 39 41 3d 3e 37 32 34 3e 32 31 3c 3b 37 2e 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 58 67 66 75 65 72 6a 64 70 6a 6e 71 6b 6d 67 6e 6c 68 6e 64 6e 60 68 5e 62 63 67 62 6a 6c 68 6b 66 61 64 68 5f 62 5a 65 62 59 61 5d 67 65 5b 65 5e 5f 68 5c 5a 53 4a 43 40 39 2b 21 1a 18 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0d 17 26 27 2f 30 3c 42 3c 43 39
 38 3b 39 36 36 3e 36 3b 3a 3e 3a 43 41 3a 39 3b 3e 3c 3b 43 3b 3f 43 40 46 3a 3d 3e 41 49 4e 4b 49 4f 51 5d 50 4d 47 4b 41 3d 40 45 49 4d 40 48 49 47 41 4b 48 3d 42 42 3c 38 46 39 3f 41 3f 37 39 38 2f 33 2d 3c 35 38 27 36 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 10 5a 67 66 6f 62 66 6a 67 65 6b 6c 64 67 67 66 69 6c 67 67 65 68 63 64 69 58 66 6d 68 66 64 66 66 60 6b 65 61 5f 5b 60 5e 67 61 65 62 58 5f 61 5e 5c 5c 5d 57 4f 52 3e 38 34 29 2b 23 15 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 20 20 32 2d 32 35 35 35 3b 35 3f 36 3f 3b 35 40 42 3e 38 42 35 36 3b 3c 38 39 3b 47 39 3d 42 35 3e 39 3e 39 3e 3a 3c 45 4e 46 49 55 4e 4c 50 4a 47 3b 47 3e 40 4a 40 4e 49 49 3e 42 42 41 3e 3b 41 3a 3b 3b 3c 3b 39 44 36 36 2f 38 36 35 35 3a 31 2f 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 12 4b 5d 68 6d 64 5b 63 62 64 65 64 62 60 69 62 61 66 6a 66 66 64 64 61 5b 64 5e 60 63 5b 66 66 62 63 5c 5e 64 64 62 5e 5d 60 61 5b 5d 58 62 5c 5b 53 56 4f 42 44 41 3c 3e 33 23 20 0e 0b 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0b 20 21 2d 37 29 39 39 3e 3c 3e 3d 3e 4a 40 44 39 36 4d 41 41 3f 3c 3e 3d 3b 39 40 3e 42 30 3a 3b 3f 38 43 48 45 38 3f 3f 43 42 4b 55 42 4e 4a 43 41 45 3f 46 3f 4b 43 4d 41 43 4d 45 40 45 42 3d 3a 36 3f 3c 40 3b 36 39 34 31 39 39 32 36 3e 35 35 38 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 49 5d 68 66 69 5f 61 66 6a 5f 69 5b 64 69 60 68 5f 64 5f 5d 69 67 6d 5c 64 65 5c 63 67 61 68 5d 66 62 5f 66 64 66 54 62 5a 60 60 64 5b 59 60 57 59 51 49 3d 41 37 32 2b 29 1b 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 14 1b 1d 29 2d 28 31 39
 3d 38 40 40 47 4e 47 4b 3e 39 3d 3c 36 42 3e 3e 3c 3c 40 42 3a 3f 3f 41 39 43 3b 3c 3b 34 40 3c 42 45 4a 4a 4b 4e 4b 4e 52 4b 4a 43 47 4f 3e 47 47 47 42 4a 41 42 43 3b 3e 3c 31 3c 38 39 3e 43 3d 35 39 2f 34 37 37 36 30 31 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 4a 5d 6d 5f 65 64 60 62 62 5d 62 69 64 6a 60 65 68 62 67 63 5f 62 66 5a 65 67 5d 66 61 62 62 66 6b 64 61 60 59 5d 59 5d 5a 5c 61 58 57 5d 50 54 57 49 39 42 3a 32 29 26 23 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 19 1a 21 23 29 30 32 33 39 35 43 48 48 4b 45 47 3d 37 32 37 3f 3f 36 3d 3d 39 39 3f 30 3f 43 45 44 41 45 3c 3e 40 3f 3f 49 48 43 41 47 49 4d 4d 41 41 44 47 48 49 45 41 3f 3d 46 46 41 40 39 34 40 2f 3e 36 39 39 39 39 37 3a 35 30 32 3b 2c 30 2d 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 3c 4e 68 66 5c 57 5d 61 64 59 55 58 60 64 62 5d 65 65 65 65 69 5e 5e 60 5d 5e 59 62 6a 61 61 63 64 62 62 5a 61 63 62 62 5b 58 57 5b 55 4f 4e 4c 49 3c 35 37 36 2e 30 1e 1b 0d 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 14 20 1e 20 2e 2b 31 36 33 3f 3e 4b 45 52 49 4b 3f 43 36 39 3a 38 39 3b 45 34 39 3a 2d 3f 3b 3c 3d 3d 3e 42 41 47 40 46 42 43 44 4c 44 47 49 41 47 4b 42 46 4c 44 46 3d 3c 42 3e 41 3b 3c 3d 3d 42 44 34 3f 34 3b 3c 35 33 37 39 30 36 33 3c 33 2d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 39 62 62 62 56 52 55 62 5d 5d 5a 60 58 5a 5f 5c 5d 5f 65 62 69 64 5e 62 53 5a 5f 68 62 63 67 63 5f 61 63 6a 66 69 59 58 5c 4f 50 4f 56 44 42 48 3c 38 35 2b 29 26 1b 17 0f 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 0e 1c 1e 1f 2b 2f
 2d 34 34 39 3b 3f 49 4b 49 4a 39 3c 38 41 3e 3a 43 3e 3b 3f 42 37 39 3f 3b 3e 47 41 40 41 3c 39 41 42 45 4a 43 46 43 40 4b 46 45 47 3e 4e 3f 45 4f 43 43 4b 4b 41 3b 44 39 43 3e 3b 3a 3a 40 40 49 3e 40 36 32 35 33 34 37 33 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 43 64 65 66 58 60 60 63 5b 59 5e 5e 60 5c 66 5b 62 5c 58 55 5c 5f 5d 62 5b 5e 6c 62 62 6e 5f 69 64 5d 67 5f 5c 62 5f 58 5c 51 51 4a 4b 42 43 40 32 30 27 28 2d 23 1a 13 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 0e 13 20 27 2d 25 2e 35 34 42 41 3d 42 44 3f 39 39 33 41 3b 35 3e 3c 3f 3d 34 3c 39 3b 39 42 39 3e 41 45 42 3f 3f 46 42 3e 40 41 45 45 4b 42 44 41 42 4a 3d 41 49 42 3f 4a 3c 44 4d 3e 43 45 43 46 3c 47 44 42 45 40 38 3e 36 34 3a 39 35 33 26 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3d 5a 5f 69 64 62 5f 5e 45 5c 5a 5a 63 59 61 5c 59 63 66 5e 6b 61 61 5e 60 68 66 68 66 65 62 5d 5f 63 65 66 56 56 54 59 53 4d 49 47 3c 3c 38 35 2e 2a 2e 24 20 1b 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 0d 13 1e 22 27 30 2e 2c 36 38 3b 3a 46 36 38 40 3b 3a 37 3a 3f 39 3e 40 3a 35 40 3f 3c 33 38 3d 3c 3f 3c 3a 3f 3d 3d 46 40 40 3e 43 46 41 43 44 44 48 3e 44 3f 3e 40 3f 46 45 45 43 48 3e 48 4e 44 47 4c 43 43 41 43 3f 3a 42 3c 36 37 38 2b 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3c 5f 67 66 64 54 56 55 5d 58 59 61 5d 62 5e 57 64 64 5f 63 60 58 5f 64 5b 60 69 65 5a 61 61 65 5d 5f 60 54 5b 5b 55 4e 46 45 43 3e 38 33 2c 2a 25 23 21 1d 1e 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0a 12 23
 21 29 2d 28 2c 33 38 35 3b 3d 41 44 39 41 39 37 47 3c 43 3f 3c 3f 39 36 43 3f 44 40 3d 3b 40 47 4c 48 4d 44 48 42 41 48 41 41 48 42 48 42 3d 43 4b 4c 4d 4c 47 45 40 48 3d 4a 4c 4b 41 4a 4e 4d 47 48 4e 43 40 41 48 49 42 39 2b 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 54 60 6f 62 61 60 65 64 5c 5f 5e 63 5e 62 64 64 60 60 5b 6b 61 5b 5a 5a 66 5c 61 61 64 5f 5b 57 63 56 5a 55 4a 41 49 48 3e 3d 32 2d 35 2b 26 24 1f 19 1e 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 0d 15 1a 20 26 2d 2c 34 38 3d 3b 3d 37 40 3b 3f 3d 41 37 39 3b 3f 39 37 47 3a 42 3e 3b 38 38 44 42 44 4a 41 3f 47 3f 44 46 45 46 41 4d 47 48 47 49 4f 49 50 4f 45 4c 4b 4d 42 46 46 46 4d 46 4e 48 46 4a 49 4b 44 4d 43 53 4b 43 32 31 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 35 54 5f 63 60 64 64 5d 64 63 5e 5f 64 52 5f 64 61 65 59 64 67 63 64 65 5c 65 60 60 62 5d 5b 5c 61 56 47 57 4e 52 45 3b 3e 3d 2d 38 29 2d 2f 22 25 1d 19 09 07 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 07 0d 14 1d 1f 22 2c 2e 2b 29 39 34 3f 3c 3a 39 3d 45 3e 3a 35 3d 42 42 40 38 3a 37 36 3f 3f 3c 43 43 47 47 4a 49 45 42 4c 4c 47 4b 4c 4d 52 4b 48 45 4d 45 44 42 3d 41 44 45 46 41 44 43 43 4b 46 4f 48 43 40 48 49 3f 4a 46 3b 3d 30 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 30 57 68 63 5c 64 62 59 64 62 65 64 64 64 61 64 62 5b 60 60 65 68 65 58 64 57 60 5b 54 61 57 59 4c 50 4e 4a 45 41 42 41 3c 28 2d 2a 20 27 21 23 1a 0f 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 0a 16 18 20 21 2e 2a 33 2e 36 38 3b 38 39 36 3f 3c 3f 3e 3c 40 41 38 3d 3a 39 3f 3e 3a 43 43 49 4c 49 51 56 4b 4f 52 4a 58 47 55 52 4b 4e 47 4d 52 4c 48 43 42 43 3e 44 42 3c 44 44 41 4f 44 45 3d 39 45 44 44 46 49 3f 43 36 24 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 32 4d 5b 6a 64 60 60 62 60 65 5f 5b 63 61 6b 64 64 63 5f 67 61 62 62 5b 5e 5e 60 5b 5b 5c 5a 54 4f 4b 49 47 3e 45 3b 3b 35 31 2f 28 2a 1f 1b 1b 17 06 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0a 18 16 18 26 2c 2d 2e 38 31 34 39 33 43 3b 38 42 37 3d 3b 44 40 3b 37 3d 40 41 3b 45 44 4b 57 58 53 5c 5e 5c 59 5d 57 58 5d 53 56 5a 55 4e 4b 47 48 45 3c 42 3b 3c 43 48 3a 3d 44 48 3c 3f 43 41 3b 38 3e 3e 3a 40 36 32 25 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 27 47 53 65 5e 61 67 61 64 58 61 61 64 66 66 65 59 5d 5f 60 5f 59 5f 5d 57 58 4f 54 50 57 4d 4d 4a 4c 4b 47 38 3b 34 2f 31 26 22 29 25 1b 19 12 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0c 12 1c 22 27 25 2e 2b 2b 34 30 3c 40 35 3a 38 43 3e 40 3a 2f 3c 3d 43 3a 35 42 43 4b 51 59 5f 60 5c 68 63 60 65 65 69 67 6a 66 5b 5a 54 57 4a 44 41 3a 3a 3f 3c 30 38 3f 45 38 46 49 3c 3f 3f 3d 3e 38 3c 36 39 37 2e 2b 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1e 45 5a 5c 5e 51 5c 61 5e 5d 5e 60 5e 59 61 5f 61 5d 5d 5d 60 59 5b 55 54 4e 55 4d 4f 4e 4c 4f 48 46 3b 32 34 33 32 33 31 29 2b 1e 1e 22 12 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 02 06 07 14 1d 1a 20 2a 31 32 32 35 39 36 37 38 3c 43 3b 3a 3b 3a 3d 44 3d 3b 3b 36 46 4a 54 5e 5a 64 66 6a 69 69 74 63 69 6c 6b 64 60 5e 5c 5f 58 56 45 46 41 3b 41 39 35 40 3c 3e 45 41 43 3e 43 3d 36 3c 32 38 3b 35 34 2f 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 22 42 51 57 59 58 55 62 5a 5f 5d 5c 5f 61 60 5d 56 59 59 51 5b 57 54 50 51 4c 4f 4a 4a 4c 41 41 36 33 35 33 35 33 2a 30 23 27 1d 1a 16 17 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0c 16 1f 1b 26 27 2b 2a 2f 2e 33 2e 3f 35 3b 36 3c 3d 3d 3e 37 40 3a 43 43 48 4f 53 57 62 68 5b 6b 6d 66 66 6f 70 70 6a 73 65 66 60 5c 5e 54 44 49 39 3b 3e 39 3b 3e 40 3b 38 47 37 41 3f 43 37 3b 3d 35 2b 32 2c 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 38 43 50 49 4d 55 51 55 53 5a 5a 5c 5a 5b 56 5a 56 4f 4b 4b 4b 53 4b 46 42 43 42 4b 3f 39 35 36 38 31 33 2d 28 2b 25 23 1e 1c 17 12 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0f 17 20 19 25 29 2a 34 2b 2a 35 37 3b 39 41 3d 36 43 3f 40 3a 3e 43 3d 4a 48 55 50 5b 64 5c 60 66 65 68 6d 6d 70 6f 6a 6c 69 62 61 58 55 44 41 3b 37 33 3f 3e 3b 3f 3a 3b 3c 38 3d 3b 3b 36 35 36 33 37 2a 1e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 31 42 42 44 4d 4f 4b 4b 49 4f 4e 4c 51 4c 4d 4d 48 4e 44 46 47 43 41 39 3e 3e 34 3c 38 30 2d 2a 2c 28 26 29 29 22 22 1e 12 0d 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 04 06 0e 12 20 19 23 27 2c 2a 33 2f 2f 34 3b 35 3b 36 3a 3e 44 3d 3b 3b 42 40 46 3e 43 4e 57 52 5b 62 64 6d 64 6a 69 67 70 6c 6d 71 65 69 5f 55 4e 46 43 3b 33 3f 43 4a 3b 3d 3c 3b 3f 3a 3b 34 3c 33 42 39 2f 27 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 28 3b 47 42 3d 44 3f 44 43 4b 4d 51 47 4e 44 44 4a 4b 3a 41 37 42 3a 39 39 33 35 36 33 30 2f 29 27 2e 25 21 29 21 1b 14 0c 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 12 15 1b 25 27 23 33 2c 2f 31 30 32 36 3d 3b 46 3c 40 39 3e 44 3f 45 48 4a 47 46 50 55 5a 56 5e 5f 63 68 6a 68 65 64 6b 69 61 63 62 4f 49 3a 3f 3a 3a 44 42 46 3d 3b 3f 3d 36 39 3b 3a 3f 3b 35 2e 2f 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 2b 34 39 3e 40 38 4b 45 37 41 4c 43 47 49 45 4a 47 3f 3c 3f 38 35 38 2e 33 3b 2a 2a 2a 2f 22 2b 29 26 29 2c 23 1b 0b 0c 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 08 0f 13 22 1c 23 1d 2a 27 30 32 2f 36 39 3b 42 35 3c 3e 3b 3f 44 41 40 3e 41 4b 4f 4a 56 56 51 52 60 5e 60 65 66 61 5b 58 5a 56 58 43 39 40 34 35 35 3f 40 3d 3d 3a 36 35 3a 37 2d 39 34 30 33 2a 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 29 38 3b 39 3b 3f 42 43 3d 39 40 44 44 42 38 3f 3b 38 32 34 33 35 29 26 26 2e 2c 2b 28 2b 21 2e 21 1e 1e 1c 17 0c 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 09 15 1c 22 21 23 32 28 31 32 2e 32 3b 38 33 33 35 41 47 46 42 3e 3e 40 48 4e 45 45 4e 50 54 60 59 5a 4e 59 5f 5d 5d 5e 4c 4e 3e 3f 3e 3e 35 35 39 3c 3f 40 3d 39 37 43 2f 2f 3d 2e 2b 29 26 17 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 30 39 44 3f 3d 37 3d 38 41 41 3e 3b 40 34 2c 2d 39 38 2d 2c 26 30 2a 26 27 2d 2a 2c 2b 2a 2e 28 1a 19 1a 16 08 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0b 0a 12 22 1b 1e 29 26 2e 28 33 33 2f 32 36 41 44 43 41 3f 48 41 45 3f 4a 49 48 52 4d 53 50 52 5c 5b 55 5b 51 4e 4e 48 43 44 3f 3b 41 43 44 41 42 40 35 3e 38 3a 39 37 32 3f 40 2e 34 2f 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 2c 38 45 44 38 47 3b 41 3e 39 38 3a 32 32 33 2c 2b 2a 30 30 25 23 25 2c 28 2a 2b 25 1e 20 1b 11 21 18 10 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 0d 1f 1e 1f 1f 21 29 26 2d 3a 32 38 33 38 3a 40 3c 41 3f 38 2e 46 3e 48 47 43 49 4c 50 4c 52 4b 4d 4b 48 4d 43 45 45 38 3e 38 37 3e 40 3d 33 36 3c 3a 43 37 3b 2f 39 3c 2b 31 31 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 22 49 48 39 3d 3a 3b 44 42 39 33 32 30 2d 28 2d 31 27 27 2e 23 29 2d 25 2c 2a 24 23 1f 18 20 11 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 11 1a 25 26 26 23 21 27 2d 33 33 38 35 39 37 3d 40 42 3c 35 3a 43 45 4e 43 3f 43 41 4b 4b 47 42 47 42 44 46 42 38 3d 41 46 49 3d 3a 3e 3a 39 3b 39 36 30 34 35 2d 2f 26 22 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 2c 39 36 41 36 34 3a 30 2f 37 28 27 2f 25 2f 30 28 28 20 27 1e 2a 25 21 22 26 20 1d 23 15 16 14 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 09 17 15 20 20 23 28 2b 30 2b 27 2d 30 3d 38 36 39 3c 3c 39 40 40 43 3b 45 44 41 47 47 42 41 3e 42 40 41 44 3f 33 3d 3d 44 43 3a 3e 37 3c 39 39 36 36 35 38 36 2b 2c 26 2c 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 26 3c 3a 36 37 34 31 30 2d 25 2d 28 2b 1a 2a 25 26 27 2a 23 2f 24 16 25 1e 27 1a 18 15 0f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 07 0c 0b 17 12 1c 26 21 29 23 28 27 2d 2f 36 37 3b 37 2f 37 38 40 45 41 3c 44 3f 3b 3d 40 44 44 3d 3d 3e 3e 42 3f 3b 38 41 3d 35 44 39 35 3c 34 30 34 29 33 2c 33 2a 36 2f 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 35 3a 2c 2f 31 29 2b 25 24 21 25 26 24 25 25 1d 23 29 24 24 20 20 20 1a 1c 15 13 0a 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 06 0f 13 0d 1b 1a 1b 24 29 1e 22 35 2d 2f 31 38 37 36 32 36 3c 39 38 3e 3e 45 35 3e 36 39 36 32 38 3a 38 39 3c 39 34 3b 3c 40 36 3f 32 30 34 33 36 2f 26 31 24 2a 26 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 14 30 2c 1f 2a 29 1e 2a 24 1b 1c 1f 22 1d 22 2d 16 20 25 24 17 1e 12 0e 11 0a 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0a 0a 0f 15 16 1e 2a 28 2c 1e 24 24 32 31 29 29 34 39 35 34 37 34 2d 36 34 3c 37 33 2e 2e 31 34 35 31 3a 2e 39 36 2f 37 34 39 31 32 2d 34 32 29 2c 27 25 21 24 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 25 28 23 1e 24 24 29 1d 24 16 1c 1e 21 24 1e 1b 1e 1a 18 1a 18 10 0e 08 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 07 08 16 1a 15 21 25 2b 21 23 26 2a 2e 2d 26 2a 25 2d 2e 2f 2d 23 27 31 2d 22 29 26 31 2e 2f 33 33 25 32 2c 30 32 2b 2c 2a 31 2d 24 2c 1e 24 23 20 22 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 16 12 0c 12 10 1e 15 14 19 1e 15 10 14 19 1a 15 1a 0e 14 0f 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 12 0a 12 1c 25 1a 1e 24 1a 1f 20 20 29 21 24 25 1c 1f 15 20 1c 1b 1d 1f 24 29 2b 26 29 1f 25 28 1b 29 2b 2b 27 20 23 28 1f 1f 24 1e 1d 16 19 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 0c 07 09 0e 09 09 0d 0b 0a 06 1a 12 0a 11 0a 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 09 16 16 14 22 1b 28 21 1c 20 21 1c 1a 1b 0f 11 0c 15 16 13 14 1f 26 1f 24 26 1d 25 1e 21 1e 24 2a 25 1e 1d 1a 17 1c 1b 1a 1d 19 10 12 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 03 0e 05 0e 09 0b 05 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 03 11 14 19 19 1c 17 16 14 10 0b 0c 06 06 05 0f 06 11 0a 19 1c 1e 1a 12 12 15 12 0c 19 13 0f 19 13 12 11 12 0a 0e 11 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 03 05 06 05 09 08 06 05 03 00 06 05 03 00 07 06 0a 0c 06 0a 07 00 06 0b 09 10 06 06 0a 00 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
