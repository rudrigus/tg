 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 06 09 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 04 06 05 03 03 06 05 03 03 09 05 08 00 06 05 03 00 06 05 03 06 06 05 06 0b 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 08 06 05 09 03 06 05 03 02 06 06 09 00 06 05 03 01 06 05 03 04 06 0a 04 0d 06 05 03 01 06 05 03 00 06 05 03 06 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 06 06 05 03 03 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 0d 0a 05 03 05 06 05 03 00 06 05 03 01 06 05 03 05 06 05 03 00 06 05 03 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 05 03 06 06 05 03 0b 07 0b 03 07 06 05 03 08 06 05 03 06 06 05 03 05 06 05 03 02 06 05 05 07 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 06 06 08 06 05 0c 00 08 05 03 09 0e 06 04 08 06 06 07 0d 06 0e 10 12 14 08 05 06 0d 09 08 10 06 05 04 01 06 0d 0c 00 0c 05 03 06 06 09 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 00 06 05 03 09 06 05 03 00 06 05 07 07 07 05 0a 06 09 08 06 06 06 13 10 1c 13 07 03 0a 0d 0d 04 0a 06 05 03 0b 0d 0b 0f 09 06 05 03 00 06 05 03 06 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 05 02 06 0a 0a 06 06 0c 0f 0e 06 09 0c 05 0d 0d 12 10 06 09 08 0a 10 10 1b 1f 0d 10 0f 16 18 0d 0b 0a 06 0a 03 11 11 0b 13 03 06 06 05 05 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 03 00 06 05 04 02 06 05 04 03 06 07 07 0f 09 0c 17 0c 08 05 05 0d 0d 11 0d 0f 06 0d 17 11 0c 17 17 25 18 14 15 21 1e 13 11 12 09 08 0a 0a 07 0e 13 10 0b 07 0b 03 06 05 03 06 08 05 03 03 06 05 03 01 06 05 03 05 06 05 03 00 06 05 06 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 0a 06 06 05 06 0b 06 08 0e 0b 06 09 0b 0c 09 0a 0d 16 1a 14 18 11 0f 13 13 10 0a 10 12 20 17 1e 21 24 13 1e 14 13 15 12 14 0f 0c 10 16 06 07 0b 04 00 0d 05 04 0e 06 07 03 04 06 05 03 00 06 05 03 03 06 05 03 01 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0e 04 08 06 05 09 0a 09 05 08 0f 0e 09 0e 05 12 06 10 11 0f 14 15 1a 18 16 22 1d 29 23 2e 25 1c 1c 2b 20 19 13 0b 14 19 1b 0c 11 13 13 0d 10 06 0e 0a 05 06 0d 03 0a 06 0a 03 05 06 06 09 00 08 05 07 00 06 05 03 01 06 06 03 03 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 04 06 0a 03 0c 09 05 0c 04 07 05 0b 0b 0e 0b 0c 10 0e 15 13 12 15 07 09 0b 19 16 23 1d 1e 24 1f 1f 29 21 31 21 20 26 14 16 12 16 14 1f 15 0f 12 1b 08 13 0a 10 15 05 05 08 09 05 06 07 06 0a 03 05 10 05 0e 08 07 06 03 00 06 05 03 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 07 06 05 0e 0f 0b 0c 1b 0c 10 14 12 12 18 18 1d 20 1b 19 1a 1d 1e 21 17 14 22 25 1d 21 19 1f 19 1f 1e 24 18 1f 16 17 19 10 15 0d 13 14 0d 14 03 0a 06 05 07 0b 0b 0b 0d 0e 06 07 10 0c 06 05 03 02 08 05 03 04 06 05 04 00 06 0a 03 00 06 05 03 00 06 06 03 01 06 05 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 08 06 05 07 0b 0e 05 07 10 10 08 0f 04 06 15 0d 0d 14 1e 20 13 13 11 27 25 2a 1c 12 19 24 28 24 23 26 39 22 20 21 27 22 21 23 27 26 26 19 2a 27 1c 15 15 12 19 11 1d 07 13 0d 08 11 0d 06 0a 0b 10 0b 05 16 0e 09 0c 07 00 06 08 05 09 06 05 04 0c 06 05 04 00 06 05 07 07 06 07 03 05 06 05 03 00 06 05 06 00 06 05 06 00 06 05 03 00 06 05 03 05 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 0c 03 0a 06 09 07 00 07 05 12 08 0c 0c 07 0b 0b 06 12 06 16 07 0a 18 13 1c 1e 16 1c 15 20 1b 13 1b 24 23 25 25 2a 26 2f 31 29 1e 21 2a 2a 21 29 25 25 34 2e 2e 29 3b 36 35 30 22 1e 20 1e 10 14 15 12 19 14 17 13 11 0d 1d 12 14 13 13 0a 0b 10 07 0c 06 0b 09 12 04 06 08 0b 06 10 08 04 03 06 05 03 06 06 09 03 00 06 05 03 00 09 05 09 0b 06 05 03 08 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 07 06 05 0f 07 06 09 08 0e 0b 0f 08 18 0a 11 0e 09 1b 15 2b 25 24 25 27 1f 1f 2b 21 2b 31 2b 1f 30 39 34 34 2f 26 31 33 2d 36 3d 35 46 4d 39 40 49 3a 3e 30 2f 2a 2b 1e 18 14 14 16 16 16 17 16 16 15 1d 19 18 15 19 0f 10 10 0c 06 0f 0d 14 0a 06 06 07 06 09 11 0d 06 09 06 05 07 00 06 06 0b 03 06 05 03 02 06 05 08 09 06 05 03 00 06 07 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0e 05 03 03 07 05 05 09 0a 09 08 06 06 08 08 07 0d 17 14 19 15 14 19 16 1a 20 3b 46 33 30 2e 29 25 28 2b 32 34 3e 39 3d 37 34 43 3b 37 3b 4b 61 75 8f 80 86 80 84 5c 4c 38 31 2a 2f 31 2b 30 2a 23 1e 22 17 24 1f 1e 1f 24 1e 1c 1e 1a 24 11 20 12 23 19 0c 14 0c 0d 10 08 07 08 0e 11 0c 0a 0f 06 05 05 07 06 0b 05 00 0a 05 05 03 0a 0b 11 00 06 05 05 03 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 0f 0a 05 09 01 0f 14 0b 0d 0d 0b 0d 10 15 26 14 1b 1a 1b 25 20 18 23 31 42 40 35 3d 39 43 53 56 52 55 53 4b 52 55 5f 58 56 55 58 7a 96 bc ca ca d9 e1 de 9e 83 69 44 49 3d 47 4c 48 50 39 30 33 32 32 35 2f 34 29 34 2e 2a 20 25 2a 21 1f 23 18 15 16 1a 16 14 0c 0e 10 10 12 17 0d 0f 07 09 10 10 0e 05 0a 00 08 05 03 0d 0e 0d 05 0b 09 0e 03 00 07 0c 05 0a 06 05 03 07 06 05 0b 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 01 06 05 03 00 08 09 10 06 07 0e 0a 0b 09 0e 0b 0f 12 12 14 16 19 17 27 20 18 1d 1a 1c 27 25 2a 42 47 4b 51 43 5b 56 5d 66 73 77 65 6d 73 76 6e 72 6e 84 ba d0 d7 e2 f3 ff ff ff f4 91 66 60 66 75 84 5e 54 65 48 3f 37 3c 40 39 33 36 30 3f 47 34 31 2e 31 35 2c 2a 23 20 1c 15 18 0e 10 0b 08 11 0b 15 09 0e 0d 1d 22 13 14 0f 0c 09 0b 05 09 0b 16 0f 0a 06 06 17 09 07 0a 05 03 08 06 05 04 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 03 00 06 06 08 0b 0b 17 09 0c 0b 18 15 0f 0c 14 0a 10 0d 0f 14 13 27 27 24 29 2b 20 23 30 35 33 51 65 64 4e 5a 6c 6a 5c 66 6d 8c 96 88 8f 9e 98 95 97 ab d1 f2 ff ff ff ff ff ff ff ff a0 75 6c 75 8d 9d 81 6b 61 4e 45 3d 4f 6d 61 3c 3c 38 40 3a 3f 41 41 4c 46 3f 30 2b 22 25 21 23 1b 18 1a 13 15 0f 0f 13 11 19 31 4f 37 11 0f 03 08 06 06 0b 0b 0c 10 0d 0f 08 14 0c 06 06 0a 03 00 06 05 03 05 06 05 03 04 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 09 07 05 07 08 06 05 08 06 11 1b 17 15 0f 16 17 11 1e 1a 1d 15 1e 0b 1b 21 2a 30 29 40 35 3c 32 2f 3b 3f 61 63 67 5a 69 7a 90 b4 bd c7 d5 d4 d3 db dc dd cb cd e4 f1 f8 f6 fb f9 fd ff ff ff ff cc ae a5 a6 9f 9d a9 92 7a 66 4c 45 64 95 96 75 59 3e 44 42 53 56 5b 51 5e 5e 50 3f 39 40 35 2b 2c 22 1f 1d 1c 21 16 13 1a 15 3e 65 3a 18 0c 09 0f 0c 06 05 0e 0a 0e 0d 10 06 06 09 13 0c 0a 09 0d 07 05 03 05 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 03 06 05 04 02 06 05 03 06 08 05 0c 0c 14 26 3b 25 12 12 08 10 17 1b 1f 18 15 1a 19 25 34 39 39 59 51 44 48 3e 4a 54 5f 64 66 65 6d 84 c7 ff ff ff ff ff f8 ee e1 cc d1 cf dd e4 fb fa f4 eb d8 da d2 dc e1 cf c6 c8 c2 aa ab bf 9f 88 66 58 53 5d 99 c2 c5 80 4b 51 4f 5c 57 5d 64 6c 6d 64 4e 4a 47 41 39 39 37 2d 23 24 24 21 1b 18 11 1a 28 2a 1f 16 19 03 10 13 12 09 14 06 15 0e 0f 0f 0f 1d 0d 0c 04 0b 08 07 0f 02 09 14 12 0a 06 05 03 00 06 05 04 02 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 02 06 05 08 0a 06 06 0b 08 06 1a 2b 1b 14 11 19 1e 19 1f 1b 21 1d 19 20 2c 46 45 3e 4b 55 4c 4b 51 5d 6d 7a 92 a8 96 6f 84 b9 e6 ff fd f7 ea e8 d9 ca ce d4 dd df ec fc ff f7 f2 ea e3 e6 ed ff ff ee f5 e4 d9 d2 ca d0 bb b7 a1 6a 72 a7 cb a0 80 5e 64 63 66 68 5e 6f 74 6d 64 64 57 63 61 46 41 2e 2c 35 2e 2b 27 19 1c 14 0f 1d 1b 1e 13 12 16 14 13 12 18 19 12 22 1f 06 12 10 19 1c 0e 0b 0b 06 05 07 0a 14 15 10 0b 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 04 06 05 03 02 06 05 06 01 06 07 03 0b 0e 08 0b 0a 06 0b 0c 08 0b 0d 0c 08 0a 18 12 0c 06 12 24 34 2d 2b 29 29 27 2d 31 58 67 5a 52 5b 5f 55 58 60 67 7d 9d db f6 cc 9d ad af c5 d1 d9 da e2 e6 f1 e8 f8 ff ff fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ed e3 dc a3 93 a5 a2 8e 8f 85 84 82 7c 87 7c 83 80 82 82 81 80 78 65 53 59 59 52 4e 45 31 2f 2c 2a 1f 28 26 20 28 27 1c 21 1b 19 17 18 19 1c 14 19 11 15 13 12 13 13 13 11 06 05 0f 15 0d 0e 13 02 07 05 03 09 08 05 03 03 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 05 03 00 06 05 03 01 06 0f 03 0a 0a 05 1b 0b 0e 05 07 11 0c 0f 10 14 0c 18 17 12 1c 2b 44 3e 30 30 39 40 3c 56 73 81 7c 74 5d 79 8a 83 8e 82 8a 91 a3 d3 ec e7 e5 fa e9 ec f6 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 de d9 c4 bf b1 a7 aa 9e 9e 9b 99 94 90 94 92 93 90 81 7a 73 6e 6e 61 59 4d 47 43 40 35 2f 2d 30 32 2f 2b 27 2d 2e 25 1f 2d 1d 1b 25 18 21 18 13 0f 15 11 18 1a 10 13 13 0a 0a 13 07 05 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 04 05 06 05 03 00 06 05 03 00 08 08 08 07 12 0e 0a 06 0a 0b 10 0c 0c 0c 0f 0f 12 13 10 21 26 36 3a 37 3c 3a 42 4f 55 7e 9d a4 a4 91 7d 9c be bb b7 be cb e0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea e0 c3 c2 b2 c0 b7 a6 a2 a5 a4 a3 9c a0 9e 9c 90 84 82 88 8a 72 5f 60 54 54 4c 44 3f 40 42 38 33 34 36 3b 2d 2f 34 25 2a 28 26 25 1c 1c 15 1b 11 12 0c 0c 0a 0a 0a 14 09 0f 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 02 06 05 03 03 06 05 03 00 06 05 0e 0a 06 12 07 0d 08 0e 14 10 0a 13 12 20 19 14 20 1d 1c 23 20 3d 4b 3e 42 3a 44 4e 60 6d 94 cc f0 f1 db c4 b0 cf f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ea e2 d8 d8 cf ca c2 be bc b6 af b0 af a8 a2 a4 a4 ab b3 a2 8e 84 77 70 66 62 59 58 59 51 51 52 55 49 40 38 3d 3e 30 2c 30 31 2d 26 26 1e 22 1f 17 13 17 15 14 07 12 10 0b 13 08 07 0d 05 06 06 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 03 06 05 03 02 06 06 03 03 06 05 09 07 0d 05 08 05 0a 05 0d 11 12 09 1b 14 15 20 1b 1a 24 2e 29 24 2d 2c 3d 4f 4b 47 3d 4b 59 6e 94 c7 fb ff ff ff ff ec e2 ec ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f9 e8 dd e1 e6 e2 da d4 da d1 d8 dd d7 d6 d8 d6 cb c6 c3 bf c2 a9 af a3 9e 99 92 8b 8a 80 7a 77 76 7a 6d 67 5c 54 4b 41 46 41 4a 39 37 2f 31 27 28 28 20 1a 18 16 22 15 0f 0e 0a 0f 04 10 0e 0b 06 07 05 04 09 06 05 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 06 05
 03 00 06 05 03 00 06 05 03 02 06 05 06 0c 06 09 03 11 06 0b 17 0b 16 12 17 1b 19 19 23 23 29 34 33 35 35 40 3f 4b 59 5f 69 7f 91 a5 ca e8 f6 f9 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec df cf d4 d0 d8 d6 cc cc cd d0 df e4 ef ed f5 fd f7 f9 f1 e7 e2 d4 cb bd ae ab a6 a0 a0 8d 95 92 8b 8d 82 7e 84 82 7e 6f 5d 67 5e 52 4d 51 44 44 3a 2e 32 29 2e 24 27 1d 1a 11 0d 0f 0d 0b 11 0d 09 07 05 03 09 06 09 04 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 08 05 03 06 0c 05 0d 00 06 06 17 16 18 0e 18 19 22 21 25 29 22 34 30 39 41 48 4c 4b 54 5d 65 6f 81 82 92 9e b3 b8 bf ca d1 e5 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e0 d8 d4 d9 d5 da de d1 c9 cb c8 d0 df e6 f8 fc ff ff ff ff fd f7 f0 e1 dc ca b7 bf c0 b6 b0 a5 a3 9f 9c 95 8c 8d 96 84 8a 83 7e 79 67 69 65 63 62 56 52 46 3f 46 36 2d 30 20 25 2a 1f 1e 15 15 18 0f 06 05 03 0b 06 0d 05 00 06 06 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0a 14 05 06 0c 0a 05 0a 17 12 1b 15 15 14 18 27 27 2e 33 36 3c 43 48 47 54 59 68 73 71 7f 89 8c 95 94 9e af b4 c0 c2 d0 d5 e4 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e3 d9 d8 e3 dc e3 dc dd d7 dc d2 ce d0 d0 d7 e6 ed ef f6 ff ff ff f8 f5 df de db d8 d6 cf c7 bb b5 b6 b1 a4 9c 90 93 98 97 8e 8d 8c 89 87 80 84 7a 78 72 70 5e 51 4d 45 35 35 3f 3c 26 26 29 18 1c 18 0f 09 08 0b 0b 0d 06 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 07 02 06 07 05 05 06 05 06 0d 06 11 14 10 20 18 17 20 2b 2a 31 37 47 52 55 4c 5c 5b 6d 75 82 84 99 9d 9f 9b a3 b3 ab be be c6 d3 db dd ec fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f7 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 e8 e1 d5 e2 e0 df e2 e0 db dc d2 cc cc ce ca d0 d3 d0 d5 e5 f0 ee f6 f3 ef f1 f1 f0 ea e1 e5 d5 c7 c9 c8 be b8 b0 9f a3 9b 98 9a a5 a5 9f a3 93 87 89 7c 7b 75 70 63 63 54 50 4b 46 33 34 37 2d 2d 21 1a 0b 10 18 06 07 06 07 0a 09 06 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 04 06 05 04 07 0b 0a 07 10 0a 1a 1f 1f 1c 21 2e 34 36 46 46 54 5f 61 6b 6f 77 86 8c 97 a4 a1 a9 ae b5 c2 cb c9 c9 cc de d8 df f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc fa fd ff ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f5 f2 e6 e9 e9 e5 e9 e4 e0 d8 da d0 d1 d3 d6 cf ca d4 cd d1 d7 dd e3 e4 ed ee f2 ef f2 fa ff f6 f5 f0 e3 de db d4 d3 c4 b8 b6 af 9f a1 ab ae a7 ad a1 9b 90 85 7f 7c 79 78 72 67 64 5e 5a 51 4f 46 43 35 2b 23 13 0f 0d 06 18 0f 10 06 07 05 0e 07 07 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 08 03 06 06 05 03 08 06 07 12 0f 06 06 0c 06 10 16 0f 18 1b 24 35 33 41 44 40 4a 5c 68 6a 6e 85 89 95 96 a2 a7 af aa b2 b7 bd c4 d3 df e1 e5 e0 e4 e9 ed f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f5 fb f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fa fb f5 ee f1 f3 e8 e8 e9 e7 e3 e4 e0 d5 d9 ce ce d3 db e4 de e1 e4 e4 ec ed f3 f0 eb e1 dd ea e0 de dc dd dc db cc d2 cb cb c5 c4 bd b3 b2 a8 ac ab a2 9b 9b 97 90 8b 88 8d 8a 89 7c 6f 62 5b 64 5b 5d 4b 33 2f 2b 1d 24 19 1f 0f 14 14 0e 08 09 09 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 05 07 05
 0f 04 08 0a 0b 0d 1a 1d 20 27 2c 38 40 59 5e 70 6c 70 85 92 9b aa b3 b0 be b2 b3 b7 be b6 c8 cf d5 d5 e1 eb f0 f7 f3 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff f4 eb f1 e8 e7 ef df e0 e3 e3 df da dc de e6 f1 ec f4 f5 f7 fc fb f2 ea df d2 cf c5 c9 c3 c1 bf b9 b6 b5 b6 b7 bd bb bc b9 bd bd b4 b7 b5 a9 ae a0 a2 9b 9f 96 9d a3 aa a0 99 8b 7e 78 6a 62 5c 4f 44 3e 27 2e 25 28 1a 19 17 1a 0c 10 06 07 04 04 06 05 03 00 06 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 08 0d 0c 0b 0d 0e 15 0d 18 1e 23 2a 3a 42 46 58 5c 5f 72 7d 93 a2 b2 bc c4 c6 cd ca d3 d0 d8 d8 db e0 dd e0 e6 f0 f2 fb fe ff ff ff ff ff ff fd e3 eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f3 ef ee ef e7 ed e5 da dc d6 e6 e7 e9 ff ff ff ff ff ff ff fc eb e1 e0 d0 d2 c5 c3 bc bb b8 b0 b9 af b2 b0 b4 bb a5 a8 ab a0 a9 b2 af ad af ab ae a8 a5 a3 b0 b4 bf ca c2 b2 ac 85 77 66 59 56 4b 45 33 2b 29 30 2a 1a 20 19 19 0c 0e 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 02 06 05 03 05 06 0c 08 03 06 05 03 01 0d 15 10 15 19 1a 2a 3a 43 4c 50 5a 61 73 7a 7e 7b 90 9a ac bf cb dc e2 e8 ef ed f0 f0 f1 e8 e7 f2 f5 ff ff ff ff ff ff ff ff ff fd f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fc fb f4 f4 ed ef e1 e9 e6 f2 f8 fb ff ff ff ff ff ff ff ff ee e9 e4 dc dd e1 d0 c9 cd c6 cb cd cb c5 c2 c3 b9 bb aa a3 a6 aa a5 97 9d a0 a8 a1 98 9e 9e af aa bc d6 e8 e6 e0 c7 a5 86 6b 4d 48 46 49 48 44 44 3c 32 30 29 1f 16 0a 08 00 06 05 09 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 0a 06 03 05 06 05 0a 00 06 12 06 0a 0a 0b
 1e 21 27 2b 45 4e 53 58 5d 63 71 86 93 92 90 91 95 9e b6 cb c6 de e6 e8 f2 f0 f3 fb fb ff ff ff ff ff ff ff ff ff fe f3 f1 eb f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fe f7 fd f8 f3 f7 fb f7 f9 ff ff ff ff ff ff ff ff ff ff f6 f5 f0 f3 ed e7 e9 e5 dc e1 e1 e2 da e1 dd de d9 c0 c4 b8 b1 b1 b1 a8 a0 99 91 96 92 94 91 a4 a3 ac c4 de e8 eb e4 c0 98 7b 65 53 55 49 4b 54 5a 4f 3c 3c 31 2d 18 0d 13 0e 0c 0c 07 02 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 0f 0c 0a 0f 1b 17 1c 24 36 41 53 5c 4e 55 5e 66 6b 81 8f a8 a8 99 9e aa ac af c5 cf cd d9 dd de e6 f1 ff ff ff ff ff ff ff ff ff f9 f6 ed e9 f8 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fa fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ff ff fa f5 f4 f4 f3 f8 fa fa ed f1 e7 d8 ce c5 ba be b4 a9 a7 9b 98 95 8e 8d 8a 87 93 98 a0 b6 c5 d0 c9 bb a0 89 6e 63 61 5b 50 44 4c 58 50 3e 37 38 20 1f 1c 16 0a 0f 05 04 06 05 06 01 06 05 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 07 09 0e 13 11 15 26 1f 22 29 25 43 5d 63 60 5c 65 66 72 83 7b 90 a8 cc db ce ba bc be c6 c9 d5 df e0 de df e5 f5 ff ff ff ff ff ff ff ff fc f4 f8 f9 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 f8 ea dd d0 c9 ca c9 c5 b8 a3 9c 91 95 8a 8b 8e 87 8d 95 9e a2 aa a7 a3 90 86 76 6e 65 67 55 59 4f 53 49 55 3f 3c 33 31 2f 25 1c 18 12 0e 06 0a 0b 03 06 07 05 09 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 02 06 08 09 0b 0a 08 14 1c 2a 46 49 3f 4e 5d
 6f 7b 82 80 83 83 85 82 8f 9c ac d1 ea f8 d5 ce ce cc d6 dc e7 eb e4 ed f8 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ef e5 dc e1 db d3 d2 c3 b1 aa a1 9b 94 8d 90 92 92 8b 91 91 91 8e 8a 80 79 74 6b 6f 6a 6e 66 63 57 55 49 4e 48 47 33 3a 30 2e 1e 16 0f 11 06 0b 02 08 05 0a 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 05 00 06 05 03 0a 06 05 0f 0d 12 10 1b 25 4e 88 87 86 86 95 b3 c6 c8 ca d1 c2 c9 bc b8 bb cc d5 e9 e9 e2 cb cc ce cd d9 e3 f1 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 f4 e9 eb e0 e8 d0 cb bb a9 a6 94 8e 90 91 93 8f 98 89 8a 85 7e 7f 7c 76 77 6e 6e 6b 74 71 77 6f 69 64 52 4b 49 4d 40 30 33 32 23 12 15 0f 05 0c 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 07 09 11 14 18 1e 24 2d 3c 71 bf d1 c4 d1 d3 f0 ff ff ff ff ff ff fd f2 f5 e6 e5 e9 e4 e3 d5 cf d0 e4 e5 ee f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff f9 f4 ee eb d5 cc c0 b8 b2 a7 9e 98 9c 92 8e 89 8b 84 85 7b 75 7a 79 76 7f 7a 81 84 8b 89 7e 7c 7f 6e 63 5e 53 4c 49 3b 51 43 30 24 1c 17 07 0f 0d 09 05 06 05 04 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 08 08 13 0f 13 0f 1d 30 36 40 5a 82 ca ed f3 ff ff
 ff ff ff ff ff ff ff fb f2 e7 d7 e0 e1 dd e4 d1 d6 e3 f2 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e9 df c0 be be b1 b0 ac a1 9d 9a 8f 8a 8a 86 7f 88 80 89 86 84 8d a0 96 99 96 91 8f 8f 76 7c 6c 66 65 5e 5f 54 50 45 3c 33 25 1b 16 0d 13 07 06 06 03 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 0c 09 05 04 06 0f 11 19 2e 4c 4d 5b 72 93 ca ed ff ff ff ff ff ff ff f3 e6 e0 e0 de de d5 d5 d0 d0 d0 d8 e8 ea fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ed e5 ca c6 b6 b3 b9 b1 aa a0 98 95 89 83 8d 86 8c 8d 96 a2 a8 a3 a2 ad a3 97 99 8e 8b 88 73 6b 6b 70 6e 75 69 5f 5d 54 41 34 24 15 14 0f 0d 0d 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 06 02 0a 06 03 02 07 05 09 14 19 1f 3e 57 69 75 72 91 ae dd ff ff ff ff ff ff ff f0 e0 cf d6 d2 d6 dc d9 d0 d3 d4 d9 df ec ef fe fc fe fd fb f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f3 e7 df cb c7 c5 c0 b3 b3 a8 9a 98 93 8a 90 95 99 a1 aa b7 bc b3 b1 a9 a4 ac 9f 9b 86 84 7a 6d 75 77 81 82 7c 70 6e 5e 5c 51 41 2d 26 17 16 0a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 03 06 05 03 0e 06 16 10 1b 2a 3b 55 70 80 91 95 ad b9 f4 ff ff ff ff
 ff fe f3 dc d5 cf d3 c8 d8 e4 d7 d0 d2 d0 db e5 ef f8 f1 f4 ec f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 eb e0 d6 ca ce c6 bf ba a6 a2 a6 9e 99 9e a6 a6 c1 c2 ca c1 bd ba b6 b7 b9 b1 a0 96 8b 7d 78 77 77 85 88 8b 83 7f 77 6e 61 50 39 30 2b 1c 17 05 05 07 06 05 03 06 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 04 0e 16 1a 2d 36 46 5f 64 79 84 97 9c af bd d7 e9 fb ff f4 f4 e3 d6 cf ca ce d1 d6 df d2 cd d1 d2 d9 df e2 e3 e4 f1 ef fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f0 e0 dd d1 ca cb ca bb b3 ac ab a9 a0 a5 b1 c4 cc cf d7 cc c6 c0 c4 cb ca c1 b8 a2 9e 8d 8b 82 83 7d 86 89 93 92 86 7c 6f 5f 4f 3f 2f 1e 14 14 0d 0a 07 06 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 01 0a 05 09 1b 23 37 43 52 5e 62 74 7e 96 a6 ad b0 b5 cb d0 d9 df d6 d5 c9 ce c0 c1 d1 d5 d4 d0 e1 ce d1 d8 d2 d7 e5 ec ee fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ec e4 d7 df ce c9 c8 c2 be b1 ba b6 a5 b4 bb d4 db d3 d8 dc d2 cf d8 d9 dd d7 c8 ba ad 9d 88 87 7c 7d 89 8f 96 9c 97 84 84 66 58 4a 38 35 27 1d 0f 05 06 06 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 09 0f 12 2f 47 52 50 67 6c 73 80 8c a2 ac a9 b4 ba bd bf c3 bc bd
 c6 bb be c2 c1 cf d3 ce d4 cd d2 d8 da e7 ec f0 ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fa ef e0 e3 d5 d4 d0 d2 c6 bc b5 bc bc c7 d4 d5 df df ee f2 ee fb ec f2 ea e9 d8 d0 bb a1 99 91 8a 7f 87 83 97 a3 98 92 87 7b 65 5b 51 3f 31 29 20 0f 09 05 05 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 05 06 07 0a 06 0a 13 27 44 52 55 5f 61 6b 6c 78 85 94 ab b3 b5 b7 bf c0 c1 bd c3 c1 bc ba c0 cb c6 c8 d0 d4 db d8 de e1 eb f0 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f8 f0 ec d8 db d6 d0 cc c4 c0 c1 bd c3 cb da e2 eb f1 fa ff ff ff fc ff f3 f2 e0 d5 c0 aa 99 96 87 82 89 84 8c 93 a0 a0 93 88 74 6f 5b 52 41 3e 30 17 0f 05 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 08 09 05 0b 12 21 37 4d 53 5f 68 69 72 72 78 84 94 9f b3 bd c2 be b8 c0 c1 bf c6 c0 c1 c4 c4 c4 ca ce d0 d5 d6 e5 e9 f2 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ed ee ea db d8 d9 d2 d2 cc c0 c1 c3 d1 da e8 ee f2 ff ff ff ff ff ff ff ff f9 de c6 c3 aa a9 9c 99 86 81 79 7a 88 9b 9e 9f 8f 81 7d 63 5c 58 48 3b 27 1e 08 0d 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 07 01 0b 0d 15 14 1e 2e 49 50 66 6d 7a 81 80 7c 88 8a 95 9f a9 bf c8 be be be c3 bb
 c3 cb ca c9 ce d0 cb d2 da e0 e2 ec f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f8 ed e8 df d4 d4 cf ce cc c5 c9 d3 d5 e8 f0 fd fc ff ff ff ff ff ff ff ff f2 d0 c7 b9 b1 a5 a3 92 84 86 78 7a 7a 8a 95 a7 a4 a4 95 89 78 65 56 46 32 19 10 06 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 06 0b 09 0d 15 1f 2e 3d 4c 60 6d 77 76 83 8c 9d 98 a0 a0 af bc c1 c6 c5 c1 bc c0 c3 c5 d0 cc cf d4 d4 d6 d7 da e4 e5 e5 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f6 f0 e3 e2 da d5 d3 d4 d2 d0 d4 d3 dd f1 f7 ff ff ff ff ff ff ff ff ff ff eb d2 cb b9 ac a8 9c 96 8b 86 7a 7c 79 82 8c 9f ad ad a5 97 82 73 69 5c 4c 37 1c 09 0b 06 05 04 02 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 05 0a 08 19 24 3d 4a 4f 62 70 72 78 8c 8f 91 a9 a5 a7 af b3 c3 c0 c2 bf b1 bf c2 d2 ca d8 d7 dd d7 d9 d4 e1 e2 e6 f1 f5 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f1 ee e4 e5 de d5 da d0 d9 d3 d4 d8 e3 ee f6 ff ff ff ff ff ff ff ff ff ff f6 e7 cf bc af aa a0 9d 95 8d 85 7f 74 76 7e 81 8f 9d a0 b8 a3 9f 8b 7c 6c 5d 4d 2e 1c 0c 06 09 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 07 06 16 27 43 4d 46 56 60 72 75 7b 7c 8a 88 96 9f a9 b2 b5 c0 ba bc b5 b9 be c6
 d4 d7 d3 de e5 ea e1 e2 e1 e9 ea ef fd fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 f1 e2 e2 d9 dc da dd e2 e2 e0 dd ee f2 fd ff ff ff ff ff ff ff ff ff ff fa de c9 c0 b5 ae a3 92 93 90 7f 7d 81 73 7a 82 85 8d 9e ae c0 b5 a6 8d 7e 6d 61 50 25 16 0f 09 03 05 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0d 08 0f 25 3a 56 55 49 48 56 68 75 79 80 85 91 9b a1 b0 b0 b7 b9 bb bb c1 c7 c6 cf d3 de d5 dc e6 ee ee e6 e1 e7 ee f0 f5 ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f3 ed eb e5 d9 df e3 dd e5 e6 e2 e8 e0 f2 fc ff ff ff ff ff ff ff ff ff ff ff e7 da c2 c1 b2 ad aa 97 92 84 84 88 7f 82 80 81 83 84 8b a0 b5 c7 b6 a9 99 7f 71 57 43 29 0c 05 03 00 06 05 03 00 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 07 06 0b 10 1c 37 4b 59 56 49 48 4f 5c 6a 7d 86 8a 9a a4 ac ab b2 b5 b8 b9 c6 cd c6 c4 d5 de df e2 e0 e5 f0 e6 ed e7 de eb eb ef f9 fa fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f7 f1 f0 e7 e4 e1 e0 dc e1 da eb e3 e9 e7 f3 ff ff ff ff ff ff ff ff ff ff ff f4 de d8 c1 be b4 ae 98 9a 8d 8f 86 8a 88 83 7d 80 85 80 81 8c 95 af c8 c5 af 9e 82 60 44 31 1d 0a 07 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0c 06 05 03 05 0a 08 07 1e 27 49 68 60 63 54 42 4d 48 63 7e 83 a0 9e 97 a9 af b5 b8 bb c4 c6 cc d2 d6 de
 e4 e7 e8 e4 f5 ea eb e9 e3 eb ed ed f8 fc fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f6 fb f7 ec ea e9 e5 e1 df e7 f4 e6 f0 f8 ff ff ff ff ff ff ff ff ff ff ff fe f2 dc d0 bc bc b6 a7 9a 8e 8e 8b 8f 92 87 84 90 84 8a 84 85 86 88 a9 cd d5 cb ad 90 66 49 35 20 0a 05 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 05 06 08 0a 04 0a 0c 14 1f 3c 56 65 65 59 53 4b 5a 4e 65 6b 86 a0 9f a7 ac b2 ae b4 ba c4 cf d0 da d3 e9 eb ea e9 ea ef e8 ed e2 ec e8 ed e8 f9 f8 fb ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f4 f8 f1 f1 f2 e0 e0 e6 de e6 e6 f6 f2 fb ff ff ff ff ff ff ff ff ff ff ff f8 ea de d6 ce c5 b3 ad 9a 94 94 94 8d 93 91 8c 88 8c 89 90 85 8b 8c 8a b2 df d3 be 9f 74 54 38 25 0c 07 02 06 05 03 00 06 05 06 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 04 0c 06 09 15 2d 48 5a 69 70 63 5a 50 5b 55 59 6a 6f 91 a4 b3 bd b1 b7 b5 b8 c4 c8 dc da df e7 e9 e7 f0 f5 f2 eb ee ee ec e5 ee f3 f1 f2 f3 ff fb f6 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f3 fd f3 ed e8 e8 ea e4 e4 e5 e4 eb f3 f3 ff ff ff ff ff ff ff ff ff ff ff ff fd f2 df d8 cb b7 b2 a7 a0 9c a0 93 92 97 93 92 8b 95 8f 8e 88 8e 88 8f 9f c8 dd cb a6 82 59 46 20 18 03 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 0f 0c 0a 0e 10 2d 53 65 76 69 6f 5f 52 59 5f 5d 63 70 8b a6 b8 bd bb c4 be bd bb b9 d7 dc e9 f0
 f5 f3 f5 f5 f7 f4 f5 ec f2 f3 ec fd f6 ee f8 fa f6 f7 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 f8 f5 ec e4 e7 e0 e9 e2 e0 e2 ee fb fb ff ff ff ff ff ff ff ff ff ff ff ff fd ee d9 dd c9 c2 b2 a7 a2 a8 9e 99 9e 97 8c 91 96 8f 94 86 92 8a 95 98 9b c6 e5 d0 b1 88 60 48 27 1a 06 00 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 03 06 06 05 05 06 0c 16 19 38 58 67 73 70 6e 68 56 58 5e 64 65 72 80 9a c0 ce d4 d7 cb c7 cf d8 dd e0 ee e4 f2 f7 f1 ef fc f1 f4 f9 fd ee f8 f4 f5 ee f2 ee f0 f5 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f5 fd f3 f4 f3 e5 e9 e0 e4 e1 e8 f2 ed fc ff ff ff ff ff ff ff ff ff ff ff ff ee ed ec d1 cb bc af ab a6 ab a6 a4 a1 a9 94 98 99 93 8f 9c 93 9e 91 94 a4 b0 e1 e7 bf 97 70 59 3d 24 08 00 06 05 08 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0b 09 0f 0d 20 30 5a 6a 75 74 72 64 5d 51 5a 5d 6d 77 7b 8c b5 d0 de e0 d5 d0 d1 da dd ec f0 ee f5 f0 f4 f5 ff ff fc fe f7 ed ec ef f0 f1 ee f0 ea f9 f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f9 f5 f6 ef e8 e7 e4 e8 e6 eb e5 f2 fc ff ff ff ff ff ff ff ff ff ff ff fb e7 e5 d9 d6 c6 b7 ac a7 a2 aa a3 aa a0 9e 9a 9b a2 a1 9b 98 9a 9f 96 99 a7 a4 d4 e4 d2 9e 6c 59 3a 23 0d 07 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 06 05 06 10 1c 1a 2d 4a 63 71 68 70 70 62 5b 61 5b 64 70 77 86 97 ae c9 d2 e1 dd da dd e3 e5 e9 f3 ed
 f7 ef f5 ff ff ff fc f9 e9 ef ee ee f2 ef f4 eb f9 f6 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f8 fc f5 ee e9 ee e9 e6 e9 e7 e3 ee f8 fc ff ff ff ff ff ff ff ff ff ff f8 e6 dc db cc b9 b9 b5 ad ab ad a4 ab a7 aa a9 a7 a1 a0 9e 95 96 9c a0 9f 9a a7 bf eb d5 ad 85 60 45 2e 13 03 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 08 08 06 09 0a 10 1c 2e 3e 52 65 73 72 6b 64 62 5a 62 64 6c 6d 7e 8a 9a b6 d1 d7 e0 dd db db db e1 ec f4 f6 f2 f1 f6 ff ff ff fd fb f3 eb e6 e6 ea ee f6 ed f7 f8 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fa fb f9 fe ed f0 f1 e6 e2 e7 e3 ea e7 e8 f1 ff ff ff ff ff ff ff ff ff ff fa eb e1 d7 cd ba bc b6 b5 ad b0 aa aa ad a9 a7 ab aa a5 9f a0 97 a2 9d a5 96 a5 ba d2 e0 b5 92 77 51 3b 22 0a 06 05 03 04 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 0b 08 07 17 19 26 3f 4e 63 6c 6e 62 62 5e 56 5d 61 6a 68 72 81 89 a8 c7 d4 d5 e4 dc e0 e4 e3 e5 e5 e9 ea fb f0 ff ff ff ff ff f6 f3 f9 f5 eb ec e7 eb f7 f5 fb fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fd f7 f4 f0 ed ed ec e8 eb e2 ec e5 eb f5 ff ff ff ff ff ff ff ff ff ff ff ed d9 cb c6 be ba b3 b5 af b0 b0 a6 ab af ae a9 99 9d a0 9d 98 9b 94 99 91 a3 9f c3 df c8 a7 85 56 3c 23 14 06 05 03 00 06 05 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 06 05 03 05 08 0d 12 21 38 4e 63 75 7c 74 63 5e 63 64 67 63 6a 70 73 7c 89 a3 cc ed ff f6 f1 e5 e7 de dc ec f0 ee
 f5 f9 ff ff ff ff f6 ff ff ff f0 ed e6 ec ee f0 f0 f5 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f5 f2 f1 f2 ea ec e6 e8 e1 e6 e4 e5 ea f4 f5 ff ff ff ff ff ff ff ff f8 f4 db cf c3 c3 bd b9 ac ae ae af b3 b0 b1 ae ac a9 a7 9d 9f 99 96 8f 99 95 9a 9d 9a a4 d6 c9 ae 89 62 44 27 10 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 02 06 19 22 33 49 56 66 76 7d 72 6d 62 63 67 72 6e 6c 70 79 8b 9c b5 c0 e3 ff ff ff f4 eb e1 e2 e8 ef f0 f7 fd ff ff ff fa fc ff ff ff f5 ea ec e6 e9 f3 f5 fb fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff fd f6 f1 f4 ec ef ef e2 ec e2 e1 e5 e8 e6 ee e4 f1 f1 ff fb ff fa fb f5 eb e2 db c5 be bc ae b8 b3 b5 ae a3 b1 af b4 af a9 a6 9f 99 9e 90 8d 95 94 90 9b 9f 99 9f c2 cd b0 9a 6a 44 2a 12 0a 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 1b 28 4a 62 6b 78 7a 7a 6a 6e 72 68 6a 73 79 76 76 7c 88 a5 c1 c8 da f8 ff ff f2 eb e3 db e2 f1 f7 ff ff ff ff ff f9 ff ff ff ff e9 e9 ee ef f4 f5 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 ff fe f6 f6 f6 ef ec ef e7 ea e8 e5 e6 e4 ed e4 ee e7 e3 e2 e5 e5 ec e2 e1 de d3 d9 c7 c0 c1 ba b6 b8 a9 b8 b9 b0 b0 a8 a9 a6 a5 a4 9a 9d 8d 9b 90 8f 95 97 92 91 97 98 ba c6 be a2 7d 5a 28 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 0c 10 20 3d 4d 69 70 7c 87 7f 71 71 70 74 78 75 72 80 85 84 a1 be bc d3 d3 ea ec eb ef e0 e4 e8 e8 ef fc
 fe ff ff ff fe ff ff ff fb ef ee ef ef f5 f6 f7 f9 f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb fb fd ee f5 f1 e9 ed e9 e3 e8 e5 e6 e4 e4 e8 df e2 e5 e4 e0 e1 e3 e3 db d6 d1 cd cb cc bc c2 bb b3 b0 b7 b1 ae a7 aa a1 9e a2 a0 92 95 99 92 8f 92 92 96 91 8c 8b 8a 95 a4 c0 bc ad 7c 56 31 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 05 05 0a 15 2d 4a 60 76 84 7f 87 82 77 72 79 77 75 80 81 82 8c 99 b4 d1 d4 db df ea de e7 e6 e9 e6 ea eb f8 f9 ff ff ff ff ff ff ff ff ff fe fb f6 f7 f5 f6 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff fc fa f3 f2 e7 e7 f1 ee e5 eb e7 e5 e1 e0 e7 e0 e4 e4 e3 df e5 d8 e1 e0 e4 df d1 cf bd ba b1 b8 b4 b6 b7 b2 ad a9 a6 a4 9e a3 9e 95 93 98 97 95 92 97 94 91 92 96 87 91 9e ba c0 b4 8e 5a 2a 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 01 06 05 04 12 18 43 51 66 86 8f 8f 94 90 75 79 78 74 7c 7f 83 83 89 9b b7 e5 df df e7 e5 e7 ec ed e9 f4 eb f0 f3 f9 ff ff ff ff ff ff ff ff ff ff fa f6 f5 ff fd ff fd f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f9 f6 f1 f0 f4 e6 ec e4 e3 e6 e3 e0 e4 e4 e6 e0 e3 eb dc da de de e5 e8 f6 f4 e1 d5 cb bd ba b3 b4 b2 b0 ad b1 b0 a1 a6 a6 a3 a4 a0 90 97 9d 9b 97 9e 9c 98 8d 84 8a 87 92 a6 c1 af 89 5d 26 0a 06 05 03 05 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 0f 11 25 38 5e 70 7e 90 9a a0 94 83 77 75 78 78 87 89 92 91 9c c1 f2 f5 ec e6 eb f6 f7 ef f1 f7 f6 f8 f9 fa
 ff f8 ff ff ff ff ff ff ff ff ff fd ff f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f4 f6 f0 e7 eb ea e3 f0 e6 dd e4 e2 e3 de e1 e6 df e0 de da db d5 d7 e6 f0 ff ff f1 e7 d8 be be b3 b3 b6 ab b2 a5 a8 aa a6 a5 9b a7 a0 98 94 a0 9a 98 94 97 97 94 8f 90 8a 92 a1 ac ab 8e 59 28 0a 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 0b 16 2a 43 66 7c 8b a3 aa ab a2 91 84 80 84 83 8e 92 8f 9d aa c9 f6 ff fb e9 e6 f0 fd f4 fb ff fa ff ff fe ff fb ff ff ff ff ff ff ff f7 fe fe fa fd fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb f2 fe fd f1 fa ec ef e4 ea ed e2 e4 e3 db df e0 df de e2 d4 db e1 d6 db da d0 db db ec f1 f0 eb d3 c2 be b6 ae b3 ad a8 ad a3 a8 a0 9e ad a1 9d 98 9c 9f 92 96 93 93 99 9b 95 9b 90 96 9c a6 a7 8a 53 26 0e 06 05 03 04 06 05 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 0d 15 2b 4d 63 7e 98 a5 b3 b1 ae 9d 93 8d 8d 8a 96 9a 9e a9 c4 df ff ff ff fa e1 e5 ea f0 f7 fd ff ff ff fd ff fb fa f8 fe fd fb fe ff ff fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fb f6 fa ef ee e9 ea e6 e7 e3 e2 e2 e0 e3 df da e0 d9 e0 e4 de e8 da d3 d5 db cf db d5 d9 d8 df d2 ce be b9 b2 b4 aa a9 a9 9b 9f a3 9e a9 ad 9f 9b 99 93 8c 8a 8c 8b 94 93 99 95 9b a1 98 9d a1 85 4e 20 0f 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 04 00 06 05 0e 1b 29 4d 67 7b 9d aa b8 b5 b1 ab 9c 93 92 96 97 9f ac bc dc f6 ff ff ff ff eb e8 ed ee f5 f5 f4 f2 fd f0
 fb f6 f1 f6 fa fb ff fd fc ff fe fa fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 f4 ff f3 f5 e8 e5 e5 e4 e2 e5 dc df df dd e2 df da dd dc d6 dd d5 d4 d4 d3 d9 c5 cb c9 d0 cf cd d1 cb bf ba b7 b5 ad ab a1 a4 a0 a1 a3 a6 a2 9b 99 9a 90 91 8a 85 86 84 86 90 88 94 8e 89 8b 91 98 7b 4f 1c 0b 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 0b 06 05 0d 1f 36 59 6b 7a 95 b3 bb c1 be ab 9e 9c 9b 9f 9e ab ae c6 e0 ff ff ff ff f9 e9 e4 ef e8 ea ed ef f3 ff f8 f5 f0 f5 f3 fa fa f7 fc ff fa fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe f7 f1 ec e6 ef e1 e0 de df d9 d9 d5 de db da e1 dd e4 d8 e0 dd d7 d8 d3 d3 d4 d4 d2 d5 c2 c8 c7 c6 c9 bf bf bc b3 ab ad b1 a4 9d a3 9c 9e a0 9f 95 9d 95 9c 8d 89 7e 86 7f 8a 88 84 87 8b 7d 80 8c 89 7b 4b 1d 09 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 05 0f 22 3f 59 68 84 9d ab ba bd b4 b2 a2 a2 a2 9c a1 a7 b1 d5 f8 ff ff ff ff f7 ee e4 e6 e6 ea e9 ea f5 f5 ee ee f0 f8 f6 fa fa ff ff fe fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff f6 f4 f7 ec e3 eb ec df da e0 d8 d8 d0 d0 d0 d6 d9 d5 d9 db da d5 d5 d9 dc d9 cc d9 cf ce cd ce cd c7 d1 c5 c1 bc b8 ac ae a5 9f a1 a3 9a 9b 9a a4 9e 9b 98 95 90 8c 8b 85 89 85 81 85 81 8b 7b 7d 7e 88 8d 6d 42 1c 0a 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 06 06 06 0f 26 37 58 79 8a 9f b0 bd b3 a7 9d a1 a9 ac a7 b2 b2 be dd f5 fe ff ff ff f1 eb e0 e1 e0 e1 e6 ef ee f6 f5
 fb f4 f6 f9 f9 fb f7 fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ed f2 f1 ed e8 ea e3 e3 e3 d8 d8 d3 d7 d6 ce d0 d4 d3 d4 d1 d0 d6 d5 d3 d1 cf d2 cd c8 cb d0 cd c3 c5 c5 c2 cb c4 c8 b5 b1 a4 a4 a7 9d a0 95 9a 9b 9f 95 9b 94 90 8b 88 8a 89 82 8b 80 80 80 7d 7c 75 87 7c 7f 89 67 39 17 04 06 05 03 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 08 0b 0b 1f 34 56 77 88 a6 be c3 c2 ad a0 a7 ab b6 c5 ca cd d5 d9 e7 f4 fe ff ff f9 e5 de de df e1 f0 e4 ec f6 ed f6 f3 f7 f9 fc fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 fb f3 ea ef eb de df de e2 dd d1 d8 c5 ce d1 c9 ca c8 d3 cd ce d1 d3 d1 c9 cd c5 d2 ce d0 cf d0 c9 c0 d0 ba c5 ba c7 c7 bd bb a6 a0 9f 9f 9c 98 95 98 8f 95 97 92 8f 90 93 87 85 84 7e 7a 80 7c 7b 7e 7d 7c 7a 85 7f 60 31 09 02 06 05 05 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 07 06 05 11 16 2d 55 75 8a ab c0 c6 c4 bb a3 a7 aa b5 c4 d1 db e2 da d2 dd e6 f5 fe f1 e2 d7 de db da e5 e2 e1 ed f2 f4 ef fa fe f4 fb fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f1 ef ec ea e0 de e1 d2 d5 d6 d1 dc cb c6 cc cc c6 c4 cc c8 c6 ca cb c6 d0 ce cb cd ca d3 c7 c6 c8 be c3 c7 c2 c3 c3 b4 c9 be bb b5 b0 a7 9e 95 9d 9b 9c 9d 93 95 94 95 91 96 98 98 87 80 81 78 87 80 7f 84 78 84 81 7a 7c 53 26 0b 06 06 05 03 04 06 05 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 11 12 14 28 42 63 81 a5 be cb cc c1 b7 b6 b3 af b5 c7 d9 e4 d9 cc cf d4 dc e1 ee e7 d5 d6 df d7 dd da e0 e6 ee
 ee ea f1 f3 f2 fb fe f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f7 f1 ef e5 e7 e2 e0 d9 d7 d6 d3 d2 d0 cc cd ce c5 bc c7 c2 c7 ca c8 c2 cd bf c8 c2 ca d2 cb c4 c0 c1 c3 be bc c7 c1 bc b5 b6 b3 ba bb b2 a4 a5 97 9c 95 96 94 9e 98 94 9c 9a 9a 98 8f 89 85 84 82 7e 83 83 7f 75 7c 7a 73 6f 67 40 27 07 04 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 0a 0e 29 40 5a 7d 98 b8 cd cc c2 b3 bd bc b7 bd c1 c7 db de c8 c2 ce ce ce db dd d6 d1 ce cb d1 db d1 dd e5 e8 e2 ee f0 ec f2 fa f2 fa f6 ff ff ff ff ff ff ff ff ff ff ff fd ff ff ff f5 fe ff ff fb ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f9 f5 f2 ea e1 e0 d7 d7 de d2 d6 cf cf ca ce cb c2 c3 c6 bf be c2 c3 bc bd c7 c1 c6 be bf c1 c8 c2 c8 c2 bb b7 b7 bb c1 ba b4 a9 ab b1 b0 b2 ad a3 99 9f 9b 95 8f 95 98 94 9a 98 8e 92 8c 90 85 74 80 7e 80 82 75 76 7c 6c 7b 76 6d 61 36 1c 09 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0a 05 0f 12 22 41 55 72 8c b3 ca d0 c7 bc b3 c0 be c7 ce d0 d6 e5 d9 c9 c6 ce d5 d0 cf d1 d4 d0 cb cb d2 d5 e0 e6 e7 e4 e3 e9 ed ed e9 f5 f4 f9 fe ff fe ff ff ff ff ff f6 f9 f9 fe fc fb ff fc fa fb fd f7 ff ff ff ff ff ff ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f9 f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb ef f0 e2 de e0 db da d5 d8 cd cf ce c0 c4 c2 bf c1 c3 be c5 b7 bb c2 c8 c4 c4 c7 be bf bb bb c7 c6 c5 b5 bb b5 be c4 bc bc ae b0 a4 ac b1 b2 a8 a1 87 9c 96 96 9d 9b 9b 9f 9d 95 93 88 85 86 80 7d 81 86 83 82 78 75 7a 79 76 70 61 4f 29 0e 03 03 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 13 1f 24 40 55 72 8d a6 bf cd c0 bd bd bb bd c4 c8 d3 d5 e9 f3 dd d8 d3 d8 d4 c9 cf d4 cd d1 d7 d2 d6 d9 df
 df e1 e5 e4 e9 e6 e9 ed f5 f9 fb f8 fa f8 fa f7 f3 f7 f6 f8 f9 f7 fb f8 f6 ff fa f5 f9 f8 f9 fc ff ff ff ff fd ff ff fa ff fe ff ff ff ff ff ff ff ff ff ff ff fe fd f4 ee ef ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd ff ea ee e6 e5 e1 e0 d9 da d7 d6 cd c5 ca ba c6 c8 c6 bb c2 bd c1 ba c7 bf c5 c2 c6 bc c3 c1 b6 c3 c0 c2 c3 b7 b0 b5 b1 b6 bf c4 b5 ac a5 ab ac ab a7 aa a0 a5 9f a6 a4 a5 a5 98 96 94 91 92 88 86 87 7b 81 84 7e 7b 7b 83 76 70 70 6a 63 48 21 12 03 01 06 05 03 09 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 10 08 0e 0c 20 37 4e 70 8a a4 bd bf b9 ad b9 b6 bc c6 c0 c5 d5 dd ed e6 e1 e4 df d6 d8 d2 d2 cc c3 cb ca d2 d4 d6 d1 d4 d9 df e0 e2 e5 e7 e0 e8 e9 f5 e6 ee f5 ed ee ef eb f2 f1 f1 f4 f7 fe f9 ff f9 f9 f9 fb f9 ff fa fd fa fd f9 fe ff fb ff fe fd ff ff fd ff ff ff f6 fb f3 f5 e6 ec df da df fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fa f5 f0 ec e0 e0 dd de de cd d3 cd d2 cc c2 ba bf bf c1 c0 bb c4 b6 b7 b5 c5 cb c5 c2 b7 ba bd ba bc bb bf c6 b0 b3 a9 b3 b9 c1 cb b7 be b2 a6 b0 a5 a9 ae b0 b2 b0 a8 a1 9e 94 8c 94 89 91 86 8d 88 8a 7b 80 7b 7b 83 79 7b 71 6f 6f 68 4e 2f 27 0f 0f 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 09 16 1e 43 55 71 8b a3 b0 c3 c0 b5 b3 c0 b5 bb bb c5 c9 dd e1 eb eb e8 e5 d6 cd c5 d0 cb c4 ce cb d1 d1 cf db d8 d2 da dc df e4 e5 e6 ed e5 e5 e7 e5 ea e6 f0 ed e3 ef ed ea f1 f3 fd fa f5 fb fa fc fc f9 ff f8 ff ff ff f4 fc f7 f6 fe f3 f8 f8 f3 ff fc f7 fd f3 f1 ea e5 de da d2 d5 e1 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe ff f5 f8 f2 ee ee da df de d4 d4 d4 d4 d1 cb ca c4 c1 c1 c1 ce c3 ba c1 b4 ba be c5 c6 ce cc c5 bf bb b9 b5 b1 b7 be b8 b1 af b3 ba be c4 be c1 bf b9 bb ac ad ab ad ae aa a0 96 95 92 8f 8d 94 91 8b 92 89 83 7d 7f 7e 7b 77 73 76 72 73 70 61 52 36 20 12 0c 0a 06 05 03 00 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 0c 1d 19 34 5d 68 83 9c b0 cc bf b4 b0 b2 be b6 b7 be c5 cb df e2 eb f4 e6 db d1 c8 ca c3 cc cc c5 d0 d5 cf
 d8 d6 d7 d7 de db e1 e2 dd ea db e0 e1 e6 e3 e5 e0 e8 e1 ea e9 ee f3 f4 f9 f3 f4 f8 f3 f4 fe ff f8 fd fb fb f7 f6 f3 f5 fc ec f7 f5 f2 f7 ef ee f4 f4 e9 e4 e4 db d4 d7 ce cd d3 de ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 f6 f1 f0 ec e4 de d7 df d8 d4 cf cf ce cc ca c2 c7 c2 c5 c6 ba c0 c1 b0 b6 bb bc c7 cf c8 cb c4 bb ba b7 ba bb be ba b4 b0 b8 af b4 bc c1 c9 b4 a7 a7 a7 a9 a6 a1 a3 a1 95 90 99 93 8d 8e 89 8a 8c 88 86 89 84 81 7b 7e 79 78 6d 76 62 6e 56 48 32 26 13 0b 03 06 05 03 02 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 08 0b 12 0e 22 35 57 63 84 a0 ac c7 be af b6 ae b7 b5 b7 b6 b5 c6 d2 dc eb e7 e5 e0 ce c6 c0 c4 c7 c2 c9 c2 cc c8 d2 d6 de d5 d3 d5 dc da e0 e2 da db df da de e0 da e0 e1 e3 de eb ed f2 f2 f0 f5 f4 f2 f6 ff fc ff fa f2 f7 f3 f2 f4 ef f0 f1 ea ec ea ee ed f1 ee eb e4 e3 d6 d2 d3 cf ce bc d0 d9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd f1 ee eb e3 e2 e0 d8 db df d4 cf cf ca c5 c8 c5 c7 c2 c3 c3 bb c0 b8 b9 bc b8 b2 b8 b9 c7 cc c9 b7 b1 ab bf b2 b4 bb b5 b5 b1 af b5 b9 b9 b7 b6 a0 9f 9f 96 a4 9d 9c a5 94 97 97 8e 8e 90 89 8a 92 87 94 84 87 83 7f 85 73 74 79 70 68 66 6b 56 50 3e 27 1d 18 00 06 0a 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 0f 1a 26 3e 52 68 7c 97 b4 c1 c0 ad b4 ae b2 b6 b8 b2 b4 b7 c9 d2 db e1 cf d1 ce cb cf cc cd ca c6 cb cc cd d1 ce ce d5 d2 da d5 d5 d0 cf d5 d0 d3 d9 d8 d6 d9 dd e7 ea e4 e6 ef e7 f8 f1 f7 fa fa fa f3 f8 f2 ef f6 ed f2 ee ea ef eb ea ef e9 e9 e5 e8 eb e8 de e0 db d4 d0 ca be c1 c9 c4 d1 f0 ff ff ff ff ff e7 e4 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc f1 f7 f8 e7 e8 e6 e0 d9 d0 d3 cd d5 d0 d0 cc c6 c6 c6 c8 b8 ba c2 bd b7 bf b8 ae b5 be b1 c1 cb c6 c0 b6 b6 be b0 b1 aa aa b2 b3 b5 b5 b3 a9 ac af ac a9 9c a6 96 9e 9b 9e 9a 95 96 96 9b 92 91 83 85 89 8f 8b 86 82 7b 84 7c 74 7a 6e 75 70 6a 67 57 55 49 33 25 0d 01 08 05 03 00 06 05 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 10 1d 2f 44 50 71 85 9c b2 c2 c8 ad a9 b3 af b4 b4 b6 b8 bf c8 cc d6 cf bc b4 b8 bd be c4 cb c5 cd c1 ca d0
 cd cd cf d2 d5 c8 d1 c8 ce cd cf cf cc d6 cc d9 da df ea e1 e5 ed f0 e6 f2 f3 f1 f3 f5 fc ef f7 ef ea e9 ef ea ea f0 ed ec e7 ea e5 e7 e5 ea e6 e9 d9 dd d5 cd d1 c5 cb c5 c0 c4 c8 de ff ff ff ed e1 d0 c1 d8 e4 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fa f2 f3 ee e9 e4 de e2 d5 db d2 d2 cf d1 cb ca cc c6 c3 c1 be be c3 c4 c5 bf c2 b7 b2 bc b4 bf bf bc bd b5 bd b7 b8 b4 ad af b0 b0 aa ae b1 a1 b2 a6 a5 a5 a3 97 9c 97 a0 95 97 93 95 8a 85 87 8d 87 88 88 81 8a 7e 7d 78 7a 78 79 73 79 77 74 6b 5e 66 5d 4d 36 26 17 07 06 05 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 1a 31 3d 56 73 82 9a ad bd bf b0 a9 a9 ab ac a6 a9 b5 c0 cf cc c7 b7 a6 a1 a4 aa b3 b0 c1 bd b8 c3 bf c2 c6 c9 cf c7 c4 c9 c4 c7 d1 c9 cf cd ce ce cf df d7 dd db dd db e5 e9 e4 ea e6 f1 ec f3 ea e4 e8 eb e4 e6 e3 ea de dd e8 e4 e2 eb e9 e9 e0 e9 e5 dd db d4 d2 c2 cb bd b5 b9 b6 b9 b7 d9 fd ff ea d3 ca b6 b0 b5 c2 cc da f0 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 fe fb f9 ef eb eb e6 e1 e1 e0 df d9 d7 c7 ca d0 d1 c9 bf c4 c1 b7 b7 bf b7 be be b8 b4 bd b2 b3 b8 b3 b7 b7 c1 bb b6 b1 ba ab ae ad a6 a6 a7 ab a6 9d a4 a1 a8 a5 98 a1 92 9c 9b 94 9d 8e 8a 8c 89 8a 87 86 8a 8b 87 80 7d 84 7d 7c 77 77 74 74 75 71 71 67 73 6b 5a 4e 2f 25 1b 0b 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 0a 18 20 39 4d 5f 7a 89 a2 b5 c3 c5 af ae b1 a8 ba ad af b5 bc c4 bd bd ab 97 97 a0 a7 ab aa b3 b2 b5 ba bb b8 c0 bf c3 be c9 c6 c0 c3 c7 cb cf ce cc d2 d1 d6 d5 d4 d8 dc dc df e8 e8 e3 e1 e8 e8 df df e2 e9 e7 e4 e7 e7 e2 e4 de e9 e5 e4 e0 e5 e2 e5 e7 e2 e3 d2 d2 d1 c9 bf b6 be b6 b8 b8 bc c7 df e4 c6 b3 a1 92 95 95 9b ab b1 b8 c2 c9 d9 da df ea ef ec f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f8 f0 f1 eb ec e7 e4 e5 e0 df dc d2 d4 cd c5 c9 c7 c6 c9 bf bf c4 bd bd bb c1 c2 c7 b5 b9 bd b1 ae b4 b3 b8 b5 b1 b5 a8 b0 a7 ad ab a5 aa a5 a0 a0 a2 a1 9e 9b 98 99 9b 9a 9a 99 9e 95 92 8a 8a 84 83 82 85 8a 81 86 7f 7a 80 80 7e 75 7f 73 6f 76 70 77 6e 6f 79 7c 6c 53 42 2c 20 0a 06 05 04 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 21 27 34 52 68 74 97 a2 b5 c9 c3 b1 b2 af a7 ac b3 b3 be c5 c2 b0 af 9a 8d 85 95 9d 9f a3 a6 ac aa a8 b3 b6
 b6 bf be be c6 be c3 ce c6 ce d0 cb d0 d4 d8 d5 d4 cf da da dc d8 da e0 e0 df e6 dd d7 e1 db e1 e1 d9 e1 e0 dc e0 df e1 e2 e0 e0 e4 e8 e5 de dd db d7 d2 c9 c2 ba b8 b4 b7 b4 b3 b5 b6 d1 cd b9 9c 80 76 71 75 74 77 7d 84 89 8f 9e 9e a6 af a8 aa ba cc de f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 f5 ef ea eb e3 db df e2 d7 d8 d3 d2 c9 ce ce c6 c0 c6 c3 cb bf be b9 bc ba b8 bf bd c5 b3 b4 b3 ab b8 a9 ab ae b0 b3 ab a9 b0 a7 a9 a3 a3 a1 a6 99 a0 a0 a1 9d 9e 96 9b 92 97 98 94 8b 8a 8e 94 8b 86 82 83 87 86 84 80 8a 80 85 76 75 75 77 7f 74 78 6e 77 78 7b 83 7e 72 59 4d 31 21 19 0a 05 08 06 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 09 1e 2b 33 51 66 85 9a ab b7 c7 bd ac aa a6 a1 aa af b0 be c6 bc a5 9c 8c 87 8c 93 98 91 90 a0 9b a3 a8 a7 a9 b8 b3 c4 b7 bf be c8 c3 bf c6 bf c2 cb ca c9 d0 cd cb db d7 de d6 df d6 da dd e1 d7 db db dd e6 e0 e2 d8 e4 e1 e0 dc de e0 e2 dc e4 df e6 e6 e7 dc d4 d2 ca be b4 b9 b7 b1 af ae b1 b0 c5 bc 9c 81 68 55 57 51 59 53 5c 59 60 63 67 77 71 7d 80 7d 80 8c 99 a5 b7 bd cd ea db ff ff ff ff ff ff ff ff ff ff ff f4 fe fc fe ff ff ff ff fb ff ff fe ff f2 f3 e7 e8 e9 e0 db d9 d3 d7 cf d5 cd cc c9 c7 c0 c4 c4 be b6 b8 bf b5 ba bb b5 b6 bd b5 b5 b4 b4 b7 ac af b4 ae ab ab ac a6 ad a4 a1 a6 a0 a3 9e 9b 9a 98 99 94 9b 9a 93 99 8e 8f 87 8e 84 87 8d 84 83 85 80 7f 7d 7f 7c 83 80 7a 7d 7b 77 72 76 77 77 74 73 75 76 7a 84 78 72 5e 4b 3c 26 1a 0d 08 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 12 17 24 27 3a 50 68 7e 92 b3 b7 c6 be a6 a8 ac a1 a8 a0 ab b5 b3 ab a0 8c 81 81 80 8c 8f 97 9a 90 9c 9e a2 a6 ad ae b0 b5 b4 bc c8 c1 c2 be c0 bd bc c7 c7 ca d1 c9 d5 d0 da d1 dd e0 dc e3 de d5 d9 d6 db d5 d1 de e0 db d8 d8 d6 e1 d6 e4 e4 e0 dd e3 e0 e2 df df d5 cb bf be bb b5 b5 ad aa a9 ac aa b0 b3 91 68 56 4b 4c 4a 4b 49 4d 49 4b 4a 4d 52 54 50 60 5d 63 6d 6c 79 79 7b 89 99 ae be cd e3 ff ff ff ff ff ff ff f2 ec f0 f8 f3 f3 f0 f6 f5 f5 f5 f8 f1 f1 f5 ee d6 de de d6 d6 ce cd c7 cc c1 c4 c5 c4 be be be c1 bd bc b9 bb bd b6 b5 b3 b9 bc ba bb b6 af a7 a7 ad a7 a7 a5 a0 a7 ac a5 a3 a3 a1 9a 98 91 9c 93 98 a4 a4 9d 91 89 92 90 92 88 84 83 86 83 83 81 77 80 7d 7d 79 81 7f 7e 7e 7a 7c 6f 78 76 75 75 71 7a 74 7c 6f 83 7e 6e 64 43 3a 24 1d 14 0e 03 03 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 11 1e 2a 34 4c 61 6c 7c 9f b1 c1 cf b8 af 9d a1 9f a3 ab af b4 a8 a0 9d 8a 84 7d 7f 80 8c 94 99 9e a6 a5 a8 a6 a7
 b0 ae a9 b4 a9 b1 b9 b3 b9 b8 bb c1 c2 c8 c8 ce d7 d2 d7 d8 d5 d9 e0 db e0 d8 d6 d4 db d3 d4 d8 dd db df e4 e4 d9 db d7 e1 db e0 db df df d8 da df cf cd c4 c2 b0 b9 ba a9 a5 a5 a9 ab b3 9f 80 5d 50 41 3a 42 3e 3f 3e 36 3b 3e 3a 40 46 4b 51 49 4a 58 59 60 65 61 6d 74 77 83 8c a2 d3 ff ff ff ff ff f6 e9 e0 de e8 e7 ef e9 ee ed f2 f3 f2 f0 e0 e2 e2 e5 d3 db d0 d3 cc c2 c7 c7 c2 be c7 ba c2 c1 bc b9 b5 bb b3 b5 b0 b3 af b7 b6 b6 b5 b6 b6 b8 b7 ae a2 a5 9e a8 a7 a3 ae a2 a0 91 98 9b 9b 98 96 92 a0 a3 9e 99 94 91 92 85 8a 89 84 91 81 85 82 7f 84 81 7b 80 7a 79 7f 85 81 81 74 73 7a 7c 74 71 72 74 70 7b 74 7b 84 77 6e 5b 42 36 27 1a 0f 08 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 07 0d 0a 26 24 3a 4d 59 6f 89 a2 b0 c7 c8 b6 a6 a1 98 9b a4 9c ac ad a4 97 90 85 84 81 8a 83 8c 8b 8b 99 9f 9f a1 9d a1 a5 a3 a6 a5 a2 a7 a9 b5 b6 bc c3 c2 c1 ce c7 ce d7 d3 d8 d1 d4 cf d7 d1 de da d4 d7 cc d0 d6 dc dd dc d9 d7 dc d3 de df e1 df db dc de dd da d8 d7 cb c8 c0 b8 ba b3 b5 aa a9 aa ad a0 a2 94 74 56 47 3f 35 3d 32 3e 34 30 30 32 30 34 3b 3a 3d 41 49 4e 55 52 4e 53 5b 62 58 68 6a 7e a0 ee ff ff ff ff ec cf dc d3 de db e9 e1 e8 e6 e8 e4 df e4 e3 e1 e1 db d6 d0 cc ca bd be bd b7 b9 ac bd b4 b9 b8 b3 ba bb b5 b8 ae b5 b6 b2 ad af b2 b3 b5 af b1 af ad a4 a2 a0 98 a2 aa ab 95 96 92 94 91 8f 94 92 92 98 9b 9c 96 90 85 88 86 7e 85 82 87 79 76 84 77 7c 80 7d 79 78 7a 7d 75 75 78 77 78 70 79 6f 70 76 77 73 75 6a 7d 7c 76 6c 58 46 30 29 14 13 09 10 0c 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 12 15 1a 27 3d 47 5c 79 89 a4 b3 b8 ca b6 a3 9d 98 a1 95 a3 aa a2 96 8c 86 7e 7b 78 7f 80 86 87 90 94 96 8e 99 97 9a 9b 96 9e 9c 9e a0 9e b2 b7 b6 b4 c3 c2 c7 cd cc d2 d0 d1 d5 d0 d5 d4 dc dc da cb d6 d3 d2 da da d4 d8 d6 e0 da db d5 d7 e0 d4 dd da d5 de d9 dc ce cb c2 c1 be b7 ae b8 ac ab a5 ab a6 a5 9a 69 51 3a 29 37 25 2a 2c 32 22 2c 22 2b 27 2f 36 37 35 3b 37 3e 42 3a 42 4f 4f 56 57 55 62 84 bb fe ff ff ff d5 d1 d0 d0 db d8 da d5 db d9 e0 d5 d5 d5 e0 d8 d7 ce d0 cf cb ca b8 b8 b7 b8 b4 b2 b2 ae ae b3 af b1 ab ad ae b0 ae a7 b5 b0 aa ad a0 b3 a7 ad a5 a9 a6 a3 98 96 ad a5 9a 8e 93 92 91 95 8a 95 91 8f 93 93 95 8b 87 84 7c 7b 85 81 7d 80 7c 81 7b 7f 7a 81 77 7d 77 7c 79 73 76 6f 6f 70 70 77 7c 78 75 74 71 6a 70 73 7c 76 6b 5e 4d 45 34 21 17 05 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 08 06 0e 1f 25 31 3e 48 5f 74 86 ac b5 bd c8 ad 9d 92 9c 9d 9c a0 9c 85 84 7b 7d 7e 77 84 7a 7c 7c 88 83 88 90 8d 93 8d 94
 94 94 94 9c a1 a2 ae ab ae ba c0 c3 c8 c5 ca d0 c9 c4 cb d4 cf d3 da cb d5 ce d1 d0 d3 cd d3 d9 d6 d7 da d5 d5 d8 d6 dc db d7 dd de d6 e3 d7 d7 d6 c6 c2 c3 b3 b6 ad ab a5 ab a7 a5 a0 9c 8e 66 39 32 2f 23 26 2a 26 25 2a 22 25 24 23 2b 29 28 2c 33 31 33 36 3c 3c 42 47 44 4d 55 56 73 95 cf ff ff e5 c6 c2 c1 ce ce d7 d4 d0 da d7 d5 d4 d0 cf d3 d2 d4 c8 cb c2 c6 bb b8 bc a9 b3 b1 aa b1 a7 a7 a3 a8 b2 b4 b3 ad a9 ac af ab ab ab ae b0 b8 a3 ae b0 a4 a4 9d a1 9f a4 a3 98 8e 90 8d 8e 91 8d 90 88 85 8d 96 96 8b 84 7c 83 7e 7f 7e 7c 80 79 7a 83 79 77 76 74 7c 76 75 6f 74 69 7d 75 7c 78 7f 78 75 7c 79 65 67 66 6a 7b 78 76 69 56 46 32 32 1c 17 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0b 12 0a 1c 31 2a 41 56 67 7a 8b a2 b9 be c2 aa 8c 8c 90 8d 8d 91 90 81 84 73 70 7d 75 73 79 7a 7d 89 8b 8c 91 92 8e 8f 9d 9a 9d 9d 98 a1 a8 ad a4 c0 b9 b5 c0 c9 c6 cc d0 c5 ca cf d2 d3 d5 d6 d2 d1 ca c7 cd cf d2 d6 d5 d7 d9 d2 d9 d8 db d6 d5 dd e2 d8 df e0 dc d1 d6 d0 c3 c2 ba b8 b6 a8 ad ab a1 a6 a1 9f 9c 8d 61 41 2e 1c 27 1b 1b 23 23 1b 21 1c 23 1c 25 1c 29 27 24 2b 2b 2d 2a 27 2e 3e 3f 44 48 51 62 86 aa dc de c1 c3 bc c2 c2 c0 c6 c8 ca d0 c6 ce cb d2 cc d3 cc c2 c2 c3 b7 c0 b6 b6 b0 b2 a6 a2 af a7 aa a6 a2 a8 aa a6 ab a5 ab a1 a4 ab a9 ad ad a7 ad a7 b0 a9 97 98 a2 a0 9f a0 95 94 90 81 86 8d 8e 90 88 88 86 8c 8c 8f 8d 7d 83 80 7c 7f 82 7d 7b 7c 7d 7b 7b 80 82 72 76 7d 75 82 7f 75 82 80 77 78 6f 7e 76 7a 71 67 69 66 69 73 71 74 68 57 46 3c 2b 21 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 07 08 1c 25 2c 41 47 58 6c 79 8d 9e b6 b9 ba 94 88 83 7a 89 89 84 86 74 83 75 76 72 7a 7b 76 7e 7d 78 85 89 90 8d 90 93 90 96 9c 93 a0 a7 a3 a4 ab b0 b6 b5 bc c0 c3 c6 c4 c7 d2 cc d5 d4 d4 d6 ce d1 c9 c9 cc ca cf d5 d0 d7 d3 d5 db cb d6 d7 d4 d8 d7 d1 dc d8 dd d5 d7 d0 cc c2 bd ae ac af ad b4 a4 a3 9a 9b 95 7d 44 32 28 1a 1a 19 20 21 19 13 10 1a 14 16 14 1a 1e 1f 1d 1f 24 29 24 29 29 34 3f 36 46 43 59 7f 90 bc c2 bd b5 b6 bb bc c1 c3 c6 c2 c5 c1 ca ca c5 c3 cb c3 c5 c0 bb c2 b7 ad b1 af ac a4 a5 a4 a6 a3 a5 a3 a6 a3 a9 ad af b1 aa a5 ab a7 a3 a3 a5 b2 a1 ad a8 a0 9a 9e 9a 9d a1 95 8c 8a 88 8a 8d 80 83 86 8b 88 85 8a 83 80 80 7f 7c 74 7b 7b 79 7e 6d 78 7e 7d 78 77 75 80 75 7f 86 7c 7b 78 79 6c 79 72 6f 7b 6f 6a 60 5c 66 5f 72 71 75 6c 5f 5a 3e 2e 24 13 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 08 16 14 20 2c 37 4e 5c 6f 85 a0 a9 b6 ab a7 86 84 73 77 7e 73 7b 79 79 79 7a 79 79 78 72 73 81 79 82 8b 8b 89 95 90 98 94
 98 9c 99 9e a7 ad a8 b5 b0 af b9 bc be bf c2 c5 c4 d0 d8 cb d0 d4 d1 ca c9 cd ce ce d3 d5 d2 d4 d2 d8 d5 d2 d0 d0 d1 d0 d3 d6 d3 d9 dd d9 ce d3 d1 c7 bd ba ae b0 ad a6 a6 9b a4 9b 96 8d 71 40 30 1f 17 2b 19 14 1e 14 13 14 19 1b 13 18 17 14 19 15 1a 1e 23 21 25 22 32 3b 36 39 37 60 83 90 aa ac b8 b4 b0 b4 af b4 b7 be c1 be c2 c6 c6 c5 be c1 b2 ba b3 bd b5 b5 b0 ab aa a9 a1 9f 9b 9e 9f a0 9e 9d a1 9f af aa b3 a7 a2 a5 a3 a2 a7 a3 ae a5 a5 b0 a8 9d 95 98 9f 9c a4 99 85 84 85 90 85 8a 88 81 81 88 87 80 82 86 84 7d 7b 74 7c 81 77 82 79 80 7d 76 7d 76 85 82 88 80 7c 78 7e 71 76 74 7d 77 6c 6d 68 5f 60 5f 5b 65 71 78 76 62 4c 44 32 24 12 17 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 03 06 0a 0d 11 1d 34 42 4f 5c 73 80 98 b9 b6 a9 8b 74 76 75 71 75 67 6d 77 72 79 77 73 7b 76 77 7d 76 79 88 7f 8d 8e 8b 90 99 99 98 a1 9e a4 a9 a0 a6 ac ba b6 b5 bd be ba c2 c9 ca d5 d1 d9 cf cb cb c8 ce c9 d1 cf ca d7 d3 d4 da d0 d0 d6 cf d8 d1 d3 d8 d0 ce d8 d2 db d6 cd c7 c1 ba c0 af ae b0 a6 a1 a0 9c 99 93 8b 69 44 27 18 16 1a 0e 0e 15 1b 17 0f 17 14 12 15 17 19 11 14 1a 22 19 1e 18 21 2b 32 36 2c 3c 50 80 9b a9 b0 a7 ac aa b0 b8 b5 b6 b9 b9 bb bb c4 ba ba b9 c0 b6 b9 b2 b4 b8 ae ac a7 a5 a8 99 a0 9e 9b 93 9a 96 8f 9c 98 a5 a8 a7 a9 a6 a5 aa a2 a6 9f a7 a1 a6 a6 9c 9b 9c 9d 9a a0 9d 92 8f 8b 8b 8b 86 85 89 86 84 7e 7a 82 80 84 7d 81 7a 87 78 80 7d 78 80 80 7e 7a 7e 79 7d 7f 76 7e 7c 72 7b 6b 70 71 6f 72 6c 65 64 65 61 5d 55 5f 6c 7a 72 73 63 4f 39 2c 19 17 09 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 05 11 1a 2f 35 3f 51 62 78 8a 9e ac b7 95 81 76 66 78 71 68 6d 6a 76 79 7a 7a 74 7d 77 74 73 81 8c 7b 8a 8a 8d 88 8f a2 9f 9f a2 a6 a2 a5 aa ab a5 b3 b2 b2 b4 bb c2 c9 c7 d0 cc d3 cd ca cd c2 cb cd d1 cf d1 c8 c5 cd ce d5 d1 cd d4 ce cd d7 d1 d0 d4 ce ce d8 c9 d1 d2 cd c5 be b9 b2 b2 a9 a5 9f 9f 9e 99 95 8b 66 34 1f 16 10 0b 07 0b 0f 10 0d 0d 09 0e 0f 0b 15 16 13 0f 10 15 12 11 16 1e 1e 23 29 29 33 4c 80 9b a1 a0 9f aa a5 a7 a5 b0 b0 b2 b7 b6 b2 af b5 bb b5 b0 b4 b2 a7 ab a6 a6 a8 a0 a1 9e 99 9d 96 99 8f 93 8d 8f 8d 99 94 9f a7 a2 9c 96 9d 9b 9a a3 98 9f 9e a6 98 9d 9b 8c 92 98 94 94 8b 87 89 86 84 84 87 7a 7a 81 7d 82 88 7e 83 84 7f 84 7a 81 7e 84 7f 7f 77 79 7d 7d 7d 81 7b 71 73 76 72 76 77 75 71 6b 62 63 68 64 5d 57 5a 53 5d 70 76 6b 5a 54 3d 2d 1f 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 11 17 25 34 42 55 65 7d 92 9e b1 ad 84 76 6c 71 73 6f 6e 70 70 73 72 77 7a 77 7d 74 73 79 7d 83 7e 84 81 93 93 98 a7 96
 9e a1 a0 9e b0 a3 b1 b1 b4 c1 b0 b7 c8 c8 cc c7 ca ce ca cb c5 c1 c8 c3 cb cd d2 d5 ce d4 cf c9 d3 d0 d3 d3 cf d0 d5 ca db d5 d6 d5 d8 d3 cb c7 ca ca c0 b9 b2 a6 a4 a8 a3 9b a5 94 8f 87 69 3c 2a 18 0b 05 14 0c 19 13 14 09 0d 0f 0d 15 11 0f 0f 0c 1a 1a 15 11 12 1c 28 25 22 35 2c 4d 87 9e a7 99 9d 9f a3 a2 a5 a5 b4 ad b0 b1 b2 b1 b9 a7 b0 b0 b1 a8 aa 9f 9f a7 a2 a7 9e 9e a0 90 8e 93 92 8a 90 8d 8b 8e 94 9f a9 a3 a2 9e a1 9d 96 9d 9a 99 a1 9e 99 91 94 9a 94 91 93 91 8d 88 8c 80 8c 81 7d 7d 79 7c 7c 84 81 82 7d 7d 7a 7a 83 7c 83 7d 81 8b 7f 7d 7c 71 7f 76 7a 78 77 7a 73 79 74 6c 6d 66 62 61 62 62 5d 56 55 56 54 67 7c 70 67 5b 47 2c 1c 1d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 13 16 29 35 47 53 6b 79 8e 9e b0 a9 91 7a 73 67 72 6e 78 76 6d 73 73 73 78 73 6f 77 7c 76 85 84 8a 86 87 92 91 91 9d 9d a2 a5 a5 a7 a5 ab a5 ab b4 b0 ba bb c3 c6 c9 c8 ca ca ca bf bf c3 bb c6 c7 c8 d1 d0 d2 ca cd cb d0 d2 d3 d3 cd cf d5 d1 d8 cf d9 d4 cc d3 cf ca cc b5 c1 b4 bf b0 a7 a5 a6 9e 9a 94 91 8d 79 4f 24 1c 0c 0a 09 0b 0e 05 06 0a 07 0c 0f 0a 0e 0d 12 0f 11 10 15 09 1c 15 1f 21 21 23 2c 3e 80 92 97 9b 99 9b a3 a1 a7 ac a9 b0 b4 ae a6 ae ae a7 a7 a9 9e ab 9e a0 a2 9a a3 a3 98 9d 92 9b 91 93 90 8c 93 90 8e 92 95 9c 9e 9e a1 9c a3 9d 95 9a 9e 95 96 9d 8e 8a 94 8d 8d 90 8c 8e 8f 89 84 8e 8a 84 83 80 7f 77 80 81 7d 85 80 78 80 89 7b 82 7e 85 76 7b 78 7e 7c 76 77 79 81 7d 72 72 75 73 73 69 68 5b 5f 63 60 5e 5e 62 51 59 5c 65 77 76 6d 57 50 36 24 1d 0c 06 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 05 12 23 2a 39 52 52 64 71 88 9f a6 a0 91 79 72 75 73 73 6e 7a 6e 66 75 73 72 7b 75 74 74 78 7b 7f 84 88 8e 94 97 8e 9a a4 a2 9f a4 a7 a5 ad a6 b2 aa af b9 bc c1 c5 cb c5 c4 ba b5 bd bc c5 c1 ba c3 c3 c5 c6 c6 cc cd d2 cf c8 cd cc d1 cd ca cb d4 c7 ce d0 c9 d1 cc cd cc c1 b9 b9 b1 a9 a9 a3 9f 99 99 90 8b 84 78 49 18 0f 0a 09 0a 0d 0d 0b 0c 07 06 05 0a 00 0c 09 0a 04 07 0c 12 0c 18 14 12 1d 1e 1b 29 39 78 93 97 8f 94 97 9f 99 a7 a0 ad a2 a1 a3 9c a6 a2 a2 a3 a0 a1 96 98 96 97 a0 99 93 91 8d 93 92 8d 92 89 88 88 89 89 8a 92 99 98 92 9e 9e 98 98 9b 8e 97 8f 89 98 8f 91 91 8f 8d 89 8b 8c 80 8f 81 81 84 7d 7f 7a 71 7c 78 82 7b 7f 81 82 7f 82 7b 7a 7c 7c 7d 79 77 7b 74 6f 6f 72 77 7a 6d 72 70 70 67 66 61 5b 5c 5f 5b 58 53 59 4e 50 52 58 77 79 6f 60 52 3f 23 15 0f 05 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 0f 18 27 3c 50 56 62 79 8e 99 b7 aa 90 7b 6c 6e 7d 72 76 73 71 6d 74 6f 7f 78 73 76 78 7e 7b 85 81 85 86 8f 90 9f 9f 9b
 a2 a6 a8 a6 b0 a2 ae a5 ac b6 b4 bc c6 c2 bb bd b7 b4 bd b6 c5 c2 be bf c4 c6 c6 cc c6 cf d2 d4 cf ce cf d1 d2 cc cc cf ce cf ca d0 d0 cb c8 c4 c5 c9 bf b5 ae b0 a3 a3 9b 99 9e 92 87 8a 74 45 10 0c 06 05 19 05 13 0e 04 03 07 12 05 04 0c 0e 0c 0b 07 0a 06 0b 0a 19 19 1f 1d 22 25 3a 7a 94 91 9c 97 96 9a 9d 9e a5 a3 9a 9b a5 9d ab a1 9f 9d 99 98 9c 92 8b 93 8c 96 99 93 96 94 8e 89 8d 91 85 8d 8d 87 90 96 8e 9c 9c 9f 93 98 90 92 8e 92 8d 92 96 93 8b 8b 8c 89 89 82 8a 8a 8a 80 84 81 87 7e 77 75 7c 7a 75 7d 7d 7d 7d 76 83 7c 7e 7d 7c 77 7c 77 74 73 75 74 6e 78 76 74 74 72 69 66 5d 60 59 5d 60 5b 5c 59 52 53 53 54 5b 68 7d 6e 60 4e 37 26 18 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 14 1f 30 46 49 5f 65 7c 92 a5 ab a8 85 73 6a 6e 79 75 79 7d 79 6f 6c 76 75 75 70 75 73 78 89 84 81 91 91 9a 98 9e a4 a5 9d a0 a7 a5 ac ab a5 ab ab b1 bb bb c0 b5 b5 b3 b8 b0 b3 b5 b2 be bd bd c4 c2 c1 c8 c9 c2 c9 cc c9 c5 d0 d0 cb c7 cb c9 ce d0 c9 d1 cd d2 c7 c6 c8 c1 c4 b6 b2 af a4 a5 a9 95 98 8f 8c 85 75 50 25 0e 06 07 08 04 06 0e 03 08 08 07 0a 05 06 0f 03 04 06 0e 11 0b 0e 0e 1c 20 1e 29 22 2a 6d 85 89 9c 91 9c 9a 9b 98 9a a5 a2 9d 99 9b 9f 9c 94 9c 9f 9f 9d 93 8d 8f 96 90 91 8d 8c 8e 90 95 89 8b 8d 87 90 81 90 8f 97 9c 98 9c 99 92 91 91 94 93 8d 93 99 90 92 90 93 87 85 91 85 86 80 84 7e 86 85 7d 7f 7f 7f 85 7d 7b 82 81 7b 7b 7d 7a 7d 7f 79 7a 7a 78 79 75 75 79 75 77 7b 75 74 6f 65 61 61 62 65 58 5d 5d 54 54 50 4d 49 55 5c 60 7b 76 5c 50 3b 29 1f 0f 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 05 10 22 2a 43 55 61 73 7b 92 a3 a9 ab 86 7a 6d 74 78 79 7b 7e 78 71 77 71 74 77 77 70 73 77 80 88 88 8e 92 97 93 9a a0 9e 9a ab a1 9f a8 ad a5 ae b5 b6 af af b1 af a9 ac b1 a8 aa b4 b5 b8 bb c2 c1 bd c0 c4 c6 ca c9 c6 c8 cf c9 cb cb c6 c7 c8 c7 c4 c1 c9 cb c4 ce c7 c9 c0 bb a7 ad b0 a2 a3 a1 94 94 8d 7e 82 7f 60 15 09 06 05 15 03 06 09 04 08 06 05 0c 01 06 05 03 08 06 0b 0f 06 16 14 19 1a 1a 1c 1d 2f 5b 8b 92 98 94 9e 97 94 99 9c 9b 9f 9c a2 9d a0 9a 96 97 97 90 8f 8d 94 91 90 98 93 8a 8b 86 8b 8d 8a 8d 8e 89 86 92 91 96 97 91 99 8d 91 91 8b 92 8a 8b 83 89 96 8f 90 90 80 83 84 85 8b 7a 7b 7e 7f 77 86 76 79 74 75 81 7e 7c 7b 81 7f 7a 7a 6e 7a 77 7d 77 76 78 75 78 76 72 6d 74 77 71 6f 63 63 5f 61 60 64 55 54 58 54 57 4d 54 4b 4f 57 5f 7c 76 6d 55 3f 2a 1e 0e 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0d 1f 25 30 45 49 5e 6e 84 8f a3 b2 a9 8b 74 6d 70 73 77 78 73 7a 7f 7f 78 76 72 74 75 7e 7c 83 84 88 8d 93 93 99 9a 95 a1
 9d 9c a3 a0 9f a4 a4 ab ad ac ad a5 a8 a9 a7 ad ad a1 a8 b5 b0 b9 b8 b0 c2 b3 c3 bc c3 c3 c2 c1 ca c7 c6 c7 bc bf ca c1 be cb c9 d2 c8 cd c4 b8 c4 bb b8 b7 b5 b2 aa a2 99 95 8f 8b 8a 7c 7f 60 23 0d 06 05 0a 05 0d 08 04 01 06 05 05 03 07 0c 0d 00 09 05 05 13 0f 05 10 14 0f 16 18 2a 58 84 91 8a 91 8c 94 94 99 96 a0 9b 92 97 97 9e 91 8d 8c 8f 95 90 91 86 93 92 8c 85 8f 96 8b 8e 7f 8d 86 8b 89 8a 98 8b 90 93 94 96 90 93 90 8e 88 94 8c 8d 8e 8c 8b 82 87 85 87 8c 7f 87 7f 85 7e 84 7f 76 7d 7c 75 78 7e 78 7e 7a 76 7b 73 7c 7b 79 7c 78 7b 71 7c 65 6b 74 6c 65 73 6a 5e 68 69 5a 60 60 60 5d 55 60 5c 57 52 51 4a 4d 52 57 5c 70 77 6d 57 45 30 21 0e 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 20 20 3d 4c 53 5b 6b 84 8d a7 a9 a7 8c 6f 6f 6c 6b 73 76 7b 73 7a 80 77 77 78 78 79 79 81 84 84 87 8c 92 94 93 99 9b 9d 9d 9f a1 9d a8 a9 b0 a6 ac a8 a8 a5 a2 a5 9b a0 a6 b2 b0 ae ad b0 b2 c3 b8 be c2 ba be c5 c2 c5 be c4 c6 c4 c4 c4 c4 c2 c4 c3 ce c9 cc cc bd c0 c4 b7 b5 b0 b1 b2 a4 9e a0 9b 93 8e 89 7f 79 63 21 0a 06 05 04 04 0d 07 0a 05 06 05 03 07 06 0a 07 05 06 09 0f 0a 0e 0e 10 14 17 19 18 1f 4b 77 8a 8d 8e 92 95 9a 90 90 97 98 95 94 92 9b 95 94 91 8c 8a 93 86 8b 8c 8a 8f 87 89 89 88 87 87 93 89 89 8e 88 93 99 99 90 91 90 88 91 90 97 93 94 95 8d 8f 8b 88 8b 8a 80 89 7f 8c 83 83 86 7f 80 76 7b 7f 7d 7b 72 7b 7b 7d 82 7d 7d 70 7c 79 7a 73 75 70 72 6d 6c 6c 70 6c 6f 6a 6c 68 6b 6d 63 64 5e 66 5e 5b 57 53 57 5f 55 59 55 4c 57 5a 6f 77 67 55 44 36 2a 0e 07 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 11 1d 27 34 46 53 66 70 82 89 a4 ad b2 84 74 69 6b 73 74 75 75 74 77 7f 7d 7e 77 7b 7c 7e 7b 84 84 88 92 8d 95 97 8f 95 95 95 95 9d 9b 9b a6 9d a4 a8 aa a4 9c 9f 9f a6 a4 a7 a2 aa aa a9 af b3 bb b4 ae b9 b9 ba b2 bc c1 c2 c1 b8 bf be c7 b4 c4 c3 be c1 c5 c4 c6 c4 c3 c2 ba ba ad ab a6 a3 a1 9b 91 95 8a 86 8b 7b 5e 22 0b 07 05 03 08 06 08 03 0a 08 05 03 00 06 06 04 06 06 05 08 0b 06 09 09 1e 0c 15 17 1a 3f 79 84 90 93 87 83 89 95 94 95 8f 93 93 90 90 8e 90 8f 8e 90 8d 8c 85 88 8d 8d 8a 8b 8f 90 8f 86 91 86 91 90 83 95 93 98 9b 95 8f 8b 94 97 9e 9b 89 94 8d 90 89 89 89 85 84 8b 80 80 76 7a 81 7f 7d 78 7a 79 74 6f 6e 71 78 72 70 75 75 78 70 7e 76 79 72 71 75 69 71 70 68 68 67 69 64 66 62 65 5f 60 5f 5f 63 5f 5a 5a 5a 5c 55 56 4b 51 52 5b 67 6f 68 5e 45 36 23 10 06 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0e 0c 19 28 37 44 4f 67 6b 7e 90 9e b1 aa 93 7d 5f 64 69 6b 6d 76 7b 7a 72 7a 77 71 84 77 7d 79 7f 84 88 8f 8c 92 99 90 8f 94
 91 9e 99 9b 94 9d 9a 98 9e 96 99 a1 a0 95 a4 a5 9f a7 a8 b3 aa ab b2 b0 b3 bb b2 af b9 b4 b6 b7 b8 b5 bc bb b8 be b9 b7 bd bb c0 c7 bb c5 bf c1 b4 ae b7 b4 a5 a9 a7 9b 9d 9b 97 93 85 86 7b 63 28 08 06 05 03 06 09 0a 04 04 06 05 03 00 06 07 03 01 06 05 03 04 06 0c 0d 0c 0a 12 15 16 45 76 8b 8d 90 92 8c 8f 92 93 99 96 96 93 97 89 8a 90 8e 93 90 8b 8d 94 8b 91 88 92 88 91 84 90 87 8c 85 8e 91 8d 9b 98 97 9d 8d 92 95 90 a0 9f a8 9d 93 90 92 88 87 84 85 86 83 81 7a 7e 79 7e 7d 84 77 6e 70 6f 70 71 6b 69 72 6f 74 73 71 76 76 71 7b 7a 6b 69 64 67 67 68 65 6b 61 5e 62 5f 5d 61 5c 5f 54 5f 54 5f 58 59 5a 56 50 4f 4e 5b 55 68 73 69 5b 48 38 2b 12 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0b 11 1e 28 3b 51 57 69 71 80 93 a5 a6 aa 96 73 68 6a 6a 69 76 6b 7b 72 72 74 78 7f 7f 7e 7f 7f 76 8a 84 81 8f 8e 8c 8e 93 99 90 9d 96 94 9c 9c a0 9a 94 96 96 96 9b a6 9e a1 9d a2 a5 a5 a8 a6 ab a9 b5 b1 ae b9 b4 b2 b4 b9 b6 bc b1 b1 b0 b6 b5 bb c1 bc c2 c6 b6 ba ba af b6 b4 b5 a9 a8 a0 9e a0 a1 92 99 88 92 82 81 68 2d 10 06 05 08 05 06 05 03 00 06 0a 03 06 06 05 03 00 0c 05 0a 07 06 09 0b 11 10 16 18 17 36 75 88 86 91 8a 8c 8d 87 94 95 96 93 94 95 91 92 89 8f 8b 8c 92 89 8b 87 8f 97 94 92 9d 8e 9a 91 8d 92 8f 8f 8f 8d 9a 98 99 90 92 98 96 9c ae a5 a6 a3 92 8e 91 89 88 87 7e 7e 84 7d 7d 80 7d 79 75 76 7a 70 75 6a 6b 6a 73 73 6e 75 6e 6e 72 76 74 73 7a 66 72 67 65 6e 64 69 65 5f 66 62 66 61 66 66 5c 5b 5b 5c 5a 59 5e 5b 57 55 59 4d 53 61 63 6e 6d 61 45 30 2e 14 0f 08 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0c 29 2e 40 52 56 68 6f 85 93 a0 a7 b4 9f 81 72 69 6b 74 76 69 70 72 6f 7c 7f 7d 7d 78 7d 80 7e 84 89 7d 80 85 90 8c 93 8c 8f 91 98 9c 97 94 96 9c 98 9c 95 94 9d 99 9d 9c 9c a3 a2 a5 a3 a4 ae a3 ae ad ab b2 b1 a9 b4 b5 b2 b3 b4 b3 ab b0 b5 b4 b5 b0 b9 bf c2 ba b7 b6 b1 ad ab b4 ab aa a5 a7 9e 91 9d 8b 84 88 87 72 32 0a 06 05 03 07 07 05 03 03 06 05 03 02 09 0e 03 04 06 05 03 03 0c 05 0d 0a 0e 15 0e 20 30 6b 8c 8b 8e 8b 87 8e 91 94 92 99 91 94 8d 90 94 8d 91 87 8f 8c 95 99 9c 9f 97 9c 98 99 98 8d 8c 90 92 91 8f 89 8e 8d 91 98 a5 9c 9d 9d a3 a3 a8 9b a0 93 88 94 7a 88 82 7e 81 7c 7a 7a 74 70 78 78 74 75 76 6d 6a 6c 74 6d 69 6b 71 6a 69 77 70 6c 6d 74 6c 65 62 65 6a 5c 64 63 5e 64 5e 60 5e 60 63 5a 5f 59 52 5f 58 65 57 58 52 58 4f 55 5e 65 6f 69 5d 4a 33 27 10 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 14 17 25 3c 4d 52 61 76 83 89 94 a7 a5 97 87 6c 64 5e 6e 6c 66 72 6c 72 78 75 7e 75 78 7b 72 7d 7d 83 85 82 84 8d 8b 8c 8c
 93 90 91 94 95 95 96 98 90 97 8f 9b 95 94 96 9d 97 98 9e 9f a3 a0 a8 ad b4 ae a5 ac ad b0 ae af ae a6 a1 b4 b1 aa a8 b1 ba a4 bf b2 ad b6 ad b4 ac a6 a9 a7 9f a5 9e 9a a0 94 94 8d 87 82 74 6b 35 0f 06 05 03 01 06 05 05 00 06 05 03 00 06 06 05 00 06 05 04 02 06 05 03 10 0a 0b 0d 16 28 64 86 87 8f 8d 89 8a 8a 8d 94 8f 8b 8e 8e 94 8f 92 91 8f 8d 8f 8f 9e 98 9c 9f a2 94 9a 9a 97 8b 8d 94 93 8d 8d 90 96 a0 9f 9e 9a 9c 9b 97 9d 9c 9a 92 8a 8a 89 81 80 82 7d 78 7a 7b 74 6e 74 75 70 72 69 69 74 61 60 6a 6b 70 66 60 69 65 6d 68 6e 66 6e 62 6d 56 61 60 5d 60 65 5d 63 5a 5e 61 5f 58 53 5c 63 51 54 55 5a 59 58 51 54 55 59 57 5f 6f 69 5c 4c 38 2b 0c 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 15 19 2b 3b 4e 58 6d 70 80 8f 9c 9d a9 99 8f 6b 68 60 65 6d 6e 65 6f 73 76 79 74 73 71 78 78 7b 82 7d 7d 7c 83 85 8b 8b 91 8f 99 8d 9c a1 92 9d 95 96 90 8e 95 93 94 9c 99 92 9a 9a 9a 9d 9d a0 a7 a7 a9 b1 aa ac a7 a1 a8 a9 aa ad ac aa a6 a7 a5 b1 b0 b1 b0 ac b5 b4 af ad a9 a2 ab a8 9a a0 a1 94 91 8e 8d 7f 84 7d 75 33 07 06 05 03 06 06 06 03 03 06 05 03 00 06 05 04 00 06 05 03 00 07 05 04 10 09 0b 14 0f 29 60 7a 87 8b 8e 89 8b 93 91 98 96 94 92 95 95 95 89 86 8d 8b 94 95 91 93 94 94 90 90 94 97 99 95 9c 8f 97 8f 9c 96 94 96 a2 a3 9f 9b 8c 91 99 8e 8c 8e 87 89 88 7a 7a 76 7a 7d 78 70 74 75 71 70 74 6f 6c 6a 69 70 68 70 6b 6b 69 6d 70 6b 66 6e 6c 64 62 6f 65 59 5f 5f 61 63 5f 62 5f 57 58 5b 55 57 54 5d 57 5f 5d 5a 55 59 55 5b 59 50 51 53 5d 6d 66 59 4c 37 2b 16 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 17 13 28 3e 47 54 67 6d 81 86 98 a2 a4 9e 8a 6f 62 65 5c 65 66 63 6c 6b 70 74 77 77 76 71 79 7c 7d 83 81 7e 80 85 80 87 89 93 99 a2 9a 95 99 96 8e 8d 94 8e 91 95 9a 95 92 96 9a 9d 9d 9f 9f a4 a4 a4 a6 a7 a4 a0 a3 ab a7 ad a5 a8 a5 a7 a7 a8 aa ad ab ae ab ab ad a6 a6 ab a4 a5 9f 9c 9f 9e 9e 94 93 90 89 82 87 7f 6d 35 0b 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 0c 03 0d 15 08 0c 17 1b 5d 7d 8d 8a 93 8c 8d 97 8f 93 9d 90 94 8e 8f 8f 94 8f 91 8d 91 87 89 90 92 8c 91 8f 94 92 92 93 94 8e 94 91 9a a1 9f 9b a4 a6 9d 99 94 8d 87 89 86 88 80 82 78 84 7c 75 79 75 73 75 6b 72 72 73 6e 6a 6a 6b 6b 66 6f 6f 62 61 66 68 77 67 6d 64 64 5f 6a 67 6d 64 59 5b 55 5c 5e 59 65 5d 5f 5d 59 5f 53 58 5e 5b 5a 57 5b 56 4f 52 55 54 51 56 5e 63 60 5e 4d 3f 2f 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 15 16 2d 42 48 5b 61 79 76 8b 99 98 98 8e 7e 6f 65 65 60 69 5c 67 5f 68 67 6d 77 72 75 75 75 7d 7e 78 7d 85 89 86 86 90 90
 93 96 98 96 99 8f 90 93 90 8f 90 8d 8c 94 90 97 9d 98 93 9d 98 9a a1 a4 aa a1 a3 99 9e a2 a3 9f a2 9d 9b a2 a1 a5 99 a3 a4 a2 a1 a6 a4 a8 9e a5 a6 a0 9e 9d 96 9e 96 98 8e 87 90 89 8c 7f 7d 73 37 09 09 05 03 02 06 0a 03 00 06 05 03 02 06 05 03 00 06 05 03 01 06 05 08 06 0a 0c 0a 13 20 4a 7b 81 87 88 81 8f 94 98 98 95 98 95 92 91 93 8d 90 90 8f 8e 90 83 88 8a 92 95 93 95 97 8a 93 96 89 9b 95 9f 9d a0 a7 a7 a0 9c 95 94 87 87 7e 80 81 79 7f 76 78 74 77 75 72 70 6d 6d 72 6d 67 6f 6e 69 73 6b 69 67 65 61 66 68 61 64 63 61 5a 63 66 5f 61 5b 59 5d 64 54 5a 58 63 52 62 62 58 59 56 55 5b 57 52 50 59 59 58 51 48 54 4e 56 53 5d 66 63 63 48 3d 2f 19 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 14 1f 2a 3b 45 58 65 75 83 8b 90 97 94 92 7b 66 61 5c 66 5e 62 64 69 75 68 70 70 6e 76 73 72 80 79 7b 7c 7f 82 87 8b 89 93 9a 9b 9f 9b 99 92 93 98 8c 93 8d 8e 95 96 88 94 9a 92 a3 9a 96 98 9b 9d a4 a9 9a a7 9f a0 a4 a3 a5 a9 a6 a1 95 99 9a 9d 9c a0 a1 a3 9e 9f 9f a2 a4 9e 9d 9e 9a 96 90 88 92 8b 80 89 82 7d 7a 6b 3d 07 06 08 03 00 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 05 0f 08 11 0c 0f 1b 48 7c 7d 8a 83 83 8b 8d 8c 96 91 91 8f 8b 96 92 8d 92 94 90 96 89 8d 92 8b 93 86 8d 8c 90 93 8f 94 91 92 92 99 95 9b 98 9a 97 92 9a 92 8e 8d 83 84 7c 7d 7f 6f 6f 6f 6b 69 72 6c 71 6a 6f 6b 6a 68 6a 66 6d 63 62 65 66 62 6a 66 65 66 5e 61 63 65 69 63 5c 5d 5e 57 60 5b 60 5f 5c 56 58 56 58 61 57 5a 5b 5f 54 58 56 54 55 53 52 55 4c 56 57 55 68 71 67 55 43 30 18 13 06 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0a 20 24 40 4a 5c 67 6a 76 8b 8c 90 94 8d 79 6a 64 68 65 65 5b 6a 60 6d 61 68 70 76 6b 6f 75 72 7b 7c 7d 80 7d 81 86 85 92 92 9a 99 94 93 8c 8f 89 96 90 85 8e 8e 92 8c 96 97 9b 96 9e 9b 9e 9e 9e 97 9e a5 a5 a3 9d a1 a5 9d 9a a2 9b 9e a0 97 99 a2 99 9e 99 9e 9b a1 a2 9a 9a 91 96 9a 9b 95 91 95 92 97 88 81 84 76 6d 42 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 08 0e 08 0e 06 17 47 77 85 89 86 86 7e 8a 8e 90 99 8d 94 8c 94 95 94 89 8f 92 89 8a 89 8f 8f 86 90 91 95 8e 96 8f 94 90 92 92 9b 96 9e a7 9b 97 98 93 85 8a 83 81 7f 7c 79 72 7d 77 6d 71 71 6a 6c 72 63 67 6d 6d 6e 6c 6f 67 60 60 65 6a 63 63 63 64 59 5e 5f 62 5b 5a 67 61 67 5e 63 5d 60 60 5d 57 5a 57 59 5a 5a 58 57 52 5e 60 5b 5b 54 59 50 5c 51 55 4d 50 59 5a 6a 5e 51 44 2e 20 0f 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 12 1c 2f 36 53 56 5f 70 7a 87 8f 95 8f 81 71 65 62 62 5d 66 54 54 5e 5e 66 6b 60 6d 6c 6e 6d 71 7c 7e 7c 80 8a 7a 7c 84 8d
 8b 99 8f 91 91 91 8b 92 8e 8f 87 94 8e 85 93 93 93 96 97 9c 9e 94 a0 9a a1 98 9b 9a 9a 9e a3 9e 9d 9d 96 9e 94 99 95 95 a1 8f 93 9a 9c 9d 99 9d 9e 91 94 93 94 98 93 8e 91 82 89 84 7d 7d 7c 6c 45 0f 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 07 0d 06 05 0a 0c 15 40 73 83 7e 84 79 87 84 89 8d 8e 94 8f 87 8f 8f 8d 93 93 84 8f 91 8a 89 87 91 91 90 95 97 8e 90 93 89 96 8f 99 9c 9e a0 a0 98 9a 8a 89 85 83 78 7c 72 7a 76 6f 6e 6a 72 72 6b 6c 66 68 59 66 64 60 63 60 62 6d 5f 60 6b 5e 64 63 62 5e 62 5d 67 5d 5b 64 5f 59 60 59 5a 5c 61 5a 5c 51 58 59 53 59 56 4e 5f 56 5f 5a 56 53 53 51 55 50 4d 4e 4e 53 66 60 6e 51 40 32 1a 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 14 18 2d 3c 46 5e 5e 6f 7d 87 89 89 8c 85 64 66 5d 60 5a 5f 60 61 60 5e 67 6c 68 61 68 7a 71 76 7f 78 83 83 87 88 85 8c 8c 90 8d 8e 90 84 89 84 88 8f 8b 8b 8e 8e 94 85 94 97 8f 97 95 98 9f 95 9e 9b a0 9c a0 98 9e 9e 9a 96 99 95 9b 92 90 94 98 92 97 9d 92 90 92 8f 96 99 8f 94 94 92 8c 8a 89 8f 90 8e 87 7c 7f 72 74 4d 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0b 0f 04 0b 18 3e 70 79 80 80 84 7e 8a 87 90 8d 87 96 8c 95 94 8c 92 90 8d 8e 89 8c 90 8e 93 90 8b 92 8f 96 8b 91 95 96 8e 9d 96 9f 9d 98 8f 95 8b 8a 86 85 7d 7d 7b 6e 71 69 65 65 67 64 6a 69 66 62 65 67 64 68 61 5d 66 63 62 62 65 64 67 63 5e 57 5f 55 59 65 5b 5e 5e 59 64 5d 57 57 59 5b 54 54 50 53 5a 57 5b 4f 59 5f 5d 5a 5b 57 50 4e 4b 4e 58 50 55 5a 5a 69 64 57 41 2e 1f 10 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 07 10 1d 27 3a 4e 5d 61 72 7c 7f 94 8d 8a 79 68 5b 62 5f 63 5f 64 63 62 61 5f 5e 6c 6d 64 6d 67 72 7e 80 83 86 8a 82 85 84 8b 90 95 92 8a 86 81 89 89 85 93 90 8d 8b 8c 8c 8a 91 99 94 9e 97 9d a1 9d a5 97 9a 9a a3 98 9c 9b 95 9d 90 9a 97 95 8d 95 8f 97 8e 94 92 90 93 95 8b 97 93 88 89 8b 8a 8c 85 88 8a 89 7d 80 7a 6f 4c 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 07 03 00 06 05 03 05 06 08 0a 08 0f 2a 71 7a 85 8b 87 8b 7b 88 92 8b 86 90 88 93 95 98 8b 94 94 93 90 93 9a 93 93 9b 94 92 98 95 91 97 93 8c 9c 9a 96 9b 9f 9f 91 91 8e 87 81 7d 78 79 76 74 73 77 6d 63 6e 65 6a 67 64 60 57 62 62 63 66 60 61 65 5e 62 66 66 67 64 64 61 62 62 6a 69 5c 5f 52 64 5f 5f 60 64 52 5d 5d 58 5e 50 57 54 52 55 58 60 63 5d 64 57 57 5e 52 54 55 56 52 5e 5a 62 5c 51 43 2d 1e 11 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 14 19 25 41 47 54 69 71 75 7d 83 8f 84 6f 64 56 56 62 60 57 64 60 62 60 61 64 62 62 66 69 6b 72 71 76 79 82 8c 7f 7e 7f 87
 93 95 89 84 86 7a 7f 84 83 87 80 8c 90 8c 8d 92 8a 96 90 9b 92 99 99 97 98 93 99 9e 93 94 97 9b 92 90 8a 88 92 93 84 92 8c 91 90 8a 90 8e 8a 7f 92 87 8c 91 8a 87 86 8a 88 85 76 75 77 76 75 70 53 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 07 06 0f 14 30 62 7d 85 82 79 88 7b 8e 85 96 8f 8f 91 96 90 88 92 8d 8f 93 90 8a 90 85 92 95 96 97 97 8f 8d 94 8b 92 92 95 9b 98 95 94 91 87 89 82 85 80 75 73 73 6a 71 6c 66 65 67 65 62 5f 5d 5b 5d 57 62 61 61 5f 5f 63 61 5a 57 5f 68 64 67 5b 5e 59 5b 61 5f 5d 5d 5c 56 58 60 51 55 58 5b 59 5b 51 54 57 5c 54 5d 5d 5f 5b 59 57 57 50 59 4c 50 51 45 5a 57 64 65 54 41 32 17 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 0c 24 37 47 56 60 6d 77 86 89 88 83 66 62 5b 59 5b 55 61 5b 5e 62 5c 65 63 64 64 70 66 6d 73 73 71 7d 77 81 84 88 91 88 86 89 7c 80 7e 7e 7c 7f 86 8a 84 82 87 88 8e 92 93 8f 97 95 96 8f 95 90 97 92 96 97 97 95 94 90 93 96 90 99 92 8c 87 91 8d 90 8e 7f 87 88 85 8d 87 80 84 8d 87 87 7f 84 80 88 82 7a 75 7a 7a 69 4b 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 0a 04 06 13 24 65 7b 8a 8b 81 7d 86 84 91 92 88 8a 89 87 8d 94 8d 8a 8b 8d 95 8d 90 93 93 94 94 94 99 90 90 90 8b 8e 9b 92 94 96 95 94 8f 88 8c 82 7a 76 77 74 70 69 72 64 61 62 69 62 64 5f 5e 64 60 61 60 60 5d 5c 62 59 5c 60 66 57 58 5a 63 58 58 60 5c 59 5b 5a 5a 61 59 5e 57 57 5d 4f 55 53 54 54 53 55 52 5b 55 56 52 56 59 5a 58 52 58 4c 49 52 55 50 53 60 5e 56 43 33 19 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 1f 3a 4f 5d 67 74 77 81 87 7f 7d 63 5e 51 5e 58 63 58 60 5b 5b 61 5a 5b 64 62 61 61 68 70 73 80 7b 7a 7e 78 87 8d 83 86 86 80 7b 76 71 76 7c 77 88 81 86 90 8b 93 8a 8f 94 9c 97 95 93 92 9b 96 95 9e 97 9e 9a 8c 95 95 8d 91 92 8b 8e 8e 8b 8d 81 84 84 88 80 86 88 8b 8b 87 7d 86 8a 8c 7e 86 85 7e 81 7e 7b 73 73 49 1a 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 06 06 09 14 1f 52 7d 80 86 84 7f 86 8c 92 8b 8f 87 84 8d 90 91 93 96 8a 88 91 98 96 97 9a 99 93 99 8e 90 8a 94 94 91 8a 94 93 8e 98 89 86 84 7d 75 75 77 75 69 6b 67 6d 63 63 69 60 6a 64 64 5f 5d 57 5f 5f 63 66 5f 5d 5c 58 5a 60 5c 5d 67 63 66 56 5d 5b 59 60 67 5e 62 57 5b 54 5a 57 5b 56 54 54 4f 5a 59 59 51 5f 5f 4d 58 58 56 5e 52 53 52 52 59 55 52 5b 5b 60 59 3f 2f 1d 0a 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 24 31 46 57 61 76 79 81 87 82 71 5f 5b 4e 59 59 60 62 57 58 5f 56 62 5e 63 66 63 65 68 6e 6f 73 6e 70 74 78 7d 7d 80
 79 80 7a 75 7b 7a 7a 79 81 76 83 7f 89 8e 89 8a 96 8f 91 8e 95 95 91 98 9a 95 8f 91 9a 92 90 97 97 94 88 8e 7d 8b 8c 86 8d 7d 85 82 8a 7b 7e 81 89 89 81 8a 7f 7d 83 75 83 7e 76 73 71 80 73 6b 56 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 0b 09 03 04 13 16 4b 79 82 84 88 85 85 8d 88 8f 8e 8c 83 91 93 81 97 8e 98 94 91 93 8d 92 90 89 8d 88 8b 88 89 8d 86 8e 89 95 93 92 8b 80 80 7e 77 77 71 6f 6b 6a 6a 69 64 64 5e 5a 63 64 5d 5f 59 5a 60 5d 61 5e 60 5a 5a 64 59 5f 60 65 5b 60 60 54 53 58 5a 54 59 60 58 5a 52 59 53 56 56 55 52 51 4e 5a 54 5b 58 5b 5d 5e 52 55 5e 56 56 50 55 46 4c 58 4d 54 58 5b 5f 52 3c 2b 15 0d 07 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 1a 2b 48 50 5f 6d 78 78 85 7a 70 52 4e 55 5a 5c 65 65 5f 60 5d 5b 59 5a 60 60 64 5f 6b 66 63 6d 66 71 78 79 7d 7a 6f 74 79 75 6d 75 74 75 70 75 7b 83 78 80 82 7f 8a 8c 8e 8d 8d 93 90 9b 8d 95 93 96 93 94 93 91 99 95 8f 8f 84 8f 8b 8b 84 89 7e 85 84 77 79 7e 83 80 83 78 70 7b 78 7b 79 78 7a 72 75 68 73 75 70 56 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 1b 52 7a 85 89 8c 7d 85 89 8b 87 88 88 85 90 86 8b 86 90 89 90 8f 93 92 8e 94 99 90 94 8c 91 87 8a 88 85 8b 8b 83 89 8b 86 7e 7a 76 6e 64 70 65 6b 63 60 66 66 60 5c 61 60 5c 54 53 56 5b 5d 5c 62 5b 5e 55 5a 59 60 55 53 5a 59 55 5a 55 5d 5f 5f 60 58 5a 55 58 5a 5b 54 55 56 50 54 54 4f 58 54 58 55 5a 5c 5c 55 5c 4c 4e 4e 4e 54 4f 59 4c 52 57 56 63 47 34 25 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 10 2d 3d 55 5a 68 7b 85 85 7a 6a 5c 4e 48 51 5c 5f 5f 5d 58 59 5d 5a 5a 60 5f 5f 59 57 66 63 68 6a 69 6b 75 77 73 75 7a 78 75 77 75 79 72 7c 75 79 76 7c 83 84 81 83 8e 89 91 8a 8e 96 8f 99 93 95 95 8d 8d 99 8e 93 91 84 84 8c 8a 8d 8a 7a 85 89 86 87 7e 85 77 7f 7b 73 7a 80 75 77 7f 73 77 6f 78 75 6b 6f 69 65 51 25 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 1a 4a 70 87 88 89 7f 80 85 8e 87 8e 8d 8e 8a 89 8b 85 91 8d 8f 91 89 8e 93 90 93 8a 84 8e 86 85 8a 83 88 82 90 7d 8c 88 81 80 7a 74 71 65 69 66 6a 64 66 64 5e 5c 62 64 5f 57 5d 59 61 5f 5d 58 58 59 55 56 5c 55 60 59 5a 59 5e 55 57 5a 58 5a 54 5f 5d 54 5d 57 59 57 55 59 51 54 54 4b 5b 4e 5d 62 5e 61 5b 4d 58 5a 55 51 4e 50 47 4f 5b 59 4e 56 5e 5d 4f 3a 1e 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 0b 25 37 4b 64 6d 6f 78 82 7e 70 5a 4f 56 51 5b 66 5e 60 61 58 55 5a 5d 5e 5b 53 5e 5b 63 6b 6c 67 70 6e 6e 6c 6e 72
 73 75 7a 78 74 74 75 76 72 78 79 83 85 81 83 7d 8d 86 85 90 89 8e 87 8e 8f 93 90 9a 90 90 8f 8e 8f 8a 81 87 84 7f 7f 81 89 7f 81 88 84 75 80 7f 7c 7d 7b 82 74 7a 81 76 6e 76 75 75 6e 71 69 68 58 2f 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 17 3f 78 86 89 85 8a 8a 86 8a 8c 88 85 80 86 8a 8b 8b 8d 86 8a 8e 87 93 8e 91 90 8c 8d 87 82 87 89 7c 85 8c 7f 82 78 76 7d 6f 70 75 68 73 70 6d 6c 6a 67 68 67 5f 56 65 60 58 5d 54 60 5f 5c 52 5f 5c 58 60 55 55 55 54 55 58 5d 54 58 59 60 59 5b 5a 5e 58 54 61 52 51 50 58 59 54 57 4c 51 56 5a 67 64 5c 5d 54 5d 51 4d 54 50 58 51 52 4f 4e 4a 54 56 5e 45 26 1d 0b 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 0e 17 2e 3b 53 69 74 80 8a 80 67 52 52 49 54 52 5d 55 64 56 5b 61 5b 59 5b 56 52 5b 54 63 64 62 56 5d 69 6d 69 69 75 72 74 6f 6d 70 73 6d 6d 72 72 79 71 7f 7b 8d 84 80 80 8e 84 8d 8c 8a 93 96 97 8b 94 89 8d 8f 8b 87 87 85 86 86 87 87 80 86 81 86 80 7a 80 80 76 75 7e 7e 72 76 79 7c 78 6f 6d 6e 73 68 6d 68 65 58 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 01 06 05 03 03 07 0b 34 6e 85 85 85 88 80 88 80 90 7f 7f 80 84 8a 8a 8d 8c 88 8b 92 8a 92 90 85 8e 8b 87 85 82 81 84 89 7d 80 75 78 72 77 76 73 71 74 63 68 6a 66 66 62 64 61 5f 60 5f 5a 5b 57 54 58 5b 5c 52 50 5a 58 5c 5a 52 53 58 53 58 59 5a 50 53 55 5a 57 56 50 58 58 57 58 50 4a 4f 54 4d 4d 50 4c 57 5b 58 5b 5a 50 59 49 50 51 51 58 4f 56 49 48 4d 4e 52 54 56 49 3c 26 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 09 15 23 3e 59 64 6a 8b 89 81 6c 54 4f 4d 55 58 59 5e 5c 59 54 57 55 53 55 59 5a 54 58 5b 60 65 60 67 6a 5e 69 67 6d 78 6d 6b 6b 6b 70 70 6e 76 76 71 7b 6f 84 7e 7d 85 80 7f 88 83 80 8d 87 8d 8b 94 8e 8c 8e 8c 8b 8a 89 89 84 80 7e 81 85 89 86 80 7f 7e 7e 7e 74 7c 70 77 74 74 6d 70 6b 65 70 70 6b 6b 6e 6b 63 57 2c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 08 07 33 67 86 87 80 8b 8a 8a 8e 87 89 81 81 8a 84 86 8f 8d 8d 8d 92 8d 91 89 92 87 81 85 88 83 85 80 7f 82 7c 7f 7f 72 71 6c 6b 69 65 64 6b 65 66 69 6c 67 69 5f 66 69 61 5c 57 55 53 5b 5a 4f 5e 58 55 52 54 57 50 53 53 55 57 56 61 55 57 56 51 4e 51 65 52 55 53 5b 56 50 54 50 55 4d 4d 50 59 57 66 55 4d 56 50 55 57 58 58 53 52 55 4b 50 52 4b 4d 51 49 36 22 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0c 23 3d 4e 65 6f 79 8b 80 73 57 53 4e 53 5e 60 61 5e 4f 53 54 61 54 5e 5b 59 57 53 5f 5d 5b 5f 61 62 66 62 5f 69
 6c 5e 63 63 64 6a 63 66 72 6f 75 7b 75 72 7b 75 7c 7d 7a 88 83 81 89 7d 8c 88 85 89 87 90 93 8e 90 8b 90 8b 85 87 84 87 85 80 7e 7e 7e 75 7a 77 77 78 76 70 74 73 6c 70 6c 75 71 72 65 6c 64 61 60 36 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 08 06 2c 64 81 7e 8d 89 86 86 85 90 7e 84 73 7b 81 83 86 88 8f 8d 8c 90 8f 8c 8c 8f 8c 83 84 7e 7e 83 7a 74 6e 70 73 6f 72 6d 66 6a 71 6c 6d 61 66 64 69 61 63 61 55 61 5c 64 56 59 5c 55 5d 54 5b 5c 57 52 53 51 54 57 52 54 58 5c 55 5c 56 57 4c 4f 59 5b 5e 58 57 5b 4e 50 4c 49 4d 58 52 53 5c 5a 5b 52 4a 59 54 53 4d 56 55 50 4f 50 4f 4f 4c 4a 51 48 3e 2a 1a 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 12 1c 2a 45 5d 6f 7c 81 7f 6e 5b 55 56 56 5b 63 67 64 5f 58 55 53 4d 58 55 54 53 4f 50 5f 52 56 5d 5c 5c 5d 63 64 61 64 5f 5d 5a 5f 62 68 64 69 62 74 70 6e 6f 76 72 7a 77 7f 75 7b 84 8b 8a 85 8a 84 81 7e 89 8a 89 8e 86 84 89 80 7e 7f 81 7a 80 7e 78 82 81 7a 77 71 75 73 72 6d 71 6a 6b 6b 70 74 6c 6e 62 65 59 35 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 11 1f 5d 88 8d 88 8e 85 81 83 81 84 84 83 7d 87 7e 88 8a 89 89 8a 8e 8b 8e 99 8d 8b 81 7b 81 78 7b 78 6f 6c 75 69 72 6a 64 6c 67 6b 69 64 67 6a 66 63 58 56 63 59 5a 55 5c 59 53 63 5f 53 5d 57 56 56 55 52 4c 54 56 58 58 59 4e 4d 57 50 55 54 54 52 52 4a 56 51 58 57 52 56 50 55 5a 55 5a 5b 54 53 51 52 5a 54 4e 4b 54 52 53 4f 4e 54 4e 48 45 4a 3e 2c 1e 0a 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 01 06 05 04 07 0c 1d 24 42 51 61 80 80 7f 74 5f 58 58 5e 60 62 59 60 59 57 57 53 55 50 5d 50 54 5a 57 53 54 5f 5d 5e 64 56 62 62 60 5f 5e 5c 5b 5f 5c 62 69 64 6f 68 68 6d 75 6f 6c 73 7a 7b 78 7b 80 82 7e 7d 7f 7d 83 82 88 88 8d 8d 84 89 85 88 8a 84 88 7b 7e 7b 77 7c 7a 77 6f 6f 73 73 67 78 6e 69 71 6a 6a 67 72 69 6e 64 56 33 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 05 05 05 06 12 27 5b 84 89 8c 7d 8a 84 85 7e 7e 82 74 82 83 83 79 7f 85 8b 8b 8b 8f 8e 9b 9e 8e 84 74 82 76 76 74 72 6d 6f 70 6c 6d 65 69 6a 6f 69 5a 6f 69 65 66 5e 58 66 5b 59 5d 5d 53 55 5f 57 55 5b 52 58 5b 57 55 50 59 53 55 54 51 55 50 47 58 5b 51 52 54 59 55 54 53 51 53 52 58 4f 59 4e 57 55 5e 57 56 54 57 5b 53 4c 55 53 55 53 4d 51 41 52 50 49 4b 2d 25 1c 04 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 07 15 17 28 47 65 72 8d 85 6f 68 5f 56 56 60 61 63 5c 54 56 50 4d 5b 57 56 55 4a 4f 56 54 5d 59 5d 5b 56 5f 65 64
 63 5e 5b 5f 64 60 5c 65 65 68 65 65 6d 71 71 7c 73 73 72 78 7d 76 75 7a 80 7e 77 7b 7d 7f 84 7e 83 7e 7e 8f 82 8d 80 84 84 80 80 7e 7b 79 7a 75 7c 74 72 6f 73 70 67 6c 6d 69 71 70 60 6f 69 65 63 3e 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 01 06 0e 21 57 82 82 84 89 83 84 81 86 7e 7f 76 7b 7d 7c 84 84 80 8a 90 87 89 92 95 94 8a 83 7e 7f 6a 7f 6b 76 6d 74 6d 6f 6d 6f 6d 62 68 6c 66 62 63 62 60 60 5e 5c 5d 5e 66 58 61 5b 57 5e 57 5c 4b 51 61 55 55 4d 56 57 53 4c 55 51 56 53 4b 50 53 48 55 5c 4a 54 55 50 56 4a 53 54 5a 51 55 52 5c 5b 55 51 59 50 53 55 55 5a 54 56 51 50 50 4f 4d 44 41 2e 17 10 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0c 06 1b 23 3c 58 72 7e 7a 72 66 5e 58 5b 62 60 5a 54 5a 5c 53 4c 4e 54 57 57 53 51 56 5b 53 55 5a 4d 54 54 55 5c 5a 60 59 5b 55 54 55 62 66 59 69 64 65 6f 6d 72 76 71 7a 77 6c 7e 78 79 74 76 7b 74 73 74 78 75 81 80 85 87 81 8b 85 80 88 80 7f 84 85 7a 7a 78 75 6f 79 6f 6d 70 75 6e 73 6a 70 6a 72 67 6d 6f 65 3a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 04 06 06 15 51 7c 83 8b 80 7e 82 83 7c 80 84 78 7f 7e 80 7a 85 88 8e 87 85 88 84 8e 90 8b 89 77 7b 72 77 74 70 6e 69 6a 69 69 69 5e 68 66 65 67 63 62 64 6e 5f 5e 63 5a 5e 5d 57 55 5b 61 63 59 52 51 4e 57 55 4d 54 4e 51 4f 4e 54 50 57 52 4a 4e 52 56 53 48 54 4e 47 55 55 4e 55 52 56 52 52 56 56 4b 5f 50 56 57 51 59 53 5a 54 52 5f 4c 56 4c 44 47 3c 26 1c 14 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 00 06 0c 0b 1f 36 53 6d 75 88 78 66 5c 60 5e 65 65 56 5a 51 5d 54 4d 51 5d 55 59 57 56 5a 55 52 52 55 57 55 58 59 5d 58 5e 58 51 54 56 60 5c 55 62 54 62 64 66 74 71 73 71 75 70 6b 71 75 73 73 76 76 74 70 72 7b 82 86 83 7f 81 80 83 8c 88 86 85 82 84 83 7f 70 7b 7b 6c 74 72 72 69 69 6f 70 71 73 77 6d 75 65 6c 5a 44 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 09 14 50 7b 85 80 89 83 80 7f 7d 7d 77 76 81 84 7b 7a 79 85 84 82 8a 7f 84 85 89 88 85 7d 77 74 7f 6b 70 6a 74 68 68 65 74 6a 66 6d 5e 68 66 65 69 68 64 5e 63 62 5f 62 62 58 5e 57 5c 58 5b 5a 55 55 4f 53 56 4e 51 4f 4e 54 49 53 49 4e 4d 5b 50 4f 50 54 4a 57 59 54 54 48 4f 4d 52 54 52 56 55 57 52 5c 55 52 4d 53 54 5e 5a 5d 58 52 55 4a 4d 2f 20 1c 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 05 03 02 11 09 0b 1a 29 3d 60 75 88 79 6d 62 5d 5c 62 5b 51 56 5e 57 53 56 4d 4e 55 54 57 51 57 51 54 58 57 52 58 54 5b 58
 5d 53 55 52 5d 53 4d 5b 54 5b 62 64 62 6c 65 61 6e 6c 6f 70 72 6f 75 6a 77 75 7c 70 70 74 73 7d 76 7a 7b 80 7c 86 89 84 85 82 83 81 80 7d 7e 7a 76 72 76 6d 76 6c 72 70 6e 70 72 6b 69 6f 6f 6b 5b 43 06 05 03 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 1a 49 80 8a 81 8a 7f 75 84 89 7a 77 78 7b 7b 77 7e 7f 86 85 84 85 86 86 8a 87 80 84 7e 76 76 73 70 73 6e 68 70 6c 69 6c 6b 61 5e 69 64 6a 67 62 61 60 5e 60 62 65 66 60 58 5d 61 60 5f 63 55 57 61 5d 58 4a 4a 50 51 4d 51 4d 51 4d 52 61 4f 4b 4e 54 53 59 4a 57 50 49 55 4d 57 4c 54 4b 56 55 55 57 56 5b 54 51 53 5b 5f 56 59 50 53 51 4d 47 2e 1e 10 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0c 0c 18 21 32 4f 68 81 7b 65 6a 61 56 60 59 56 53 52 5b 4e 4d 51 58 52 50 4f 50 55 54 51 53 51 54 4c 50 4f 5b 52 52 54 4d 52 54 4e 5d 56 5a 60 60 5e 55 68 64 65 64 66 6e 6f 66 6e 70 6d 72 6b 6f 67 71 80 79 7d 7b 75 75 8a 87 8c 84 87 8b 8d 84 7d 77 7a 77 78 74 71 74 70 69 6f 6f 6c 6c 6d 66 69 6d 6e 6d 63 31 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 05 12 44 7b 84 85 88 7f 82 7c 80 79 79 78 7f 82 77 83 7c 7b 84 7f 7f 82 7c 7a 85 82 7f 6f 7e 6a 73 68 69 65 65 5e 65 69 63 65 64 65 62 5c 67 5b 5a 6a 5a 5a 64 5d 5f 60 60 64 57 5d 57 5d 60 60 58 53 59 55 51 49 4b 4a 4e 4f 52 4f 4e 4f 44 51 49 4c 54 52 4e 51 4f 55 4d 4c 50 53 54 51 52 5d 52 52 58 55 5b 54 52 51 50 59 5e 5b 57 5d 53 54 37 2f 15 16 06 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 09 11 14 21 33 56 6a 7f 6d 60 63 4f 59 55 57 55 52 54 4e 55 5a 46 50 4c 4d 56 4b 51 4f 4c 52 54 52 56 57 5a 53 59 51 4a 53 4c 4f 54 50 5c 55 57 5d 5a 61 64 65 6d 6a 6e 60 6f 66 68 72 6f 6d 6e 6a 74 70 77 75 6d 7f 81 7e 7f 8a 80 80 83 84 82 86 74 76 72 72 6b 6d 6f 68 6b 6b 73 6b 61 6b 69 69 6e 68 69 5d 32 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 15 3f 7f 84 85 86 7b 7c 7e 7e 77 78 81 83 82 81 7a 84 7b 7c 78 7b 7e 7d 7f 81 84 7b 78 78 6e 69 69 65 60 66 5c 6b 62 62 62 5d 5e 61 61 56 59 60 61 61 58 5d 5b 60 5e 55 65 54 5f 63 57 5f 57 5b 55 55 50 4d 4d 53 4b 4a 4c 51 4d 52 4a 49 48 4e 50 54 51 54 48 4c 47 49 50 4e 56 4e 51 51 55 53 57 54 54 53 55 56 54 51 57 54 51 50 4e 50 44 38 2e 0b 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 08 11 0a 13 18 1e 33 4b 63 76 6d 60 5c 56 56 4f 58 58 54 56 5d 57 49 50 50 4a 52 53 52 58 4e 51 53 54 4c 54 53 55
 50 56 56 5a 57 53 52 54 53 54 53 59 5e 57 5a 5f 67 6b 64 69 65 69 74 66 77 6c 6f 6e 67 6f 71 78 79 70 75 7b 7e 87 81 83 8a 84 82 87 80 75 73 75 74 6d 70 6a 6a 66 74 6b 6a 6b 6f 6e 6d 6a 6b 63 69 48 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 05 17 39 78 81 8b 85 84 7f 80 76 7b 7b 81 86 89 7c 85 78 81 7f 76 7d 80 7d 81 84 7a 82 77 70 72 6a 68 62 63 65 5d 5f 60 61 5f 62 61 63 5c 54 63 58 5e 63 60 5b 5b 60 5f 63 5b 5f 5e 54 5b 5e 53 5e 55 50 56 54 56 50 4f 55 4e 50 4e 4d 4d 52 47 52 54 4c 57 4f 4a 52 53 56 55 50 5c 58 50 5c 53 59 5c 54 59 55 51 59 5b 5b 62 53 55 57 4e 50 42 3b 22 15 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 0e 10 0a 16 1c 31 3f 59 64 61 5c 57 52 54 54 51 4e 50 59 54 48 4d 4b 4d 50 4d 4a 4a 4d 4c 51 50 55 4f 56 55 53 55 5a 4b 55 53 52 4e 4f 4f 4c 4c 4c 51 5d 5a 60 5c 5e 63 64 66 65 69 68 6b 6d 75 6f 63 63 6f 72 6b 70 76 75 7d 7b 85 81 86 87 82 83 7a 7a 7a 75 73 6b 69 69 67 6b 67 66 64 6d 70 6c 65 74 6c 6f 67 50 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 11 3e 72 89 8c 86 83 75 80 79 7f 84 7d 87 8e 8c 86 7b 76 73 73 7d 74 76 81 7f 7b 76 70 75 6b 6c 68 5e 63 5b 58 5f 5e 5a 5b 5b 5a 61 60 61 5a 5c 60 5f 59 59 5c 59 5e 60 56 5e 51 54 51 58 52 5d 4e 53 55 4e 4f 50 55 56 50 4e 4e 52 50 4d 52 57 50 51 55 57 52 4f 52 4f 5d 5a 56 55 4e 50 59 54 55 54 55 50 58 5d 5b 58 5c 60 59 4c 4f 45 44 3a 1c 10 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0b 05 03 10 0e 16 23 2b 4d 56 59 4f 49 4a 54 54 51 54 4c 4e 5a 49 45 4e 49 49 45 48 42 42 51 4f 45 52 4c 4f 4f 55 53 51 4f 54 56 54 43 51 49 5f 4a 4c 57 60 56 57 55 5d 5a 63 66 5f 65 64 69 69 74 5b 6a 68 70 73 68 69 70 7d 74 77 7b 81 8a 83 7e 84 7d 80 70 78 75 6a 68 6c 5f 69 65 68 6a 68 69 6d 6d 6a 6f 6d 68 54 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 33 70 86 80 89 81 82 7b 7c 7d 7e 70 85 81 81 89 83 7a 77 6d 6f 76 78 7d 75 7c 7f 75 6b 65 6a 5f 65 67 64 62 5f 64 59 69 59 5e 62 5d 60 5b 5d 5b 5b 5f 5e 4e 4f 54 4d 58 4d 5b 56 52 56 59 55 4d 4b 48 51 4b 51 54 4f 52 4f 4f 51 4a 4d 4d 4a 52 53 52 5b 4b 52 53 54 59 55 60 5f 4f 57 51 57 57 57 53 59 63 5d 60 59 5b 52 50 47 44 4a 40 2d 17 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 06 10 13 12 13 1d 26 34 36 46 4c 51 4a 4d 4f 51 50 4e 4b 56 55 4c 47 4b 43 4a 4a 44 48 49 47 48 49 4e 41 42 44 4f
 4c 53 53 55 55 56 52 5b 4d 4d 55 53 4b 50 56 5e 5b 5e 58 66 60 67 61 5b 69 67 67 6b 6a 6a 6d 70 6e 6b 66 73 6b 76 7c 77 7f 7a 80 7d 75 7b 73 75 6e 6f 6d 6e 62 6e 67 64 66 62 72 6b 6e 64 6c 6b 66 54 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 2c 70 83 8a 87 7e 81 86 88 78 77 76 81 82 80 87 83 7e 80 72 6f 72 75 78 73 6e 78 72 76 67 68 65 60 5f 67 60 5e 60 5d 5d 5b 5b 5e 59 59 58 61 57 58 5c 5e 57 56 5b 52 52 49 57 51 4a 4c 4d 57 57 52 56 53 4f 50 52 4d 4e 56 55 57 4f 4f 4f 53 4d 52 55 54 52 57 4f 55 5b 56 56 5b 53 57 4d 51 59 52 55 5d 63 5b 5c 60 58 56 54 46 49 4b 3b 2f 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 0a 0d 0a 15 16 17 22 2c 28 3e 49 49 42 49 53 4f 4a 4d 49 49 48 4e 4e 43 4a 4b 41 42 3f 49 45 4e 44 46 43 42 4a 44 48 51 4e 4f 52 4d 4e 58 4f 52 4e 53 4e 52 58 53 5b 59 55 57 59 60 61 62 65 60 61 6e 6c 69 6d 65 6d 6e 6d 70 73 6a 6e 74 7e 7a 7d 7d 71 77 72 6d 75 6c 6b 69 58 69 68 6d 60 6b 71 6b 6d 69 67 69 5e 5a 24 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0b 2d 66 83 84 83 82 7b 80 78 74 78 77 80 7e 7d 80 89 7f 83 78 77 71 72 7a 74 73 77 73 6d 66 69 67 6a 66 63 5f 60 5e 58 57 5b 5c 5e 5b 59 56 55 56 58 57 55 51 50 5a 55 53 50 56 4d 4a 50 4d 4d 58 4f 51 4b 50 52 4a 53 53 50 55 50 56 51 54 52 51 5e 57 5b 4e 4e 53 54 50 5b 59 58 4a 58 5e 54 57 58 58 56 55 5d 64 63 5b 55 52 4b 44 41 3f 25 11 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 11 13 25 25 33 35 41 4a 45 4f 47 43 49 46 44 4d 42 48 3a 3c 46 3d 4e 46 45 3d 40 40 3f 44 3e 43 3f 49 3f 4f 44 4e 46 47 4b 4d 4d 4d 51 48 4f 4a 46 5b 52 54 59 5d 52 5b 5a 5f 61 61 5a 6c 5f 60 63 68 62 62 6f 6a 74 65 6b 75 72 76 72 6f 6e 70 75 6c 74 68 6b 65 62 6b 65 66 67 67 6c 69 66 61 67 6c 68 5b 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 24 5b 7d 84 86 81 78 78 7d 6e 7f 70 78 75 73 7c 7d 81 82 7d 70 73 6b 6c 6e 6b 78 71 6f 6b 65 6c 5f 62 61 5e 5e 5e 56 58 56 57 64 5c 56 5e 60 4e 52 58 57 51 52 55 4f 50 4d 57 52 4b 4d 4a 54 4e 51 59 55 4e 50 5e 52 57 55 53 55 4a 52 52 4f 55 53 4b 57 47 4b 55 53 53 53 52 58 54 59 56 4d 5d 4c 53 5c 5a 5c 60 5b 5a 54 50 4d 45 48 35 23 0c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 06 0d 14 13 14 20 30 31 39 41 4a 42 47 4b 41 4a 44 42 49 44 4d 3b 45 41 43 47 48 3e 3b 4a 3f 3c 40 3d 4c 46 4d
 3d 44 43 48 4d 4d 47 52 56 4f 55 4e 4e 51 53 53 54 4f 4f 55 59 57 56 63 63 5f 60 5e 64 67 6a 5c 64 65 61 67 5f 64 6d 71 75 6e 6f 68 72 6e 6d 71 73 6f 6e 6b 69 74 72 64 64 68 65 64 64 6f 73 6f 63 5d 2a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 19 57 80 7b 84 77 7e 7d 7d 74 72 71 75 78 77 75 77 80 7f 85 7a 71 77 6b 6d 6d 6d 69 6a 67 6f 63 61 5e 5b 64 5f 55 5c 59 52 5b 5f 59 51 56 58 62 5b 56 54 51 4f 58 5b 53 50 49 50 50 4d 4c 54 4f 4f 53 4a 4a 56 56 4b 51 5a 4b 56 55 5a 55 57 58 5e 52 59 4f 4e 55 4e 53 55 56 59 51 50 5c 55 5b 58 5b 5a 54 56 5d 5d 52 59 50 4b 47 3d 35 1f 0e 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 03 10 20 20 21 25 3c 3e 4a 4c 44 48 43 42 44 47 43 38 3b 42 45 42 43 38 41 3f 45 3c 4b 40 48 46 46 45 40 45 46 42 45 4c 47 43 4e 4b 4c 4a 52 51 46 4f 51 50 4e 58 4c 51 58 5b 5a 5b 5d 5f 5e 5e 5b 66 62 68 60 5a 5b 61 64 6c 67 6b 69 70 6d 6a 6e 6f 6c 71 67 6a 73 6d 70 6b 67 60 60 65 6d 63 6b 6d 68 6c 5b 28 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 1f 4b 72 76 84 7b 73 74 77 73 72 73 72 7b 6c 71 72 6d 82 7c 77 70 76 6e 6c 6a 6a 6a 6a 63 64 62 64 5e 5b 63 5f 59 5d 56 5b 58 61 5a 59 50 5b 57 4f 50 56 52 48 4e 4f 4a 4b 56 56 53 4e 4e 53 4c 4c 56 4e 46 48 57 52 55 4e 52 57 47 53 50 52 55 5d 55 59 4a 4f 45 48 5b 4b 4d 4e 51 52 50 53 59 52 58 58 58 59 5a 59 60 4c 53 43 46 3f 2c 24 06 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 09 0b 0f 0f 17 1e 21 32 39 34 42 45 49 44 3e 42 47 47 3e 49 44 45 3c 47 44 3d 3d 44 48 3f 3f 47 4c 3f 40 42 3b 42 40 43 46 40 41 4c 44 52 4f 4e 4b 50 50 4a 51 51 51 53 4e 48 58 5a 57 63 61 59 5b 5e 62 64 69 66 54 59 60 62 57 60 63 61 6a 6b 64 69 68 60 6c 70 6b 69 68 6e 6d 68 6a 5c 62 5a 60 62 66 66 67 64 60 32 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 18 46 74 78 7a 7f 76 7a 74 70 67 6d 6f 70 70 71 6e 77 70 79 7a 74 70 6d 69 6a 63 6c 61 65 6b 66 67 61 62 5f 50 5e 5b 50 54 57 54 4e 54 51 53 52 50 52 51 51 54 52 46 52 53 54 4a 52 57 49 5a 57 53 54 58 53 50 50 4b 55 50 52 50 4a 50 53 54 50 50 4e 4c 53 4b 52 4c 4e 50 51 54 50 4e 56 55 62 5c 54 5d 5e 5b 56 5a 55 55 4c 44 3a 38 20 0d 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 09 15 11 12 20 2b 33 39 49 45 45 49 3d 3e 44 40 46 42 43 47 3f 3f 36 3c 3b 3f 44 46 41 43 46 4a 41 47 47
 3f 44 4c 39 44 41 47 4a 4d 46 51 54 55 4f 4a 4d 4d 4e 4f 53 4a 4f 55 4e 59 55 57 55 5c 5c 69 4e 33 45 63 61 5c 59 57 5d 60 66 62 5d 59 5e 5e 64 6e 67 6f 65 62 65 68 61 67 5d 5d 5d 64 6b 60 61 6b 5e 37 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 19 51 76 76 7e 76 74 7a 70 75 72 70 6d 73 6d 6d 6f 6d 75 6e 74 77 72 62 6f 70 63 63 67 64 64 5b 60 65 5b 5a 5b 52 52 5a 52 60 55 4e 48 4a 54 58 4e 4c 57 4d 50 55 54 55 56 55 54 52 4f 52 5a 4e 52 56 55 56 4e 50 4b 4b 4a 56 4f 52 51 54 5b 51 47 50 4b 4d 4f 51 4e 52 4e 52 56 58 52 59 59 5a 54 58 55 59 66 5e 5c 5b 50 51 3c 3a 37 20 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 07 10 11 14 1c 1c 25 39 37 41 46 44 48 48 41 47 3e 41 46 44 43 45 3c 43 40 43 43 42 44 45 40 42 45 41 45 40 40 42 43 45 45 46 47 49 46 49 52 4a 56 4f 45 4e 51 45 4f 4b 51 53 4e 49 59 50 52 5d 55 5e 5b 5a 5f 60 61 59 54 5a 5a 5a 61 5b 59 5f 5a 5c 5e 59 5b 5f 60 68 6c 6d 6c 72 66 64 62 5f 57 61 63 64 62 5e 3a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 05 0e 43 6a 71 76 76 74 73 75 6f 71 69 71 72 5f 6d 6d 6a 71 6d 75 72 68 67 61 61 5b 5e 62 66 60 61 63 5e 57 56 5d 62 5a 50 56 5b 56 55 55 59 5a 53 53 55 4b 48 56 56 52 4c 52 4b 5e 50 50 57 5f 4c 55 56 53 56 4f 56 51 48 4c 49 5b 49 54 43 55 4e 50 57 52 4e 52 55 4a 50 50 55 4e 4e 5d 54 54 5c 5b 5d 54 5d 62 5d 66 60 54 54 45 3b 2f 18 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 03 0c 10 17 21 24 2f 32 43 44 45 4e 4d 42 4a 45 39 43 41 43 43 45 43 41 3b 43 3e 43 35 44 44 40 47 3e 44 3f 3e 41 3d 42 4d 40 45 48 44 44 42 4d 54 48 4b 4f 4e 4e 46 4e 51 4a 50 54 57 51 59 55 53 63 5c 55 51 55 5b 4c 55 58 4f 5e 5e 5b 5c 54 5b 58 5d 62 5e 5d 5d 65 65 63 6e 62 61 5e 56 5d 64 56 63 62 5b 3e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 10 3b 69 72 7e 7e 6e 79 6f 72 77 69 6e 66 69 63 6b 69 71 65 6c 65 64 64 64 63 5f 5c 63 55 60 5e 5d 5d 59 4f 59 55 58 57 52 5a 50 53 50 51 4d 53 57 4a 51 44 4f 55 54 4f 51 55 58 51 50 51 58 4a 52 4c 4f 4a 56 48 53 44 4f 52 4d 51 52 4e 50 4d 52 53 54 4b 51 50 50 50 47 51 52 4e 57 53 5c 5c 50 50 5a 54 5f 67 66 61 48 47 3b 3a 27 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 16 1d 2f 21 28 2e 41 40 46 4b 45 49 42 40 3d 44 3d 45 3d 41 3a 35 3f 41 47 40 46 41 3f 40 3a 47 44
 3c 40 4d 3e 48 41 44 43 42 47 44 45 42 50 4f 50 48 48 4a 53 43 49 43 49 50 55 4c 4a 54 4e 57 56 58 51 54 5a 51 4f 50 54 50 57 5f 5b 56 55 4c 54 5b 5f 5d 61 5d 65 5f 67 69 61 65 65 5f 5c 61 58 59 53 30 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 10 38 6f 72 77 75 74 73 77 70 6c 63 69 66 69 63 67 66 64 6a 69 65 60 62 62 62 5b 59 59 53 57 59 57 52 58 57 5c 59 58 55 59 56 52 4c 4f 53 4f 48 53 53 51 4c 50 4b 4a 50 58 51 53 5d 59 5b 50 52 55 51 51 4a 48 51 53 4e 4f 55 58 4e 58 51 52 55 57 55 57 58 50 54 4a 53 50 54 54 53 55 57 5e 57 54 55 50 58 68 65 65 55 50 49 46 31 1f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0d 15 0e 13 22 27 2f 39 42 43 43 4a 46 49 41 44 49 3e 3b 44 3f 3e 3d 38 45 3f 45 3b 43 41 40 45 3c 44 45 45 3e 48 42 42 40 44 4b 48 43 46 4c 48 4a 48 4d 49 50 47 4b 4b 49 4a 4e 4d 42 50 54 51 53 56 53 57 54 5f 58 50 5a 54 5c 60 51 58 54 52 52 5c 4e 4b 4c 5a 5e 63 65 66 63 64 61 62 65 53 58 5b 5a 59 59 36 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0a 0d 2d 6b 7b 7e 73 76 77 70 62 68 65 68 5d 6b 61 66 68 77 64 5f 62 63 56 5b 59 59 5b 5f 5c 60 51 59 5d 56 5a 56 54 56 57 58 52 54 52 48 52 4e 4d 56 4e 4b 4d 51 47 50 54 50 5d 53 50 56 53 53 48 4e 50 4f 4b 4f 53 4d 54 55 5e 62 5c 5f 4e 57 54 59 4f 4f 54 5a 59 56 56 52 52 50 52 57 58 5a 59 4e 4e 55 5c 65 6a 62 65 58 47 44 32 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 06 10 1e 1b 27 3b 3b 42 45 47 43 3b 45 3b 44 4a 43 48 42 47 3a 42 3b 41 3d 41 3f 45 44 41 44 3e 4a 45 3c 3f 43 41 46 46 48 3e 48 4b 46 47 48 44 44 4d 45 53 4e 49 4d 4c 48 4a 50 54 5a 48 45 4c 4d 56 55 54 54 51 50 52 51 5e 4f 49 4f 50 58 55 55 50 55 58 54 52 54 57 55 5b 5f 65 6c 60 60 54 59 58 55 34 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 32 68 71 6e 76 70 72 6c 61 65 64 6d 60 60 61 5f 64 65 60 5e 56 62 56 57 5b 5c 59 5b 56 54 4c 57 4c 5a 5f 58 5e 5a 4e 5c 53 4d 54 51 54 54 52 4f 4c 51 51 4d 55 51 49 4e 52 57 49 4b 48 53 4c 4b 4d 4a 49 4e 4a 50 4f 51 56 69 62 5f 58 4f 5b 56 50 59 4e 56 53 55 57 55 50 5d 53 52 50 4e 53 53 4d 4c 50 66 6a 65 5b 4b 49 3e 20 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 13 13 19 29 33 3d 43 46 45 41 48 4e 43 4b 42 42 44 42 40 42 40 36 43 3c 4a 3c 40 42 41 40 3d 3c
 3e 40 47 39 44 42 40 43 47 45 45 46 3f 45 44 46 55 4a 43 50 49 4a 51 48 55 47 46 48 4b 4a 4b 4b 56 4c 51 56 58 4e 52 55 53 4a 55 49 49 54 4a 54 4f 4b 53 57 5b 55 58 5b 62 57 5a 60 62 5f 54 59 56 57 44 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 2a 62 68 70 6d 66 65 69 66 6b 5f 6c 69 67 5f 65 69 63 68 5d 5d 59 55 60 53 57 56 54 55 55 53 54 57 4e 59 52 4d 53 52 59 5d 56 47 4f 5b 4c 50 4e 42 52 4c 45 52 45 51 4f 50 53 47 54 4f 4f 4e 50 54 4b 49 4a 48 4b 52 5a 4d 60 60 5c 55 4b 4a 4f 5b 56 56 50 57 50 52 54 58 51 4e 4d 4f 56 51 47 56 5c 60 64 66 57 55 44 43 2f 1e 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 0e 12 20 23 21 2c 44 37 40 46 4b 3e 44 49 50 41 47 44 4e 3a 3a 42 3a 43 42 4a 47 46 44 41 41 40 3b 44 46 41 46 43 44 44 45 40 42 47 41 42 4b 44 47 45 43 4c 50 47 51 55 4d 4e 49 4c 4a 4e 48 4a 48 4e 4c 4d 51 50 50 4f 52 52 4b 50 54 4e 4f 4d 56 4e 54 4e 54 4f 5e 55 54 53 5d 5c 62 62 61 5b 5b 50 4c 3f 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 21 5d 68 6f 76 6a 72 6f 66 68 60 60 60 62 68 6b 6c 5e 5e 60 5a 5b 51 5f 5c 63 50 4f 58 54 4e 55 56 5b 55 4f 58 57 55 59 54 5a 4c 59 4c 55 56 4f 50 4a 55 4e 4b 4e 53 4d 54 4c 4a 52 44 53 4d 4a 59 4c 40 47 49 59 5a 5a 55 54 52 59 51 50 52 4f 51 57 52 52 5d 57 50 50 54 58 56 50 53 56 5b 4f 5e 61 64 64 65 58 53 4a 3c 28 15 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 0a 16 13 1f 26 2c 3d 3f 3f 48 40 41 49 4a 49 44 3f 4a 46 42 43 3c 46 43 45 45 40 47 43 41 41 4a 3d 3b 4d 42 45 46 45 42 43 49 45 43 4b 4b 4a 43 49 43 40 45 45 41 4b 4a 4c 49 48 50 4a 48 4b 45 4a 52 51 54 54 59 4e 4b 4b 4c 49 55 49 4d 48 49 4a 4a 50 51 52 4e 54 4c 55 52 53 56 5b 5e 5e 5c 58 55 51 43 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 26 52 68 71 71 6b 6a 65 65 6c 67 65 65 63 6b 62 67 64 5c 60 5b 5e 52 5c 57 5b 55 4d 58 53 4f 4f 4f 58 4c 5a 54 5c 56 5a 58 53 53 50 45 4d 4e 50 50 4e 46 44 53 4e 50 51 4e 49 4c 4e 4d 4c 4b 43 41 4d 4a 59 49 53 53 52 4a 56 4f 49 48 4b 5b 4f 54 5b 52 4e 50 49 4c 4b 4d 54 55 54 5c 66 5d 5a 64 63 69 68 61 58 4c 48 39 1c 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0a 15 18 1f 28 34 44 3e 45 46 3b 44 43 48 45 46 3d 4a 3e 41 3f 49 46 41 46 41 48 46 45 43 3c 44
 4c 46 41 43 3f 4a 43 44 41 3f 47 4c 3d 40 48 4e 42 49 49 4d 42 4d 4b 49 4c 47 48 4c 4a 48 47 4b 48 4e 4c 4e 4a 4b 4f 4f 4b 4b 4f 4a 45 46 47 4e 4c 46 4d 4d 4a 4f 58 4e 52 52 57 5c 59 61 50 55 4c 50 47 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 25 47 63 62 6e 6e 64 67 65 64 65 63 64 64 61 6f 62 6f 55 5c 59 58 57 53 53 50 4f 57 52 4e 53 54 4d 4b 4c 4d 59 50 50 51 52 4b 52 4a 4c 51 4c 4b 49 49 4b 47 4d 4d 4c 48 43 45 43 50 4a 4c 53 4d 4d 50 47 48 45 4c 4f 52 4e 4e 4f 4c 4a 55 54 50 55 4b 4f 53 4e 4f 51 56 57 57 5d 61 62 56 5f 5f 66 71 70 67 59 4c 50 3f 34 17 06 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 0f 1c 1b 28 34 3f 43 47 44 40 3f 48 46 45 46 44 46 40 44 49 4a 47 45 40 3e 44 44 42 41 45 4c 42 3f 42 3e 3d 45 40 43 45 4c 47 3e 3c 49 4b 4b 4a 41 46 51 47 43 4f 46 47 4d 4a 4f 47 4a 46 52 4d 4d 47 46 4b 4d 4a 4f 4f 49 4e 48 46 4e 3f 4c 4c 45 47 4e 4f 52 52 4b 47 52 4b 57 55 5b 5b 54 52 53 42 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 1f 4d 69 61 6c 66 61 63 65 69 5f 5f 65 62 64 69 67 64 5b 5f 55 59 57 56 5c 4d 52 57 55 5a 52 61 4b 4e 51 54 59 57 50 4e 52 48 4a 4f 51 52 50 54 45 50 49 4d 53 4f 4d 51 4f 53 4b 49 4a 54 51 44 4a 4b 49 52 4b 51 52 52 4c 58 4c 4b 53 4b 47 54 52 58 4d 56 56 50 56 5a 51 63 5e 6b 66 62 63 5f 62 6c 67 68 57 4e 50 35 2a 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 0a 13 25 29 37 37 38 48 41 3c 42 38 44 3d 44 3d 3c 48 4a 49 46 4a 48 3e 44 43 41 42 3d 3e 48 4b 4d 3d 42 45 44 42 42 42 49 41 49 49 4a 4a 49 4b 48 47 4d 42 4c 4d 45 4a 48 46 4e 4b 53 51 4c 49 4b 4b 44 46 46 4a 4f 4d 45 4b 4f 49 52 41 4a 49 45 45 49 3f 50 49 51 48 50 51 50 58 52 4d 48 4a 45 41 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 16 51 61 69 66 61 65 61 60 62 5e 5e 67 67 60 61 5c 66 5e 5f 60 58 56 53 57 5b 51 52 57 53 51 5a 52 54 4e 57 50 57 49 53 52 48 4b 49 48 50 4d 51 55 4d 4d 4b 51 50 44 4b 4c 4b 4d 4c 4a 45 4d 4c 4d 4c 49 58 53 4b 52 4f 44 50 4c 50 4c 56 51 4d 55 54 4c 52 4b 4e 58 55 60 5c 5d 64 5f 55 5a 63 72 74 6d 60 50 55 43 2c 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 03 19 1d 21 29 3b 47 41 3e 44 45 41 3e 44 41 40 42 42 4b 43 45 42 44 3f 3e 3f 45 45 41 43 40
 3a 45 3a 40 3d 40 41 45 46 4e 46 44 48 47 47 44 42 43 4f 4d 46 4a 4c 44 42 46 3e 46 41 4a 44 47 47 45 45 47 45 4e 4a 50 48 46 4b 4b 45 4a 45 48 47 41 47 43 49 47 43 46 49 4a 52 4b 50 56 56 47 4c 40 47 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1a 54 5f 65 6d 65 68 5d 55 61 54 5f 5c 64 61 5f 64 65 6a 64 5d 60 5e 59 55 53 4e 52 51 4e 53 54 47 58 51 50 4c 51 4e 4f 4e 4e 47 48 51 49 4d 4c 51 4f 4b 4a 42 58 47 44 4a 4d 47 4a 49 4e 53 50 4e 47 4c 47 50 4e 4a 4c 46 49 42 4a 4d 4d 4d 49 4c 54 4e 4f 4a 4a 4c 58 50 5d 61 58 5d 54 5c 60 6d 6b 54 5a 55 41 37 20 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0e 12 14 21 2e 37 41 43 43 42 3b 44 3d 44 39 3d 43 45 47 52 44 44 46 44 41 49 48 3c 3e 3f 38 41 44 3b 3e 3c 40 45 3e 47 3e 43 42 42 47 48 43 46 45 4d 48 4b 47 4a 45 49 48 4d 49 47 4a 4d 41 4b 4c 4b 4d 3f 49 4c 4b 4d 4b 50 4d 44 4a 50 48 52 44 4a 4b 4a 47 43 3f 46 54 50 51 53 4f 4b 4c 44 3f 43 1a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 01 17 44 63 62 6b 66 63 63 64 5e 58 5b 6b 60 62 64 66 64 68 60 5f 65 58 58 58 54 51 53 49 4f 4d 4d 55 48 52 4e 59 54 46 4d 48 52 44 44 4d 49 50 4b 54 53 56 51 4a 4a 4b 4a 47 49 49 54 4d 52 4d 47 55 4e 4b 51 4b 47 50 52 4c 4e 46 4a 52 4f 4d 53 4d 57 4e 4c 4b 51 51 5f 53 65 58 4f 4e 50 65 68 72 67 51 4e 4e 40 37 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 12 14 19 30 37 39 42 43 3f 3a 42 41 3e 4d 43 47 46 3f 40 45 41 49 3f 3e 4c 41 48 49 3d 40 3e 47 3b 47 3f 40 41 44 47 4e 3c 44 43 46 49 4d 4a 47 4a 43 42 4d 45 47 4c 4a 51 48 46 41 46 4f 45 49 50 44 4a 46 44 45 48 52 48 50 45 47 4b 45 48 4f 47 48 49 50 49 46 46 3f 4e 46 48 4f 4a 4e 49 47 3d 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 10 42 5f 67 69 66 66 67 64 5a 57 5f 5a 60 62 64 62 5c 56 67 5e 63 5d 5f 5e 5b 53 55 4e 52 4c 55 51 4e 52 4f 51 4a 50 52 48 4e 4d 4e 56 4b 49 50 4e 4e 4b 48 4c 4c 4b 46 44 4b 44 4a 51 4f 4b 4a 53 51 52 57 4e 48 48 59 51 4e 4b 4c 48 4a 4b 4d 49 4e 56 54 50 55 5c 5f 5b 5b 4c 57 52 58 5f 65 5b 5d 4b 49 42 35 2a 08 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 08 13 14 26 2a 36 44 46 44 48 48 4e 44 3a 3a 3a 44 3a 41 3a 3e 44 3d 43 3b 41 3a 38 3e 40
 47 3d 46 40 44 45 3d 42 3e 39 45 49 43 42 42 44 53 41 4f 47 49 41 43 4c 48 4c 4e 45 42 43 43 43 47 40 44 46 42 43 45 44 47 4f 50 48 49 44 44 45 41 40 46 44 44 4e 43 43 40 43 3d 51 4b 48 3f 43 45 46 3e 20 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 11 41 61 64 6b 64 62 61 61 60 61 60 5a 60 60 5f 56 62 62 5a 63 5f 61 5e 52 51 4d 56 55 4c 53 53 4d 4a 4d 4f 4d 52 44 40 4c 4c 4b 46 4f 51 52 44 50 4b 45 4d 4c 46 47 4f 42 47 49 4b 45 54 4c 59 55 50 54 52 49 49 3e 4a 4c 46 48 4d 53 51 4c 50 43 54 54 4d 59 59 5c 5d 65 5e 52 4e 4c 57 60 5f 53 48 44 46 36 2a 1b 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 11 14 11 1d 2a 2f 42 41 42 44 44 3f 42 3b 42 4b 42 42 3a 42 44 45 3e 41 48 43 49 45 40 3d 42 3c 45 44 3c 40 41 3e 3c 48 42 3e 46 48 46 46 48 4a 4d 47 40 4e 4a 4b 4d 47 4e 51 43 47 4f 44 49 46 48 47 47 43 50 4e 43 46 4a 44 4c 4d 49 4f 44 4b 4b 45 4a 4f 43 48 4b 4a 47 4d 47 4a 4c 44 49 44 3b 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 3b 64 62 65 64 60 60 5b 54 52 5f 5c 58 5c 5a 5d 60 63 65 5b 64 62 5a 58 55 54 5a 52 54 52 56 51 50 51 56 52 4b 42 4e 4a 47 4e 49 57 52 51 53 45 4b 4e 46 4b 4f 4c 4b 4b 46 4c 52 51 5a 52 4e 62 5e 55 4e 46 47 58 4c 4a 47 4a 4e 50 52 4b 4f 51 54 52 50 54 62 61 64 68 56 52 4f 4d 59 59 4d 49 51 3d 3d 3b 1e 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 0a 11 11 26 26 32 44 3f 3e 47 44 41 40 38 3e 41 39 39 39 3c 3f 3c 45 47 3f 42 41 43 41 41 43 43 3e 46 3d 44 3d 43 3b 46 45 41 44 4a 41 4f 44 42 46 53 40 41 53 49 4d 57 45 55 4b 47 40 47 4f 43 4f 48 41 44 43 46 4c 47 4b 47 44 49 47 50 45 49 4d 40 4c 4c 46 44 49 47 4a 53 44 52 4b 44 43 40 39 18 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3a 61 6b 68 72 61 63 5a 58 55 59 61 5a 5c 5a 5b 5b 5a 5e 5f 64 5e 5a 55 5a 50 5a 54 56 53 52 55 51 5a 56 52 54 4a 4a 52 4d 48 44 4e 4b 4a 4c 4b 45 55 50 4f 51 49 45 4f 4e 3f 5a 51 54 5a 53 5c 5e 51 4d 4d 4f 50 4d 4d 47 50 4b 4d 4a 4b 50 55 53 57 58 61 5e 6d 6d 64 57 4e 49 4c 50 4f 4f 4e 46 3e 31 2a 18 10 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 07 0d 11 14 20 2e 36 3c 41 44 38 3a 36 41 48 38 44 3d 44 3d 38 42 3d 42 3c 3b 3b 42 44 40
 47 3b 3d 3c 45 43 40 3c 40 41 43 43 43 48 4a 48 47 47 45 47 3d 51 47 48 47 4d 51 4c 4b 49 4f 48 3e 46 44 44 4d 44 44 48 45 49 46 4c 48 45 4d 4e 4c 43 47 48 45 46 46 48 47 45 46 49 49 4c 44 44 42 3d 39 25 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 2d 58 62 6f 68 63 62 5b 5d 56 58 65 54 57 5f 55 59 61 5b 63 5e 5b 5e 5c 5c 4a 53 59 5a 4d 58 52 4e 52 4c 4d 4d 48 49 4b 4e 4f 4a 4d 54 4b 54 52 51 4c 54 57 54 55 4c 4d 52 4d 4f 56 55 55 50 5a 50 4b 52 50 4c 4e 4d 56 4d 4b 4d 51 46 4f 51 4e 5b 54 4d 59 6b 68 6b 69 5c 44 4f 4c 50 4f 40 47 45 36 26 0e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 05 00 0b 07 10 15 1e 2e 38 46 48 43 42 38 39 3f 40 46 3d 40 37 3c 3b 40 41 46 48 47 45 42 3a 40 45 44 41 36 38 3d 3e 41 3f 3e 42 3a 44 40 47 48 44 45 3d 4e 41 50 46 43 43 46 42 4b 47 4a 40 48 46 40 48 43 47 47 48 48 47 3a 4e 40 4c 51 4c 4a 4a 48 42 45 47 3e 44 44 4d 4c 49 48 46 45 45 3f 3f 3c 48 31 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 2c 58 6a 6b 69 67 68 5c 5c 4c 54 55 56 5a 56 56 63 58 59 55 58 5c 5c 53 59 57 5c 53 58 51 52 53 56 53 53 4f 54 4b 49 55 4f 51 4a 51 4b 4a 4f 4e 53 4d 4d 56 53 5c 53 51 54 4e 4b 4d 4c 4b 48 50 4b 4a 50 4e 4e 5c 58 53 4f 52 50 55 49 4b 50 48 54 51 5e 62 77 71 63 55 4d 4b 49 4d 4b 4d 45 44 38 2c 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0b 09 12 16 1e 28 36 39 36 37 3f 3e 42 43 3e 3c 3f 3c 3b 3c 3e 3e 42 48 4c 45 43 45 4b 45 41 3e 47 44 3c 3a 3d 3e 40 40 3e 42 48 3e 41 45 4d 43 47 44 47 46 48 45 45 4b 45 4e 49 49 49 48 4d 42 43 48 48 41 42 44 48 4a 46 44 4d 46 42 4b 4a 4e 44 47 48 47 3e 44 4e 4a 4a 4b 45 4d 44 3f 42 44 3c 28 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 28 55 66 66 69 62 65 55 5f 4f 53 4e 50 55 5b 53 59 53 53 5c 5d 64 57 61 5f 55 54 53 5e 5b 5a 55 50 50 50 53 54 4c 4b 55 50 47 4f 4a 52 54 55 58 53 4e 59 54 65 5d 5a 4e 4b 47 4c 50 4c 4f 51 45 49 48 50 4f 56 4b 52 4f 53 50 57 50 54 4e 4e 4a 51 58 5f 67 6d 69 5e 56 50 4f 4e 4c 4b 47 47 3b 35 27 14 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 18 1c 2c 3a 3c 36 3b 42 41 40 45 34 3b 41 38 3d 3a 39 41 4e 4b 42 4e 45 43 47
 47 3e 43 45 3a 3e 42 3d 44 44 44 42 43 3f 3e 47 4c 46 42 4a 48 4a 40 40 52 48 4b 49 44 4e 4a 47 48 49 41 44 3f 45 40 44 4a 3a 3b 3f 40 43 43 49 41 4d 49 44 4e 40 49 52 4a 4c 44 48 4e 4d 47 43 40 47 42 32 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 26 50 5d 6e 5c 5d 5b 58 56 5a 57 5d 57 51 59 55 59 50 56 5a 5c 5d 59 60 57 5a 60 57 59 56 5c 59 51 56 50 50 50 49 47 44 49 51 52 4b 55 57 54 57 53 58 5a 5e 64 57 5c 4c 44 42 4a 41 49 44 41 46 40 46 47 4d 4a 4c 4c 49 45 47 45 51 48 4a 4f 50 52 5a 59 6e 65 53 50 51 4f 49 49 4b 4d 48 41 3c 32 13 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 10 11 28 30 39 36 3a 40 38 3e 42 39 3d 41 3a 37 36 39 3f 45 43 3d 4c 3c 3c 49 3a 44 41 3b 3c 40 36 40 42 3b 42 3e 47 38 46 45 49 40 46 4b 44 44 46 49 45 48 47 3d 48 46 49 49 48 47 44 44 44 42 42 40 41 43 3c 48 42 43 4f 43 46 40 42 40 45 47 47 46 45 4a 45 4b 4c 47 47 4a 42 48 3a 3e 29 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 22 4e 5d 64 5f 5b 5b 53 51 52 54 58 56 51 51 58 53 5a 59 65 5b 58 5a 55 59 5e 5f 55 54 55 56 53 51 51 59 50 48 4d 48 54 4c 4c 47 51 5c 5e 5f 64 5f 58 4f 59 54 4d 54 4d 49 48 47 44 4f 43 46 41 44 45 4b 47 46 4b 4e 47 4c 3d 4d 40 44 41 52 54 55 59 67 59 5a 58 50 4b 45 4f 4f 4f 48 45 42 33 27 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 06 09 12 16 1e 28 39 3b 40 3d 42 40 3e 44 3c 40 3b 3c 38 41 3e 3b 43 41 45 44 44 3f 44 41 47 43 43 40 41 41 42 3e 43 46 47 3b 4c 42 4b 45 40 4c 47 3f 48 45 44 4d 44 4a 52 3f 4a 4d 47 4c 4d 46 40 40 39 48 43 40 41 44 3e 39 4b 48 43 4d 4b 47 4c 3c 47 4b 3f 43 4e 50 46 47 51 4e 47 47 49 44 36 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 1e 45 5b 69 60 60 61 5d 5a 4c 59 57 52 57 50 61 5e 5c 5a 53 54 5e 55 5d 5f 55 55 4f 54 55 59 5b 53 52 50 51 4e 4e 4a 4a 46 49 4e 5d 61 6d 60 5b 59 52 52 56 50 4a 4d 4a 3e 48 43 46 46 43 44 45 48 46 4c 49 45 48 50 4c 4d 44 4b 49 45 4a 49 4b 53 5a 5f 5a 5d 54 4e 54 47 47 47 52 41 45 36 26 1d 13 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 18 24 2d 3e 3d 38 43 3d 3d 43 44 42 3b 39 37 3a 37 49 3a 38 3f 3a 33 39 47
 3e 46 37 3d 3b 41 38 44 43 3e 44 43 46 49 47 3e 3f 46 3e 41 47 45 48 44 45 43 40 4a 4a 4b 4b 4a 40 4b 48 45 3d 43 44 3f 40 38 42 3b 3f 43 41 40 45 43 44 4a 47 49 46 41 46 41 4a 42 40 4c 4c 4a 47 42 3a 35 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 43 59 5a 65 57 56 54 5d 52 5a 55 55 5c 55 57 4f 59 58 55 5b 5b 5f 55 53 52 58 55 57 5f 49 53 53 5a 50 4e 53 45 4f 49 44 4a 57 57 66 63 60 5d 5e 4e 4b 4b 4e 47 49 41 47 42 3c 46 43 4c 48 4b 40 46 4d 49 44 4e 44 47 45 4e 49 43 52 45 4a 4b 56 5b 5d 56 4b 51 4b 51 45 46 48 45 3f 42 3c 22 1f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 1c 1d 2c 3c 35 37 42 45 4d 42 44 3f 3c 39 3e 34 3b 44 3b 38 3c 36 41 3a 35 40 42 43 43 3d 46 3c 42 45 43 40 41 44 48 3f 3a 3a 3b 3a 45 44 43 48 38 43 45 46 46 47 47 43 4a 48 46 4c 46 3f 42 47 41 41 46 4a 41 3e 3c 41 44 3c 41 42 49 49 4b 47 41 46 41 44 48 4b 42 49 44 45 43 3e 27 0e 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1a 49 52 5a 57 58 5e 55 56 54 5d 5b 56 4e 56 5d 56 5b 56 55 5e 53 5f 54 59 53 52 5a 57 54 59 48 4f 4f 4a 44 50 4e 4c 48 49 51 51 58 58 5d 5e 52 54 49 45 47 44 46 44 48 49 42 42 3e 47 49 4b 4b 47 43 41 4d 45 48 4f 46 45 45 49 53 43 4e 50 4a 55 52 54 55 4b 53 53 3f 46 4a 40 46 3d 41 20 1f 10 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0b 0d 21 28 32 41 3c 3e 42 49 42 49 43 3d 30 39 40 38 3c 42 3c 40 37 38 3d 3a 45 42 3e 3f 3e 45 45 45 40 45 40 45 43 4c 43 3d 44 39 45 42 3d 42 42 41 47 50 3e 49 4b 44 4a 46 46 45 44 4b 3f 3d 3f 42 42 3f 39 38 47 3d 44 46 49 41 42 42 47 49 47 3e 42 3c 4f 49 49 44 42 45 3f 42 3e 33 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 1c 31 5b 62 52 57 54 53 53 52 56 55 4d 52 56 53 59 58 5b 63 58 5b 5a 51 57 54 51 5b 52 58 54 4e 52 56 54 59 56 51 46 51 52 51 4e 54 54 5a 56 4d 4b 4a 44 4d 44 46 43 48 44 46 41 42 47 4b 44 4a 46 48 4d 4a 48 4f 50 4e 43 46 4a 3f 45 47 45 4e 4d 55 4e 4e 47 46 44 47 49 44 4b 4c 3d 34 29 14 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 0d 16 21 24 34 36 37 45 42 50 4e 44 3b 41 3a 3a 3f 41 40 3e 3d 37 3d 3f 36 45
 3f 46 37 38 37 47 3f 47 43 4a 39 43 3d 47 48 3d 43 42 3f 4a 45 3b 41 44 46 3e 46 47 41 4a 46 50 56 4e 53 4d 40 4f 44 44 43 42 3a 44 49 43 36 39 41 3e 42 43 3f 42 41 38 46 39 3d 41 43 4c 47 41 39 40 3e 36 14 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 35 55 55 5c 59 50 53 58 50 59 56 59 59 52 58 5c 58 5c 57 58 5a 5c 57 62 52 5b 4e 4d 48 55 48 46 4d 4d 52 49 4d 4d 53 53 51 52 53 59 4a 4b 4d 32 4e 49 3f 49 40 41 42 4c 46 48 46 47 44 46 4b 49 40 47 44 46 4f 4e 43 48 4c 47 4b 46 46 50 4f 4f 53 4d 4a 47 49 50 4c 45 42 45 40 42 2d 1f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 0d 1d 19 27 32 36 3e 48 3d 44 48 3d 3c 38 38 37 39 31 3c 3a 3e 3a 34 36 38 41 38 34 3e 38 40 3c 3a 41 41 42 49 42 3e 44 41 49 47 40 43 47 40 43 36 3f 41 48 47 41 45 47 44 4a 4c 51 54 4a 40 3a 41 40 43 3b 3e 41 3d 3c 45 45 42 36 40 39 3e 3f 35 3d 46 43 45 40 3b 3e 3e 3e 38 3c 38 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 36 49 51 57 51 50 56 4b 4b 52 53 4a 51 50 56 59 59 5c 5b 5e 5e 58 56 4b 4d 50 50 4b 4f 4f 4e 51 43 4f 4e 52 47 4e 51 47 4f 5b 51 52 55 48 4b 4c 3c 41 42 40 39 46 3e 44 48 46 41 4b 49 46 4e 52 47 49 47 45 42 4a 3e 4e 45 45 4a 47 4b 4b 4e 4b 49 46 47 4b 4e 45 42 43 47 4b 46 2f 23 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 0b 12 26 28 2a 3c 43 4a 45 3c 47 3d 39 3b 2f 3b 35 42 3f 38 36 3b 36 3c 3b 36 3a 3f 38 38 46 3c 42 3c 43 42 42 3a 42 3c 44 49 4d 41 3f 41 44 42 41 3b 3f 42 3d 44 48 4b 43 46 4c 51 55 4b 46 47 40 3e 41 36 45 43 3a 3a 3f 43 3b 3e 3f 40 41 3e 43 3a 3f 3d 3c 37 41 3e 3d 39 35 36 3b 13 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 2d 49 54 53 50 51 52 51 4f 4b 56 4b 5a 52 4b 5b 58 5f 5f 58 59 52 57 54 4f 55 4a 56 48 52 46 4a 4a 4f 4c 50 54 50 54 54 4d 54 57 4e 4c 3f 49 43 3c 45 41 4c 49 42 4e 48 47 51 46 47 46 40 44 46 48 41 40 44 4f 48 46 48 48 42 4d 49 45 4b 49 51 4a 49 50 3f 49 4b 46 44 47 43 38 32 20 0c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0e 12 1c 26 2b 39 39 41 40 45 3c 44 3e 3c 3d 3d 44 3b 3e 39 3f 41 39 3d 36
 37 3d 3a 38 37 3e 37 3c 3b 42 3d 44 43 3c 3b 40 45 43 40 44 3b 3e 43 41 46 3a 3d 3e 42 49 4c 4b 46 4b 4b 58 48 45 3c 45 3d 3b 3e 43 44 46 37 41 3e 3e 38 44 44 3b 41 42 3c 38 47 3a 3f 40 40 37 39 3b 31 32 11 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 34 47 52 4f 4a 4b 4a 58 50 4f 52 4b 4e 53 52 54 5b 5f 56 55 52 52 53 54 4d 50 4b 4f 4c 4e 52 40 4e 53 51 4f 4c 4f 51 4e 59 55 52 4c 43 46 41 49 44 48 46 3d 47 4a 49 46 48 49 47 43 4c 3e 40 44 3f 49 4a 46 44 44 45 46 42 4a 48 45 48 4f 4c 45 4a 52 51 47 52 45 44 48 3b 41 34 25 16 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 06 05 10 12 1b 24 38 3c 3e 3a 44 3f 3d 42 3e 36 2b 36 3b 34 40 36 37 37 34 33 3b 35 3e 35 3b 37 32 40 41 3e 39 44 35 35 3b 3f 3b 3c 40 4b 3a 40 44 37 3e 3a 3c 37 3d 39 3d 44 4c 43 41 4b 43 3e 43 3f 40 37 45 3c 3d 43 37 42 3e 3d 32 35 3d 3e 3d 3c 41 3c 3b 3c 3b 3c 3a 46 39 3a 2f 34 1c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 26 41 3f 4a 58 4e 4d 4b 4a 51 53 4f 47 50 4f 53 58 5a 57 4e 56 4f 4b 51 53 51 4f 4d 4c 4b 45 4a 46 47 4b 44 4f 4e 4c 51 4c 4e 55 51 4a 41 41 41 45 3d 40 40 4a 46 47 42 44 41 3b 42 44 46 4e 49 42 46 3d 46 4c 49 3f 47 45 41 3d 51 4a 49 48 45 4f 4c 47 47 40 42 4a 44 3c 36 28 20 09 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 13 1a 21 26 31 33 34 3e 34 45 44 44 44 3d 3f 37 41 3b 3f 44 32 3f 39 3d 3a 3c 3b 3a 43 37 3b 33 33 4a 42 42 3f 3a 3e 3f 3f 3b 43 40 47 36 41 42 43 38 43 47 46 38 3f 3f 41 3e 43 4c 38 41 3b 36 38 41 3c 45 3b 43 39 43 38 39 43 3c 39 43 41 3e 3b 36 40 3c 40 3a 35 3b 35 31 38 36 1a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 1f 45 4f 50 53 4b 4b 4f 4a 53 4f 55 4b 51 55 5d 53 5f 52 54 56 4e 54 4a 50 4a 49 54 52 56 48 4e 4f 44 4b 53 4a 54 48 57 52 51 54 4f 4d 36 42 3d 43 43 4a 44 43 4f 48 4d 45 43 40 46 44 45 42 46 41 3d 3e 47 40 48 4b 46 4a 41 44 3f 48 44 4a 46 41 48 4c 4c 4d 46 43 40 2e 30 24 13 07 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 13 11 23 29 31 39 34 3b 2c 47 44 3f 3b 39 3a 39 3f 3a 35 3b 3b 33 37 3c
 3a 36 3e 38 3a 3d 37 40 34 34 3d 3c 35 42 3e 3e 3d 3d 42 45 40 49 4c 49 3e 45 3a 3b 39 33 40 3c 41 42 45 44 41 42 3f 44 49 46 47 41 43 49 37 40 41 3f 3a 42 3b 3e 40 3b 3e 3b 31 3c 38 38 3c 40 3b 33 38 2a 1d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 26 48 56 51 4c 4f 4c 51 4c 58 49 54 52 50 53 54 52 5c 60 56 5b 4f 52 57 4e 54 53 4e 51 53 44 50 4f 46 4f 4b 4c 4f 51 57 53 50 4a 42 40 3b 41 40 43 4a 3f 42 4a 41 48 4f 48 3d 4c 47 46 40 45 47 3f 41 46 44 45 47 40 41 44 43 53 45 47 4e 41 4f 45 4d 47 48 4d 4a 3c 44 39 25 25 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 17 15 20 25 2e 36 39 39 38 36 39 48 37 3d 3e 35 41 39 39 34 36 3a 38 33 37 31 3b 3d 34 34 31 38 33 34 33 37 3f 3e 36 3c 3d 3a 3c 43 3a 4a 4c 4c 48 43 45 3b 3d 3f 3e 3f 46 44 3b 3b 41 42 45 47 3f 3e 41 42 43 43 40 3b 3a 38 42 40 3d 3e 38 33 3f 2d 3c 34 37 36 37 38 34 38 2f 19 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1f 3e 51 52 51 49 4e 47 3d 53 50 48 48 4e 52 57 4e 4d 4f 54 56 53 4f 54 55 58 57 5c 4d 4b 4e 46 48 41 4d 56 4b 50 4f 51 4d 4b 3e 44 47 47 43 41 41 3f 49 44 42 46 49 4a 43 41 45 4b 46 50 40 46 44 46 47 41 42 44 3b 3b 3f 45 3d 3c 40 48 4e 48 43 45 40 3f 40 36 3e 37 26 24 0c 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 09 0e 16 25 33 36 38 3e 3f 3d 3b 36 41 35 37 36 38 3a 3d 34 31 39 35 37 3a 31 39 35 3d 32 3e 36 3d 3c 42 37 37 3b 3b 39 3a 43 34 3b 3e 36 44 42 42 3e 3d 3d 41 3f 45 3f 45 3e 40 42 4a 42 45 49 43 48 4d 3f 42 44 3b 3c 37 37 3d 3a 3c 36 38 3a 3a 3e 3f 2e 3a 2f 36 39 31 2e 32 25 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 26 47 55 4e 4a 4e 4e 46 52 4f 4b 46 45 48 56 51 53 50 56 4d 4e 50 4e 51 52 5b 59 5f 58 4f 4f 3f 45 48 53 4e 4e 54 4e 49 49 49 4f 4a 4e 3e 3e 45 3b 3d 3f 4a 3f 40 4d 45 46 47 41 41 42 3a 41 41 44 42 40 3d 41 46 3f 33 3e 46 41 42 43 47 40 45 4a 40 47 44 44 3c 3a 39 25 15 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 08 0e 14 2d 26 2c 33 39 36 3b 35 3e 3d 37 49 46 35 3d 42 3a 34 3c 3c
 37 3b 37 35 36 34 3c 3c 38 3b 34 39 36 3f 3d 39 40 3b 39 3d 42 38 3a 42 3d 40 48 41 3f 41 3c 39 41 40 41 46 43 47 45 44 4d 4f 4e 4e 3f 4a 37 3e 45 3b 3d 44 42 3a 33 3c 32 3b 35 32 32 30 39 37 42 37 38 30 1e 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 18 3f 4b 4f 4e 55 4c 51 55 50 4d 47 51 52 55 4f 4f 54 54 54 50 5a 50 58 53 52 4e 55 55 4e 51 4a 4a 56 4b 4b 56 47 50 4a 42 4c 41 41 4a 48 42 49 43 45 40 46 44 4a 4d 41 44 3e 41 49 46 45 45 47 40 44 41 40 3f 3c 3a 49 45 46 49 40 43 45 4a 43 41 3f 44 44 3d 3d 32 2d 22 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 0b 13 1d 2a 30 31 3a 43 3d 3a 37 37 45 40 43 42 3b 3d 36 3d 3d 40 32 37 3c 36 3e 3b 36 37 39 36 36 36 34 3f 3a 34 3c 37 3c 3c 32 39 38 3c 37 42 39 3d 41 46 3f 3e 3d 43 3e 3c 3f 43 4a 47 51 4e 53 4e 47 4b 38 39 3d 39 36 42 32 38 40 32 37 38 36 38 2e 37 36 35 39 34 2e 35 22 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 39 4e 45 53 49 47 50 49 4a 50 51 51 50 4f 39 4f 4e 50 55 4d 56 50 4f 5b 5f 58 66 57 55 4e 4b 54 51 53 4e 4d 49 3f 44 49 4c 4d 40 42 43 4b 49 45 43 47 41 45 46 47 44 41 45 40 43 45 40 36 45 3a 49 4a 41 44 3a 41 44 46 4f 44 46 44 41 43 44 41 48 48 45 40 2f 2d 22 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 14 17 29 31 40 38 41 43 3c 38 3a 3d 3c 3e 39 3b 3e 38 38 3a 38 38 3e 38 35 39 38 37 35 3f 32 38 40 39 38 36 3a 3c 38 3e 3c 38 32 3e 3e 3b 30 36 3a 39 3b 3a 37 3b 38 37 41 3d 3e 42 45 4a 4d 52 50 4e 4a 37 39 34 31 33 32 37 38 36 34 39 2f 38 3d 33 35 38 2f 30 2e 35 32 20 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 38 4b 4d 51 50 4b 52 4f 51 4a 50 42 45 45 4e 4c 4d 55 53 56 51 4b 57 5c 59 5e 5a 51 53 54 4a 4d 55 50 43 4a 49 4a 43 48 4c 41 4b 50 4d 4a 44 46 46 45 43 43 40 42 3d 40 40 3e 47 45 44 4a 43 3e 42 3d 42 47 3f 49 40 36 42 4a 41 3f 49 45 4c 44 39 3c 38 2f 38 29 15 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 07 14 13 21 32 33 38 40 43 3e 38 37 41 45 45 42 37 3d 39 35 36 3e
 36 3b 3a 34 32 37 39 35 39 3b 42 44 38 3e 36 34 44 3a 3e 3f 38 3b 35 32 3e 3b 3f 39 38 36 3a 43 44 3f 44 3b 41 3d 3e 49 42 47 51 4a 4e 44 36 39 3d 3a 3b 3c 37 35 31 37 2d 36 3a 38 30 37 39 37 31 33 3a 2e 23 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 33 50 50 53 4e 45 4b 43 47 50 49 4c 4e 55 54 4d 51 52 58 53 57 58 56 56 5b 55 64 5a 50 4c 49 53 47 4d 4d 4f 4c 47 45 54 48 50 4e 47 40 4a 4b 45 47 3e 40 48 41 3f 42 3d 3c 4a 40 3b 42 45 44 45 43 44 47 50 41 45 48 43 49 48 4c 44 4d 4a 46 3d 35 3b 3b 3e 26 20 1a 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 15 21 27 35 45 46 4d 44 3e 37 38 40 45 3f 42 42 34 42 36 37 34 36 36 39 36 3d 3d 3e 3a 3b 36 3f 3b 3f 3a 3e 34 33 36 3d 34 32 41 35 3c 36 36 33 32 3b 39 3a 3e 33 32 3d 33 39 3d 3e 42 3f 4c 47 46 42 3e 40 37 3c 3b 33 3c 39 3d 30 37 36 35 3d 34 3b 33 33 36 35 35 2c 29 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 34 4f 4d 51 46 49 4c 41 44 44 44 4e 51 48 52 50 4d 52 5a 4a 55 56 54 59 50 5b 61 5b 5b 58 4b 55 50 51 52 4e 4e 4d 54 4e 3f 54 4c 54 49 41 46 48 3a 49 3c 46 4b 40 45 42 43 3e 45 4e 3e 48 47 3e 40 47 44 4b 4e 59 52 52 54 4f 54 59 55 51 48 3e 48 37 3a 32 1f 20 0b 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 19 1d 2c 44 45 49 43 40 36 39 40 38 3b 3a 35 3e 39 39 38 37 37 35 32 3a 39 33 30 3c 34 40 3b 38 36 3b 44 3a 37 31 37 3c 3c 3a 34 33 2e 2f 37 37 32 36 36 36 36 38 37 32 2f 3a 3e 3a 41 45 44 47 3e 36 34 3b 33 31 30 2c 31 36 39 39 31 34 32 32 3a 36 3e 37 30 2e 30 25 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 2d 4a 47 47 49 47 4a 46 4c 42 40 4c 4f 45 52 4e 53 53 58 59 58 58 53 4c 51 55 5d 5e 58 4b 56 49 55 50 4c 59 4f 52 46 4c 4c 4d 49 49 4d 4c 48 37 3f 3f 37 40 3e 44 43 3d 48 47 4a 4a 4a 42 44 45 50 59 60 59 59 4e 68 59 5a 6a 55 66 5b 5b 54 47 46 36 35 2a 1f 15 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 0b 1b 2e 33 51 53 48 42 38 3a 3d 39 44 43 3b 34 37 31 31
 35 3a 35 37 34 3d 36 3e 37 3a 3c 3e 39 39 36 3d 3a 3b 3a 39 3b 3c 33 38 34 30 39 36 31 36 35 3a 38 31 38 3c 32 34 3a 33 41 35 42 41 3a 3a 34 39 3e 3a 37 32 34 34 35 3c 35 31 37 36 33 41 36 36 31 2b 34 31 28 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 31 41 41 4f 47 43 4e 3c 41 4a 4b 4a 4c 52 4e 53 4d 4b 53 50 5b 53 52 4e 4e 58 52 54 56 4f 54 54 59 56 5a 5b 57 53 4e 4e 4c 4e 48 52 4b 4d 44 45 44 40 46 3d 3b 45 46 41 46 4c 49 4c 51 4d 56 55 58 5b 62 6b 69 65 65 64 6a 68 69 6b 60 5a 48 23 32 37 36 25 16 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 1e 26 40 42 52 5a 4a 3d 3c 38 3d 3d 2c 3b 37 2f 3e 34 37 35 3d 35 30 3a 3d 3a 37 42 39 37 3b 33 43 3a 35 3c 33 3a 35 3d 3a 35 30 36 37 39 30 38 33 34 3b 38 30 39 3a 36 36 3a 38 37 3d 32 38 3c 39 37 35 34 37 37 31 37 31 34 39 3c 30 32 38 38 2d 31 36 34 2f 29 29 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 26 3c 41 4a 49 4a 47 3b 3b 4a 45 4b 54 4e 52 46 4d 4d 4f 4f 50 4f 42 47 49 4c 4d 49 53 53 4f 53 4d 54 52 5a 52 55 52 55 56 55 48 4d 4b 44 48 3e 3d 46 44 40 45 45 45 47 56 4e 61 56 60 5a 65 64 6d 72 72 7d 6a 68 73 6c 6d 6e 6a 63 65 5b 56 48 3e 2d 2c 1b 0b 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 10 1b 2b 3d 4b 4e 49 48 3c 35 38 34 3a 40 39 36 3a 39 3c 36 3a 35 3a 3a 3b 35 3b 34 35 3a 36 3e 40 34 36 31 3e 38 39 34 28 35 36 3b 34 2b 37 30 32 34 33 35 34 2f 39 34 2f 33 34 39 39 40 3b 31 35 35 3b 32 31 32 2c 2f 35 33 2a 30 35 37 2d 38 3b 30 33 33 31 2f 25 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 42 45 46 40 40 42 3e 47 43 43 39 46 4a 48 4a 4a 4b 46 3f 46 43 45 45 45 49 4f 49 4f 4c 4f 4c 57 52 54 55 51 58 55 54 49 47 49 4c 4e 4d 4c 47 4c 43 4a 54 50 52 4e 52 5a 5e 66 67 6c 79 71 6e 74 73 7c 76 78 74 74 6c 6a 6d 68 6c 5e 60 54 44 43 27 1c 13 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 16 25 37 47 54 55 42 38 3e 32 3c 36 34 34 31 3c 39
 3c 3a 2e 36 3a 3d 34 35 3a 40 3e 3b 3d 3e 39 39 36 39 3e 37 34 35 34 35 3e 34 34 32 28 33 32 36 39 30 35 37 38 33 34 3e 2c 32 35 35 30 2f 2d 31 3a 36 3a 30 37 34 33 39 30 2e 36 34 33 38 35 36 32 35 32 2a 2b 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1f 38 3c 43 43 37 48 40 46 42 43 41 3d 4a 44 4a 46 45 45 47 48 43 3e 43 43 3e 4c 4b 4b 49 4e 4d 50 50 54 56 4d 4f 45 47 4a 4b 4e 4f 49 51 47 50 49 4f 54 61 5e 65 72 68 7a 72 75 74 72 75 77 77 74 75 71 6f 76 77 6d 6b 71 6a 6d 6b 5c 61 54 45 38 24 18 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 1b 2d 38 42 4a 4f 41 3f 38 34 35 39 34 36 38 32 32 2f 2d 36 3c 36 37 3a 30 37 37 37 36 37 36 37 30 3d 33 37 33 35 38 37 37 31 39 30 36 31 35 36 33 30 37 3b 29 34 35 2e 2e 36 36 38 31 3d 2e 35 30 2f 38 35 2e 39 2e 33 35 30 34 34 34 2f 2e 3b 2b 36 34 36 29 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 37 44 44 3d 3a 3f 3c 3a 41 39 3c 42 3c 42 3e 45 44 45 45 45 41 47 45 3f 3f 40 42 4e 48 46 44 46 48 55 4b 49 47 4a 50 4f 54 51 4e 56 54 58 5b 5f 66 6b 6c 72 72 70 6b 76 7a 83 7b 75 79 73 72 7a 74 75 70 6d 67 6f 64 6f 64 68 60 63 62 4d 3f 36 1b 0b 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 0e 14 23 35 42 48 4b 47 3a 32 2f 32 37 32 36 3d 32 3b 37 35 34 38 32 32 32 35 39 2d 36 37 35 3e 33 2f 36 37 3c 35 3d 39 32 3d 38 38 34 33 33 2c 35 31 39 2f 34 39 2c 2b 33 2d 2f 34 33 36 35 31 35 33 30 32 31 35 2f 33 31 2f 2c 36 37 32 38 31 32 34 31 38 33 30 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1b 34 42 3c 3b 3c 41 3a 3e 38 3b 42 41 3c 3c 39 3d 3c 3c 42 3e 3e 42 3c 44 3c 40 42 3f 42 3b 3f 45 3d 49 49 45 44 48 4f 50 52 5d 62 60 67 6b 67 6b 75 76 7b 6b 76 75 78 75 78 74 76 71 76 73 70 6c 74 6d 6a 6b 60 69 64 6b 74 64 65 5d 56 4a 39 22 14 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 19 27 2e 45 4a 4d 3d 36 37 32 35 41 3b 36 35
 3d 33 3a 3e 2c 39 34 39 38 3f 34 38 38 3a 36 3c 36 34 36 3c 32 35 32 36 39 3b 35 32 30 34 31 35 2a 2d 32 39 2e 30 35 32 39 2f 34 33 2c 34 30 34 38 2e 37 33 2e 2f 32 36 31 2a 38 3e 44 35 35 34 33 39 33 35 2c 1d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 31 44 45 3c 37 3e 32 38 3e 3d 35 3b 35 38 36 3e 3e 45 3c 44 3b 3b 42 44 35 3c 35 41 3a 40 41 3d 43 4a 4c 50 55 56 5c 67 65 68 76 73 75 75 75 7c 7b 74 7c 76 7a 77 77 79 75 7e 7c 77 74 69 6a 71 71 64 6c 6b 66 6f 64 60 69 64 5f 5d 55 43 28 1c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 15 2c 3b 43 4a 3c 3a 35 33 3a 33 38 2e 34 33 3b 38 36 37 36 35 36 37 39 36 35 3c 3b 32 40 35 36 39 37 34 35 3a 37 40 35 37 2f 30 35 30 36 37 36 34 30 32 32 32 2c 32 2e 31 34 34 34 2c 2d 33 35 2f 35 38 2d 33 2c 35 32 34 41 40 42 37 33 38 37 34 39 36 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 15 32 42 3e 3c 2e 3b 34 32 32 37 39 31 42 3d 2f 36 40 3a 3d 41 3d 44 42 39 3a 3e 3b 39 3f 39 43 4e 44 4b 51 5f 5a 68 6f 72 7b 83 80 7d 75 7e 7c 79 7e 78 81 7b 76 7d 7a 75 74 75 77 73 73 6b 6f 6f 67 68 68 6c 6c 66 5b 6a 63 5a 5f 59 4b 39 1a 11 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0f 23 22 37 41 3c 39 36 35 30 33 30 2a 31 37 42 31 39 32 3a 37 30 35 39 34 35 32 3b 31 35 2b 36 31 36 35 31 39 37 37 3b 2e 34 32 2c 2f 32 31 2f 2d 2e 35 31 2a 35 2f 28 25 32 2c 2f 31 35 30 2e 2d 30 31 39 2b 29 35 2c 2f 32 3d 3c 39 37 35 34 34 38 34 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1a 2d 2f 39 3e 34 3b 31 34 33 32 35 39 3b 3b 35 30 38 3d 3d 3d 32 3c 3a 3a 36 3b 3d 41 3a 3e 42 51 58 60 62 6f 6a 7d 76 78 7e 7f 84 79 7e 80 7f 7d 7c 78 7a 76 73 79 74 70 70 6d 6c 65 69 6e 64 63 68 60 67 73 6b 66 61 63 64 60 55 4d 3c 28 17 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 19 22 2f 33 3b 39 41 3a 39 37 2f 3b 35
 33 36 35 3a 35 39 33 36 34 35 31 2f 31 36 3a 36 32 34 3e 35 39 39 31 34 39 34 2e 2c 28 30 35 34 2f 2e 2d 30 36 37 2c 2b 2f 2e 2d 36 2f 2e 21 2c 33 32 37 39 2c 33 2b 2d 32 32 2d 2c 33 34 36 38 35 34 34 40 2a 1a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 34 31 34 37 32 3e 37 36 3b 37 37 30 35 2f 3a 3b 39 36 3d 33 2c 31 3e 3f 37 3b 38 49 48 4a 55 63 6c 74 79 7b 84 83 7c 7c 84 85 7f 78 8a 79 72 79 7d 7a 73 74 77 7a 71 6f 6f 67 6d 66 6d 5f 64 62 59 5d 5c 63 6a 62 5c 62 60 5c 51 3a 2c 21 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 12 19 1f 34 2a 3c 34 33 3f 38 35 3a 34 37 3c 39 36 35 37 2d 39 35 3c 35 2d 33 34 2d 30 39 2f 2f 38 30 36 2e 37 36 2e 2f 2d 35 34 30 2f 2c 35 30 37 2d 33 33 30 39 30 34 2c 2c 34 34 2e 36 2b 2e 30 2d 2c 30 2d 2b 31 36 36 34 35 32 27 33 2f 31 30 2e 1c 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 2b 33 3a 3b 32 38 33 31 3a 3a 2e 3d 32 38 38 32 36 3a 35 36 39 36 37 39 44 4a 45 4a 55 66 6d 73 7d 7c 76 7c 7a 74 87 84 80 83 7f 7b 84 77 78 7b 75 76 71 76 72 6e 72 69 6f 64 6d 66 65 48 5c 5f 5e 60 68 5f 64 68 5f 5a 55 54 44 30 1a 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 11 1f 22 2d 31 39 39 35 37 2f 33 2d 3c 38 34 3d 3a 39 38 2d 2f 34 30 39 33 36 30 3a 2f 3c 34 32 2c 2e 32 2d 32 3a 32 35 2b 2e 2b 30 2a 30 2f 28 1e 34 29 31 2e 29 30 30 33 2b 2f 28 2b 2c 2c 35 2c 2f 31 25 2d 26 26 2c 2f 2b 21 25 2e 2d 36 2c 2d 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 1d 33 32 34 2a 39 28 3f 3a 2e 33 32 33 3d 3f 38 35 36 36 36 36 3f 46 42 48 55 56 64 73 72 7f 7f 7d 80 7d 7a 85 7b 80 7c 7e 7a 79 74 75 7c 78 73 74 71 6b 70 63 65 67 61 63 67 5a 5f 65 5e 65 62 56 5b 5f 5e 5a 64 53 50 48 3c 2b 1b 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 11 1e 30 2c 2e 32 40 35 3a 36 38
 34 3b 3a 37 37 33 33 31 33 30 38 34 37 33 33 2f 29 32 30 34 38 36 34 2f 2b 2d 31 34 30 31 2c 31 2d 31 33 35 2b 25 26 2d 2f 37 2c 26 2a 26 30 2e 2c 26 2e 29 2e 30 2d 25 29 2d 31 37 2a 27 2c 27 28 29 29 27 21 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 26 34 35 32 28 2c 33 30 29 35 2e 2f 36 2e 32 3d 31 34 3d 36 46 4c 4c 54 56 65 64 78 78 79 7c 81 7f 7c 85 7e 84 84 80 7f 74 80 82 7c 7d 72 6f 6f 6e 70 68 70 69 65 61 61 65 5f 60 57 65 55 5c 5f 57 54 5b 5b 59 53 50 4c 40 3b 20 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 06 13 25 27 36 2f 3a 37 39 39 2f 39 2f 38 35 39 3e 38 35 3c 38 31 32 36 32 37 3a 2c 2e 31 3a 30 36 31 33 34 34 36 32 28 2d 2d 36 31 2e 30 31 2e 2b 30 2c 2e 25 2f 2d 2a 2f 30 2b 29 26 2a 2a 2d 2e 2b 1e 29 29 31 2e 25 2a 25 2a 26 2a 25 26 28 22 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 2f 35 3a 32 2c 31 34 30 2e 33 33 34 35 36 31 3f 3d 44 35 4e 52 5b 67 72 71 83 7b 70 81 7c 86 7e 7d 7f 7d 7d 7e 7b 80 71 75 7c 6e 7d 72 6a 6f 6c 6c 6d 65 69 66 6a 63 59 65 59 5e 5b 59 59 62 5e 58 5f 58 57 51 4a 41 36 24 11 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 1d 20 2b 2d 2f 38 37 36 35 37 39 3e 3b 3c 46 39 3b 33 2f 34 32 34 34 38 3b 32 35 36 37 2f 34 29 30 37 30 34 29 2c 28 2d 2e 31 30 35 30 24 29 2a 2f 32 2a 26 30 2a 23 26 2a 2e 2e 28 26 29 2a 30 29 28 25 2c 28 22 31 25 24 29 23 21 26 19 20 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1d 29 33 2e 2d 32 2b 2f 31 27 31 36 30 35 35 38 3b 46 4f 54 5c 64 60 6f 7a 76 79 75 7a 7d 79 7c 7d 7f 79 74 76 72 70 71 6f 71 6f 6c 70 6c 69 69 6b 64 5c 61 5e 59 59 5b 54 5d 59 57 54 5f 4d 4e 52 4f 61 50 52 49 3b 32 23 10 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 17 25 28 31 2e 2e 35 34
 38 36 32 3c 39 38 35 36 3d 3a 32 33 33 2f 2f 37 32 3d 31 35 33 35 37 2a 32 2d 2b 30 30 21 24 39 2e 2f 2e 32 30 2e 26 29 2b 29 26 2b 2c 2f 21 29 22 27 24 20 26 2a 28 26 2a 26 24 2a 29 2d 24 2c 21 20 25 23 26 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 18 2b 27 30 2f 2c 24 2e 29 20 30 34 2e 3f 3e 3d 47 50 5a 5a 66 76 63 70 79 75 6b 74 6c 6b 71 6e 76 74 6a 6b 6f 72 6e 64 72 6e 6d 64 64 6b 5d 63 61 5f 5c 5a 53 51 55 54 4f 57 58 4b 4d 4a 55 56 55 4f 49 45 3a 3b 20 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 13 19 24 30 33 39 38 3a 33 37 3a 3d 3b 44 39 36 3c 36 38 33 2f 3c 34 2e 35 34 31 35 2b 34 36 34 30 31 2f 34 39 34 34 27 28 28 34 2f 27 23 2d 32 2b 2b 2c 27 21 29 23 2a 28 24 23 24 29 2a 29 24 2d 20 2d 29 21 27 24 29 21 24 20 24 24 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 10 24 27 27 35 2f 2c 2c 2f 2e 2f 3c 42 50 4a 57 50 5b 61 66 6a 68 66 6a 69 68 6d 6e 69 68 69 6d 6b 68 65 67 5e 5a 6e 61 66 5b 62 62 5e 55 56 5f 5d 59 54 55 52 52 4a 50 4e 4f 46 47 49 4f 47 51 50 40 44 39 29 21 12 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 13 1e 26 2d 29 2f 33 38 3a 33 3b 3f 3d 30 30 36 40 32 30 36 38 36 37 33 33 37 36 2c 35 30 2f 32 2d 28 34 30 26 2f 31 35 28 29 2b 2a 2f 2a 25 25 22 28 26 25 21 15 1a 25 21 1e 26 24 2c 27 28 2a 2a 1e 29 23 23 27 1f 21 1e 26 22 19 1e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 1d 26 1f 1e 23 23 24 26 27 36 3b 4c 48 49 52 5a 50 4d 53 5b 5d 5b 60 58 5e 5d 5c 58 51 51 56 5f 55 54 53 54 57 58 4f 55 4d 4f 4f 4c 4a 46 46 45 45 44 45 4a 40 3e 4b 49 42 46 45 44 4b 3b 39 3a 36 30 26 1e 0e 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 10 1d 1e 2e 2c 2c
 39 3b 31 32 33 37 39 32 31 33 30 32 2c 30 35 32 2f 30 34 35 32 32 2e 25 2c 2f 2c 29 31 24 27 2d 33 23 26 2c 1e 22 23 24 29 21 22 23 18 15 08 14 13 14 1a 1f 22 26 28 23 25 1c 22 23 16 1f 22 22 1e 18 1a 1e 16 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 16 18 16 14 22 22 2b 2f 33 39 36 36 39 38 38 35 49 43 3e 46 43 44 39 45 44 3e 3b 34 40 3c 3b 3c 39 3b 35 37 33 35 37 3c 38 3c 38 41 32 33 34 34 38 32 30 34 30 2f 2e 3a 32 32 35 31 2d 30 2a 1f 13 09 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 1a 14 2b 2d 2f 30 32 33 35 3e 3e 34 38 35 36 38 32 29 30 34 3a 33 31 3d 34 34 2f 31 2b 2f 32 2b 2c 2a 25 26 30 2b 21 2e 25 30 28 21 28 26 21 20 21 0f 0c 06 0f 11 11 15 1f 23 1d 22 25 1c 24 1f 21 1b 1e 21 1d 16 16 15 11 13 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 10 0d 11 13 18 23 25 24 23 26 31 27 30 2b 2e 27 2b 2c 26 30 2a 2f 2d 21 25 2d 25 29 2a 2c 28 2b 29 29 29 23 25 26 25 27 25 28 26 2e 23 1e 2c 21 27 22 22 2d 22 20 1d 22 26 1e 19 1e 12 13 0d 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 16 1b 1b 24 34 35 32 32 34 38 31 33 38 38 35 34 37 32 34 34 2e 32 39 39 2e 2d 32 2a 37 33 2a 26 29 25 27 25 25 1d 28 27 27 24 27 24 23 22 1d 19 12 03 06 05 09 04 10 0a 16 1c 1f 1f 15 15 17 12 09 13 0d 0a 13 0f 0c 0a 0c 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 06 0d 11 1e 1d 16 12 18 16 17 14 11 22 1a 16 16 1c 1a 1f 1e 18 25 1c 1a 11 15 15 12 13 1a 18 14 17 17 12 10 15 18 1c 1e 11 15 1a 10 0e 16 14 19 13 19 1a 19 11 11 1a 0b 13 0d 03 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 19 17 27
 27 2d 2b 32 30 2b 34 36 36 32 2b 32 2f 2f 2a 30 35 31 38 33 2d 33 27 2c 26 24 22 22 26 15 28 1f 1b 17 1e 25 19 19 13 14 1a 18 0e 09 04 00 06 05 03 00 06 05 0a 0b 06 0b 0a 04 06 0c 05 0c 06 05 07 00 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 0a 05 03 04 06 05 03 03 08 05 05 00 06 05 04 0c 06 13 05 06 07 13 0c 04 06 07 03 05 06 05 09 02 06 05 0d 01 06 05 03 0a 06 08 0a 06 06 07 03 04 06 09 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 11 20 21 2d 2b 29 2f 2f 38 39 38 36 33 34 2d 2f 31 2a 28 26 2a 28 27 2a 23 21 25 1c 12 14 1a 1b 17 19 1a 21 19 19 11 18 12 14 0c 0c 0d 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0e 21 20 24 25 2c 25 2c 35 36 30 2f 24 33 24 29 22 22 20 25 29 22 1d 20 1e 16 12 11 0b 05 0d 0a 0e 0b 0e 0d 0f 08 00 0b 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 0a 0a 14 1d 1d 24 25 2a 25 30 20 29 25 23 1f 21 17 15 1a 0f 10 12 19 08 0d 04 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 0f 0f 20 1a 13 20 1b 1f 1e 11 16 0f 0c 0b 09 06 09 04 04 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 03 00 06 0f 07 12 07 05 08 08 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
