 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04 05 05 05 05 05 05 05 05 05 05 05 05 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 03 03 03 05 05 05 05 05 05 04 04 04 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03 04 04 04 04 04 04 03 03 03 04 04 04 04 04 04 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 08 08 08 07 07 07 05 05 05 05 05 05 04 04 04 04 04 04 05 05 05 05 05 05 07 07 07 06 06 06 05 05 05 05 05 05 05 05 05 05 05 05 04 04 04 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04 05 05 05 07 07 07 05 05 05 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 06 06 06 0a 0a 0a 0e 0e 0e 0c 0c 0c 09 09 09 08 08 08 07 07 07 07 07 07 09 09 09 08 08 08 0b 0b 0b 0a 0a 0a 08 08 08 09 09 09 08 08 08 06 06 06 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 05 04 04 04 09 09 09 0a 0a 0a 07 07 07 05 05 05 04 04 04 04 04 04 05 05 05 05 05 05 04 04 04 03 03 03 04 04 04 05 05 05 05 05 05 04 04 04 04 04 04 04 04 04 04 04 04
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 05 05 05 05 05 05 04 04 04 04 04 04 05 05 05 07 07 07 0b 0b 0b 0e 0e 0e 12 12 12 11 11 11 0d 0d 0d 0d 0d 0d 0e 0e 0e 0c 0c 0c 0f 0f 0f 0e 0e 0e 10 10 10 0f 0f 0f 0e 0e 0e 12 12 12 0f 0f 0f 0e 0e 0e 0b 0b 0b 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 07 0b 0b 0b 0a 0a 0a 09 09 09 07 07 07 05 05 05 05 05 05 06 06 06 06 06 06 05 05 05 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 03 03 03 05 05 05 05 05 05 07 07 07 0b 0b 0b 08 08 08 06 06 06 07 07 07 0d 0d 0d 12 12 12 16 16 16 1b 1b 1b 1b 1b 1b 1c 1c 1c 19 19 19 1b 1b 1b 21 21 21 25 25 25 21 21 21 1b 1b 1b 1d 1d 1d 23 23 23 2f 2f 2f 2d 2d 2d 2b 2b 2b 25 25 25 1c 1c 1c 19 19 19 15 15 15 10 10 10 0f 0f 0f 11 11 11 15 15 15 10 10 10 0c 0c 0c 0c 0c 0c 09 09 09 07 07 07 09 09 09 08 08 08 05 05 05 04 04 04 05 05 05 04 04 04 03 03 03 04 04 04 04 04 04 04 04 04 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 06 06 06 07 07 07 06 06 06 05 05 05 05 05 05 07 07 07 09 09 09 0a 0a 0a 0b 0b 0b 0c 0c 0c 0d 0d 0d 11 11 11 16 16 16 1e 1e 1e 26 26 26 30 30 30 40 40 40 56 56 56 5f 5f 5f 66 66 66 91 91 91 88 88 88 76 76 76 5d 5d 5d 65 65 65 89 89 89 90 90 90 90 90 90 7b 7b 7b 66 66 66 54 54 54 5a 5a 5a 5b 5b 5b 48 48 48 3e 3e 3e 37 37 37 29 29 29 1f 1f 1f 19 19 19 15 15 15 10 10 10 0c 0c 0c 0d 0d 0d 0c 0c 0c 09 09 09 05 05 05 05 05 05 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04 04
 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 05 05 05 05 05 05 07 07 07 09 09 09 08 08 08 08 08 08 08 08 08 0c 0c 0c 11 11 11 13 13 13 15 15 15 16 16 16 20 20 20 30 30 30 48 48 48 60 60 60 7b 7b 7b b4 b4 b4 e0 e0 e0 f6 f6 f6 ed ed ed ca ca ca e0 e0 e0 d7 d7 d7 d2 d2 d2 d1 d1 d1 db db db d8 d8 d8 ba ba ba be be be c7 c7 c7 a6 a6 a6 92 92 92 98 98 98 a1 a1 a1 9d 9d 9d 8c 8c 8c 7c 7c 7c 71 71 71 71 71 71 5c 5c 5c 3e 3e 3e 2e 2e 2e 1d 1d 1d 15 15 15 10 10 10 09 09 09 05 05 05 04 04 04 03 03 03 03 03 03 04 04 04 04 04 04 04 04 04 04 04 04
 03 03 03 03 03 03 03 03 03 04 04 04 07 07 07 0b 0b 0b 09 09 09 09 09 09 0a 0a 0a 09 09 09 09 09 09 0c 0c 0c 14 14 14 1c 1c 1c 21 21 21 31 31 31 54 54 54 75 75 75 79 79 79 90 90 90 b3 b3 b3 b3 b3 b3 ae ae ae b2 b2 b2 b8 b8 b8 d6 d6 d6 fe fe fe fc fc fc eb eb eb e0 e0 e0 f6 f6 f6 fb fb fb dc dc dc c8 c8 c8 b5 b5 b5 a4 a4 a4 99 99 99 9f 9f 9f aa aa aa ae ae ae a6 a6 a6 a0 a0 a0 b1 b1 b1 c5 c5 c5 d6 d6 d6 a8 a8 a8 7e 7e 7e 81 81 81 6d 6d 6d 42 42 42 1f 1f 1f 0d 0d 0d 06 06 06 05 05 05 04 04 04 04 04 04 04 04 04 04 04 04 03 03 03 03 03 03
 04 04 04 04 04 04 04 04 04 05 05 05 09 09 09 12 12 12 13 13 13 10 10 10 0c 0c 0c 0e 0e 0e 10 10 10 16 16 16 22 22 22 39 39 39 57 57 57 8c 8c 8c 9d 9d 9d b2 b2 b2 c4 c4 c4 d3 d3 d3 e7 e7 e7 e4 e4 e4 cf cf cf c4 c4 c4 be be be bf bf bf d9 d9 d9 e3 e3 e3 dc dc dc ce ce ce d5 d5 d5 d2 d2 d2 c7 c7 c7 c4 c4 c4 bf bf bf b9 b9 b9 b4 b4 b4 b3 b3 b3 b7 b7 b7 b9 b9 b9 ba ba ba b7 b7 b7 bc bc bc db db db e4 e4 e4 b8 b8 b8 a9 a9 a9 b5 b5 b5 b5 b5 b5 a9 a9 a9 78 78 78 2f 2f 2f 15 15 15 09 09 09 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 04 04 04 07 07 07 07 07 07 0a 0a 0a 11 11 11 1b 1b 1b 1c 1c 1c 1b 1b 1b 17 17 17 16 16 16 1c 1c 1c 2e 2e 2e 51 51 51 73 73 73 99 99 99 ba ba ba ce ce ce e7 e7 e7 f7 f7 f7 fd fd fd fc fc fc f7 f7 f7 e5 e5 e5 cf cf cf c0 c0 c0 b7 b7 b7 bb bb bb c2 c2 c2 c4 c4 c4 c8 c8 c8 cc cc cc d2 d2 d2 d1 d1 d1 d7 d7 d7 cd cd cd c3 c3 c3 b9 b9 b9 ba ba ba bb bb bb bd bd bd c1 c1 c1 c1 c1 c1 c9 c9 c9 d1 d1 d1 ce ce ce c5 c5 c5 bd bd bd b5 b5 b5 aa aa aa af af af ae ae ae 74 74 74 2f 2f 2f 12 12 12 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 09 09 09 0c 0c 0c 10 10 10 14 14 14 1b 1b 1b 22 22 22 21 21 21 25 25 25 26 26 26 26 26 26 41 41 41 6a 6a 6a 7f 7f 7f a7 a7 a7 e0 e0 e0 e7 e7 e7 ec ec ec f5 f5 f5 fa fa fa f8 f8 f8 f8 f8 f8 fc fc fc f2 f2 f2 e0 e0 e0 cd cd cd bf bf bf bb bb bb c5 c5 c5 cc cc cc cd cd cd d0 d0 d0 d4 d4 d4 d8 d8 d8 e6 e6 e6 e2 e2 e2 d7 d7 d7 c0 c0 c0 bc bc bc c5 c5 c5 cf cf cf d5 d5 d5 d0 d0 d0 d1 d1 d1 d2 d2 d2 ca ca ca c3 c3 c3 c1 c1 c1 c3 c3 c3 c1 c1 c1 b4 b4 b4 ab ab ab 85 85 85 6a 6a 6a 34 34 34 0d 0d 0d 05 05 05 04 04 04 04 04 04 03 03 03 03 03 03
 0f 0f 0f 12 12 12 19 19 19 1e 1e 1e 24 24 24 28 28 28 27 27 27 29 29 29 31 31 31 50 50 50 9d 9d 9d c0 c0 c0 cb cb cb eb eb eb f9 f9 f9 f3 f3 f3 f2 f2 f2 f6 f6 f6 f8 f8 f8 f9 f9 f9 fc fc fc fd fd fd fc fc fc f3 f3 f3 e0 e0 e0 ce ce ce ca ca ca d4 d4 d4 db db db d6 d6 d6 d5 d5 d5 d9 d9 d9 e0 e0 e0 f3 f3 f3 f4 f4 f4 ea ea ea ce ce ce cf cf cf df df df eb eb eb ee ee ee ed ed ed e5 e5 e5 dd dd dd d8 d8 d8 ce ce ce ca ca ca c5 c5 c5 c3 c3 c3 b8 b8 b8 af af af 90 90 90 81 81 81 79 79 79 25 25 25 09 09 09 04 04 04 04 04 04 03 03 03 03 03 03
 16 16 16 1a 1a 1a 20 20 20 25 25 25 2b 2b 2b 2e 2e 2e 2e 2e 2e 36 36 36 59 59 59 c9 c9 c9 f7 f7 f7 ee ee ee f7 f7 f7 fe fe fe f0 f0 f0 e6 e6 e6 f8 f8 f8 fb fb fb fa fa fa fd fd fd fe fe fe fe fe fe ff ff ff fd fd fd f1 f1 f1 e2 e2 e2 d9 d9 d9 d8 d8 d8 e2 e2 e2 e1 e1 e1 de de de e5 e5 e5 ef ef ef f6 f6 f6 f8 f8 f8 ee ee ee e0 e0 e0 ea ea ea f9 f9 f9 fd fd fd fd fd fd fd fd fd fa fa fa f2 f2 f2 eb eb eb e0 e0 e0 d2 d2 d2 c6 c6 c6 be be be b0 b0 b0 a5 a5 a5 9c 9c 9c 8b 8b 8b 8b 8b 8b 5f 5f 5f 17 17 17 05 05 05 04 04 04 03 03 03 03 03 03
 1c 1c 1c 21 21 21 26 26 26 29 29 29 2d 2d 2d 32 32 32 37 37 37 4d 4d 4d 9d 9d 9d ce ce ce f5 f5 f5 fd fd fd f8 f8 f8 e9 e9 e9 d2 d2 d2 d2 d2 d2 ed ed ed fd fd fd fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 ee ee ee e2 e2 e2 e1 e1 e1 f0 f0 f0 f7 f7 f7 f7 f7 f7 fb fb fb fb fb fb f8 f8 f8 fd fd fd f7 f7 f7 f5 f5 f5 fc fc fc fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc f6 f6 f6 eb eb eb e1 e1 e1 d6 d6 d6 cd cd cd b8 b8 b8 a2 a2 a2 96 96 96 8c 8c 8c 92 92 92 8c 8c 8c 37 37 37 09 09 09 04 04 04 04 04 04 03 03 03
 1e 1e 1e 23 23 23 2a 2a 2a 2d 2d 2d 2e 2e 2e 34 34 34 41 41 41 76 76 76 a8 a8 a8 a5 a5 a5 be be be d7 d7 d7 d3 d3 d3 d3 d3 d3 da da da db db db eb eb eb fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fc fc fc fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd fb fb fb f4 f4 f4 f0 f0 f0 e8 e8 e8 d8 d8 d8 c4 c4 c4 b1 b1 b1 a1 a1 a1 97 97 97 99 99 99 93 93 93 4f 4f 4f 12 12 12 07 07 07 04 04 04 03 03 03
 20 20 20 26 26 26 2c 2c 2c 2d 2d 2d 32 32 32 3e 3e 3e 57 57 57 8f 8f 8f a2 a2 a2 a9 a9 a9 b4 b4 b4 cf cf cf d8 d8 d8 dd dd dd eb eb eb f8 f8 f8 fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fd fd fd f9 f9 f9 f4 f4 f4 ee ee ee e1 e1 e1 d1 d1 d1 bf bf bf ac ac ac a1 a1 a1 9a 9a 9a 8c 8c 8c 66 66 66 2c 2c 2c 0e 0e 0e 06 06 06 03 03 03
 21 21 21 24 24 24 2d 2d 2d 30 30 30 3b 3b 3b 54 54 54 6a 6a 6a 92 92 92 a9 a9 a9 b8 b8 b8 bb bb bb d0 d0 d0 e2 e2 e2 ea ea ea f7 f7 f7 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f9 f9 f9 f1 f1 f1 e8 e8 e8 de de de d0 d0 d0 c1 c1 c1 b0 b0 b0 a4 a4 a4 90 90 90 73 73 73 68 68 68 3f 3f 3f 0e 0e 0e 03 03 03 03 03 03
 1e 1e 1e 22 22 22 2c 2c 2c 32 32 32 42 42 42 64 64 64 7f 7f 7f 8a 8a 8a a1 a1 a1 c1 c1 c1 c7 c7 c7 d3 d3 d3 e6 e6 e6 f7 f7 f7 fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd fb fb fb f6 f6 f6 ee ee ee e2 e2 e2 d2 d2 d2 c3 c3 c3 b4 b4 b4 a8 a8 a8 97 97 97 79 79 79 6a 6a 6a 63 63 63 44 44 44 11 11 11 03 03 03 03 03 03
 1b 1b 1b 24 24 24 28 28 28 2e 2e 2e 3d 3d 3d 67 67 67 85 85 85 7f 7f 7f 8d 8d 8d b5 b5 b5 c8 c8 c8 d4 d4 d4 e5 e5 e5 f7 f7 f7 fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fa fa fa f3 f3 f3 ed ed ed eb eb eb e3 e3 e3 d6 d6 d6 c8 c8 c8 ba ba ba ab ab ab 9f 9f 9f 84 84 84 69 69 69 61 61 61 60 60 60 48 48 48 13 13 13 03 03 03 03 03 03
 18 18 18 21 21 21 25 25 25 29 29 29 38 38 38 63 63 63 80 80 80 7c 7c 7c 81 81 81 9d 9d 9d bd bd bd ce ce ce db db db ed ed ed fb fb fb fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd fd fd f1 f1 f1 e1 e1 e1 da da da d9 d9 d9 d8 d8 d8 d1 d1 d1 c5 c5 c5 bb bb bb af af af a0 a0 a0 8f 8f 8f 6c 6c 6c 62 62 62 5f 5f 5f 5e 5e 5e 49 49 49 12 12 12 03 03 03 03 03 03
 19 19 19 1e 1e 1e 1e 1e 1e 24 24 24 36 36 36 65 65 65 87 87 87 7b 7b 7b 78 78 78 88 88 88 a5 a5 a5 c5 c5 c5 d4 d4 d4 e5 e5 e5 f5 f5 f5 fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f8 f8 f8 e1 e1 e1 cc cc cc c4 c4 c4 c4 c4 c4 c3 c3 c3 bd bd bd b5 b5 b5 ac ac ac a1 a1 a1 95 95 95 75 75 75 65 65 65 60 60 60 5b 5b 5b 5d 5d 5d 46 46 46 11 11 11 03 03 03 03 03 03
 17 17 17 17 17 17 18 18 18 1c 1c 1c 32 32 32 67 67 67 84 84 84 73 73 73 77 77 77 7f 7f 7f 8c 8c 8c a9 a9 a9 ca ca ca e0 e0 e0 f1 f1 f1 fb fb fb fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe ef ef ef d3 d3 d3 bd bd bd b1 b1 b1 ae ae ae b0 b0 b0 ad ad ad a3 a3 a3 9b 9b 9b 94 94 94 7c 7c 7c 68 68 68 63 63 63 57 57 57 4f 4f 4f 55 55 55 46 46 46 17 17 17 05 05 05 03 03 03
 10 10 10 0e 0e 0e 11 11 11 17 17 17 27 27 27 61 61 61 79 79 79 6f 6f 6f 77 77 77 80 80 80 85 85 85 8d 8d 8d a6 a6 a6 ca ca ca e6 e6 e6 f5 f5 f5 fb fb fb fd fd fd fe fe fe fe fe fe fe fe fe fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe fe fe fe fe fe fe fe fe fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa fa fa e4 e4 e4 c6 c6 c6 b0 b0 b0 a3 a3 a3 9b 9b 9b 9b 9b 9b 99 99 99 92 92 92 8c 8c 8c 7d 7d 7d 69 69 69 69 69 69 60 60 60 51 51 51 4c 4c 4c 4f 4f 4f 48 48 48 20 20 20 06 06 06 03 03 03
 09 09 09 09 09 09 0c 0c 0c 12 12 12 23 23 23 55 55 55 6d 6d 6d 6b 6b 6b 76 76 76 81 81 81 81 81 81 85 85 85 8f 8f 8f a1 a1 a1 bc bc bc d6 d6 d6 e9 e9 e9 f1 f1 f1 fa fa fa fa fa fa fa fa fa fa fa fa fd fd fd fe fe fe ff ff ff ff ff ff ff ff ff fd fd fd eb eb eb cb cb cb cd cd cd ed ed ed fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe fe fe f2 f2 f2 d7 d7 d7 b8 b8 b8 a4 a4 a4 98 98 98 8e 8e 8e 87 87 87 81 81 81 7f 7f 7f 74 74 74 67 67 67 66 66 66 69 69 69 59 59 59 4f 4f 4f 4b 4b 4b 4f 4f 4f 4e 4e 4e 24 24 24 06 06 06 03 03 03
 04 04 04 05 05 05 07 07 07 0f 0f 0f 23 23 23 45 45 45 61 61 61 6c 6c 6c 72 72 72 80 80 80 80 80 80 7e 7e 7e 82 82 82 8a 8a 8a 94 94 94 a7 a7 a7 c0 c0 c0 d7 d7 d7 e6 e6 e6 f2 f2 f2 f4 f4 f4 f4 f4 f4 fa fa fa fe fe fe ff ff ff ff ff ff ff ff ff f2 f2 f2 a3 a3 a3 63 63 63 78 78 78 b3 b3 b3 eb eb eb fd fd fd ff ff ff ff ff ff ff ff ff ff ff ff fc fc fc e8 e8 e8 c7 c7 c7 a9 a9 a9 96 96 96 88 88 88 7d 7d 7d 74 74 74 6c 6c 6c 65 65 65 5d 5d 5d 5e 5e 5e 62 62 62 63 63 63 59 59 59 4e 4e 4e 4c 4c 4c 52 52 52 56 56 56 24 24 24 05 05 05 03 03 03
 03 03 03 04 04 04 08 08 08 10 10 10 2e 2e 2e 51 51 51 61 61 61 66 66 66 67 67 67 72 72 72 75 75 75 75 75 75 77 77 77 79 79 79 7f 7f 7f 8b 8b 8b 9d 9d 9d b9 b9 b9 d4 d4 d4 e8 e8 e8 f3 f3 f3 f2 f2 f2 f6 f6 f6 fc fc fc fe fe fe ff ff ff fe fe fe e9 e9 e9 7c 7c 7c 40 40 40 53 53 53 79 79 79 b7 b7 b7 ef ef ef fd fd fd ff ff ff ff ff ff fe fe fe f5 f5 f5 d7 d7 d7 b4 b4 b4 97 97 97 82 82 82 73 73 73 68 68 68 5d 5d 5d 52 52 52 4b 4b 4b 4f 4f 4f 55 55 55 59 59 59 5d 5d 5d 53 53 53 4d 4d 4d 4c 4c 4c 55 55 55 53 53 53 1c 1c 1c 03 03 03 03 03 03
 04 04 04 09 09 09 08 08 08 08 08 08 25 25 25 56 56 56 5b 5b 5b 5d 5d 5d 64 64 64 67 67 67 6e 6e 6e 6d 6d 6d 6c 6c 6c 6f 6f 6f 73 73 73 7b 7b 7b 89 89 89 a2 a2 a2 bb bb bb d4 d4 d4 ec ec ec f5 f5 f5 f7 f7 f7 fb fb fb fe fe fe ff ff ff ff ff ff e6 e6 e6 6b 6b 6b 30 30 30 42 42 42 56 56 56 7d 7d 7d b5 b5 b5 ef ef ef ff ff ff ff ff ff fb fb fb e7 e7 e7 c4 c4 c4 a7 a7 a7 89 89 89 73 73 73 64 64 64 4f 4f 4f 42 42 42 3d 3d 3d 40 40 40 46 46 46 4b 4b 4b 50 50 50 55 55 55 54 54 54 4f 4f 4f 4f 4f 4f 57 57 57 44 44 44 10 10 10 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 04 04 04 1a 1a 1a 52 52 52 61 61 61 63 63 63 5d 5d 5d 63 63 63 65 65 65 5e 5e 5e 61 61 61 64 64 64 67 67 67 6e 6e 6e 79 79 79 88 88 88 a1 a1 a1 b9 b9 b9 d0 d0 d0 e2 e2 e2 ef ef ef f8 f8 f8 fe fe fe ff ff ff fd fd fd e1 e1 e1 64 64 64 25 25 25 2f 2f 2f 3b 3b 3b 53 53 53 74 74 74 c4 c4 c4 fe fe fe fd fd fd f0 f0 f0 d0 d0 d0 b3 b3 b3 9e 9e 9e 86 86 86 64 64 64 46 46 46 37 37 37 33 33 33 35 35 35 3a 3a 3a 3f 3f 3f 45 45 45 47 47 47 4d 4d 4d 50 50 50 4f 4f 4f 50 50 50 4c 4c 4c 26 26 26 06 06 06 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 04 04 04 10 10 10 46 46 46 5d 5d 5d 5d 5d 5d 5f 5f 5f 63 63 63 61 61 61 5c 5c 5c 61 61 61 64 64 64 64 64 64 69 69 69 75 75 75 77 77 77 78 78 78 8d 8d 8d a6 a6 a6 b5 b5 b5 c2 c2 c2 d2 d2 d2 e5 e5 e5 f1 f1 f1 f4 f4 f4 e1 e1 e1 79 79 79 18 18 18 1d 1d 1d 27 27 27 38 38 38 4c 4c 4c 89 89 89 f4 f4 f4 eb eb eb d1 d1 d1 b9 b9 b9 a5 a5 a5 8b 8b 8b 68 68 68 4a 4a 4a 39 39 39 32 32 32 32 32 32 33 33 33 33 33 33 35 35 35 39 39 39 3f 3f 3f 47 47 47 4e 4e 4e 4e 4e 4e 4c 4c 4c 39 39 39 14 14 14 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 04 04 04 0c 0c 0c 2f 2f 2f 53 53 53 56 56 56 57 57 57 5c 5c 5c 59 59 59 57 57 57 56 56 56 5b 5b 5b 61 61 61 6c 6c 6c 75 75 75 73 73 73 6f 6f 6f 72 72 72 78 78 78 7d 7d 7d 7f 7f 7f 83 83 83 90 90 90 9a 9a 9a 9f 9f 9f 99 99 99 5e 5e 5e 12 12 12 13 13 13 16 16 16 23 23 23 33 33 33 5a 5a 5a c1 c1 c1 b4 b4 b4 9c 9c 9c 86 86 86 6f 6f 6f 5c 5c 5c 4b 4b 4b 41 41 41 3c 3c 3c 37 37 37 32 32 32 2f 2f 2f 2d 2d 2d 31 31 31 36 36 36 3d 3d 3d 44 44 44 4a 4a 4a 4d 4d 4d 4a 4a 4a 28 28 28 07 07 07 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 1b 1b 1b 3f 3f 3f 4f 4f 4f 4d 4d 4d 4f 4f 4f 4f 4f 4f 51 51 51 52 52 52 55 55 55 5a 5a 5a 5b 5b 5b 60 60 60 68 68 68 6b 6b 6b 6c 6c 6c 67 67 67 60 60 60 5d 5d 5d 5d 5d 5d 61 61 61 67 67 67 62 62 62 5b 5b 5b 39 39 39 0d 0d 0d 0d 0d 0d 0a 0a 0a 0f 0f 0f 1d 1d 1d 31 31 31 6a 6a 6a 68 68 68 61 61 61 58 58 58 4e 4e 4e 48 48 48 42 42 42 3b 3b 3b 35 35 35 31 31 31 30 30 30 2f 2f 2f 2d 2d 2d 2d 2d 2d 34 34 34 3a 3a 3a 43 43 43 4a 4a 4a 4d 4d 4d 3d 3d 3d 15 15 15 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 19 19 19 33 33 33 4a 4a 4a 4c 4c 4c 4a 4a 4a 49 49 49 4a 4a 4a 4a 4a 4a 4b 4b 4b 4a 4a 4a 4c 4c 4c 4f 4f 4f 53 53 53 57 57 57 5d 5d 5d 5b 5b 5b 55 55 55 52 52 52 51 51 51 57 57 57 53 53 53 4c 4c 4c 45 45 45 2c 2c 2c 0a 0a 0a 0a 0a 0a 06 06 06 05 05 05 0a 0a 0a 1c 1c 1c 45 45 45 4b 4b 4b 4f 4f 4f 4f 4f 4f 4a 4a 4a 45 45 45 3d 3d 3d 39 39 39 37 37 37 34 34 34 31 31 31 31 31 31 2f 2f 2f 2f 2f 2f 35 35 35 3d 3d 3d 4c 4c 4c 52 52 52 47 47 47 29 29 29 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 15 15 15 2c 2c 2c 43 43 43 49 49 49 47 47 47 44 44 44 47 47 47 4a 4a 4a 4b 4b 4b 49 49 49 48 48 48 4b 4b 4b 4d 4d 4d 4d 4d 4d 52 52 52 53 53 53 4f 4f 4f 4b 4b 4b 4a 4a 4a 4a 4a 4a 45 45 45 3e 3e 3e 38 38 38 26 26 26 08 08 08 07 07 07 05 05 05 04 04 04 04 04 04 0c 0c 0c 34 34 34 3d 3d 3d 45 45 45 4a 4a 4a 4d 4d 4d 48 48 48 3f 3f 3f 38 38 38 37 37 37 31 31 31 2f 2f 2f 31 31 31 31 31 31 30 30 30 37 37 37 4a 4a 4a 50 50 50 4b 4b 4b 3c 3c 3c 11 11 11 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0c 0c 0c 22 22 22 37 37 37 42 42 42 41 41 41 41 41 41 44 44 44 48 48 48 49 49 49 47 47 47 45 45 45 46 46 46 4c 4c 4c 4b 4b 4b 49 49 49 49 49 49 49 49 49 45 45 45 42 42 42 3a 3a 3a 33 33 33 2e 2e 2e 29 29 29 1b 1b 1b 05 05 05 04 04 04 03 03 03 03 03 03 03 03 03 05 05 05 28 28 28 37 37 37 40 40 40 47 47 47 48 48 48 44 44 44 41 41 41 39 39 39 37 37 37 31 31 31 2c 2c 2c 2b 2b 2b 2f 2f 2f 30 30 30 33 33 33 39 39 39 3c 3c 3c 39 39 39 1d 1d 1d 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 18 18 18 31 31 31 3c 3c 3c 41 41 41 42 42 42 45 45 45 46 46 46 44 44 44 42 42 42 44 44 44 43 43 43 46 46 46 4a 4a 4a 4a 4a 4a 4b 4b 4b 4b 4b 4b 42 42 42 39 39 39 30 30 30 29 29 29 25 25 25 25 25 25 1b 1b 1b 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 21 21 21 34 34 34 3e 3e 3e 43 43 43 43 43 43 44 44 44 41 41 41 34 34 34 32 32 32 2c 2c 2c 27 27 27 29 29 29 2d 2d 2d 2e 2e 2e 2e 2e 2e 2f 2f 2f 34 34 34 2a 2a 2a 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 07 07 07 25 25 25 38 38 38 3c 3c 3c 3e 3e 3e 3e 3e 3e 41 41 41 41 41 41 42 42 42 42 42 42 41 41 41 42 42 42 46 46 46 47 47 47 47 47 47 47 47 47 3a 3a 3a 31 31 31 2d 2d 2d 27 27 27 26 26 26 28 28 28 1e 1e 1e 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1c 1c 1c 33 33 33 3f 3f 3f 46 46 46 46 46 46 41 41 41 3c 3c 3c 31 31 31 2e 2e 2e 2d 2d 2d 2c 2c 2c 32 32 32 37 37 37 2f 2f 2f 30 30 30 32 32 32 33 33 33 14 14 14 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0f 0f 0f 2e 2e 2e 39 39 39 3a 3a 3a 3b 3b 3b 3d 3d 3d 3d 3d 3d 3d 3d 3d 3e 3e 3e 3f 3f 3f 40 40 40 41 41 41 40 40 40 3e 3e 3e 3e 3e 3e 37 37 37 30 30 30 2c 2c 2c 29 29 29 29 29 29 2a 2a 2a 1f 1f 1f 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 19 19 19 37 37 37 43 43 43 4a 4a 4a 47 47 47 3d 3d 3d 35 35 35 30 30 30 31 31 31 31 31 31 2f 2f 2f 2e 2e 2e 31 31 31 33 33 33 35 35 35 36 36 36 24 24 24 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 32 32 32 39 39 39 3a 3a 3a 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 3d 3e 3e 3e 3e 3e 3e 3f 3f 3f 3d 3d 3d 3a 3a 3a 38 38 38 32 32 32 2f 2f 2f 2d 2d 2d 28 28 28 29 29 29 25 25 25 1b 1b 1b 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 1d 1d 1d 3b 3b 3b 47 47 47 4c 4c 4c 42 42 42 39 39 39 36 36 36 34 34 34 33 33 33 33 33 33 33 33 33 33 33 33 35 35 35 36 36 36 38 38 38 2c 2c 2c 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 33 33 33 37 37 37 3a 3a 3a 3a 3a 3a 3a 3a 3a 3b 3b 3b 3c 3c 3c 3d 3d 3d 3c 3c 3c 3b 3b 3b 3a 3a 3a 37 37 37 32 32 32 2b 2b 2b 25 25 25 25 25 25 23 23 23 23 23 23 1b 1b 1b 07 07 07 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 38 38 38 42 42 42 43 43 43 3d 3d 3d 39 39 39 37 37 37 36 36 36 39 39 39 38 38 38 37 37 37 37 37 37 37 37 37 37 37 37 2c 2c 2c 0d 0d 0d 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 1e 1e 1e 34 34 34 37 37 37 38 38 38 38 38 38 38 38 38 3b 3b 3b 3c 3c 3c 3d 3d 3d 3d 3d 3d 3b 3b 3b 3a 3a 3a 36 36 36 31 31 31 2b 2b 2b 2a 2a 2a 27 27 27 25 25 25 1c 1c 1c 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 16 16 16 34 34 34 3b 3b 3b 3d 3d 3d 3e 3e 3e 3f 3f 3f 41 41 41 40 40 40 3e 3e 3e 3d 3d 3d 3a 3a 3a 3a 3a 3a 39 39 39 2f 2f 2f 11 11 11 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 24 24 24 35 35 35 38 38 38 38 38 38 38 38 38 3a 3a 3a 3b 3b 3b 3b 3b 3b 3c 3c 3c 3d 3d 3d 3b 3b 3b 39 39 39 36 36 36 33 33 33 32 32 32 2d 2d 2d 2a 2a 2a 1d 1d 1d 08 08 08 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 16 16 16 36 36 36 3c 3c 3c 40 40 40 43 43 43 43 43 43 41 41 41 41 41 41 41 41 41 3e 3e 3e 3c 3c 3c 3a 3a 3a 30 30 30 13 13 13 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0b 0b 0b 26 26 26 36 36 36 38 38 38 38 38 38 38 38 38 39 39 39 39 39 39 39 39 39 3c 3c 3c 3c 3c 3c 3a 3a 3a 39 39 39 38 38 38 38 38 38 33 33 33 2e 2e 2e 21 21 21 09 09 09 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 19 19 19 3b 3b 3b 3f 3f 3f 41 41 41 42 42 42 43 43 43 43 43 43 42 42 42 40 40 40 3d 3d 3d 3a 3a 3a 30 30 30 15 15 15 04 04 04 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 12 12 12 2f 2f 2f 39 39 39 3a 3a 3a 38 38 38 39 39 39 37 37 37 37 37 37 39 39 39 39 39 39 39 39 39 39 39 39 39 39 39 39 39 39 37 37 37 31 31 31 26 26 26 0b 0b 0b 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 3d 3d 3d 3e 3e 3e 40 40 40 42 42 42 42 42 42 45 45 45 45 45 45 3f 3f 3f 3a 3a 3a 2a 2a 2a 0d 0d 0d 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 19 19 19 38 38 38 39 39 39 37 37 37 39 39 39 37 37 37 38 38 38 38 38 38 39 39 39 3b 3b 3b 38 38 38 38 38 38 37 37 37 35 35 35 34 34 34 27 27 27 0c 0c 0c 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 18 18 18 42 42 42 48 48 48 52 52 52 5b 5b 5b 62 62 62 68 68 68 61 61 61 41 41 41 1c 1c 1c 08 08 08 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 17 17 17 2f 2f 2f 37 37 37 38 38 38 38 38 38 38 38 38 39 39 39 38 38 38 39 39 39 3a 3a 3a 37 37 37 37 37 37 36 36 36 33 33 33 29 29 29 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 23 23 23 6a 6a 6a 72 72 72 76 76 76 75 75 75 6e 6e 6e 5b 5b 5b 37 37 37 0e 0e 0e 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 0d 0d 0d 26 26 26 34 34 34 37 37 37 3a 3a 3a 40 40 40 43 43 43 46 46 46 48 48 48 47 47 47 46 46 46 46 46 46 45 45 45 3b 3b 3b 16 16 16 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 25 25 25 71 71 71 6d 6d 6d 68 68 68 5b 5b 5b 41 41 41 1d 1d 1d 06 06 06 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 06 06 06 16 16 16 2c 2c 2c 3d 3d 3d 53 53 53 61 61 61 6b 6b 6b 70 70 70 71 71 71 72 72 72 73 73 73 71 71 71 60 60 60 24 24 24 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 1b 1b 1b 5e 5e 5e 54 54 54 42 42 42 22 22 22 0a 0a 0a 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 09 09 09 19 19 19 33 33 33 4a 4a 4a 5a 5a 5a 63 63 63 67 67 67 68 68 68 69 69 69 68 68 68 58 58 58 21 21 21 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 10 10 10 34 34 34 1b 1b 1b 09 09 09 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 08 08 08 13 13 13 23 23 23 30 30 30 42 42 42 4e 4e 4e 52 52 52 51 51 51 46 46 46 1d 1d 1d 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 04 04 04 09 09 09 10 10 10 12 12 12 10 10 10 0c 0c 0c 05 05 05 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03 03
