 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 05 00 06 05 03 00 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 06 06 05 05 08 06 08 06 0b 06 05 03 00 06 05 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 03 06 05 03 00 06 05 03 02 06 05 04 00 08 05 06 03 06 05 03 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 03 07 05 0a 0d 07 08 04 09 0c 05 03 09 06 05 05 01 06 05 06 0b 06 05 03 05 06 05 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0e 06 05 03 04 06 05 06 04 06 05 05 0f 08 05 04 00 09 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 01 06 05 04 06 09 0d 11 11 0d 0f 0b 15 11 0e 07 0e 0d 0e 08 10 10 0a 19 12 0b 05 07 05 0d 0a 09 05 06 09 07 03 06 05 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0b 05 03 00 06 05 05 04 06 0a 04 06 06 0b 03 00 11 0b 0f 02 06 05 03 09 0d 0a 0c 14 11 10 04 01 06 05 06 03 06 05 03 00 06 05 03 02 06 0a 03 13 14 11 11 0e 0e 16 1d 23 26 25 24 33 29 25 20 1f 18 23 22 2b 27 26 15 20 22 1d 1b 1d 24 1c 11 16 0f 0d 0e 0b 10 0d 0e 0e 06 05 0b 01 06 05 03 07 06 05 03 03 06 06 0a 10 06 05 03 09 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0b 0b 05 12 09 0b 12 0e 17 13 11 11 0a 12 16 18 1d 24 30 39 34 32 14 11 16 0f 19 0b 0b 08 10 05 06 05 03 06 06 0b 14 17 2d 30 29 2c 2b 35 3d 48 44 47 4b 4b 4f 45 3e 31 30 3c 37 3d 37 39 37 38 39 40 36 39 35 2e 2b 2e 2d 25 1c 20 20 1f 1e 19 09 05 06 10 10 0a 0f 00 0c 0d 0a 02 10 05 11 0b 0c 0b 04 09 06 05 03 05 06 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 05 06 09 06 05 03 0a 09 05 09 05 0d 0b 0a 14 18 17 1c 1f 1c 1f 28 29 25 28 26 35 44 50 6d 6d 5a 3f 3d 34 2d 36 3a 35 2a 2e 24 11 06 05 04 17 1f 10 19 36 45 57 4f 51 57 53 68 66 74 70 62 63 50 4f 3a 45 39 39 34 38 3c 2e 3a 41 3a 3b 42 39 38 44 3a 36 2b 2b 33 32 36 37 30 32 2e 25 23 18 17 0c 0d 1b 21 22 1a 1a 19 11 19 1b 06 10 06 06 0d 08 07 05 06 05 03 03 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 07 01 06 05 07 0e 0e 0e 0c 0f 0f 14 12 1e 1e 20 20 29 2b 2c 36 39 36 43 47 4f 54 53 5b 72 77 8b 92 8c 6c 57 48 44 40 46 45 4e 4d 4e 43 32 11 11 14 2c 35 3b 3e 41 4d 4e 4f 59 5e 63 68 73 73 67 57 52 4f 42 3a 41 39 35 3a 3b 49 36 3c 3a 3c 3d 3c 47 3e 3d 3b 3f 42 3e 41 42 37 3d 43 4a 4d 6c 67 4a 41 38 2f 3a 37 36 2f 2a 25 25 1b 20 1c 1d 16 13 13 14 13 14 06 05 0c 11 09 08 0b 00 07 05 03 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 00 06 05 03 07 06 06 0a 0f 07 13 11 0c 10 14 12 0b 11 14 1d 23 1e 2e 33 35 31 42 35 46 53 51 64 60 67 6b 6c 77 7f 82 81 9e a5 a8 a2 86 6c 54 4e 50 4c 4e 49 55 55 54 52 42 33 28 34 3f 48 51 4a 47 4e 50 4c 50 56 53 57 5f 5e 5a 4e 4a 4c 40 49 43 3e 45 3b 3b 39 3d 3a 3a 43 43 41 3e 37 40 43 41 47 3f 41 3e 43 44 49 47 4c 69 8b 8e 79 66 5b 5c 59 4f 47 51 3e 3e 48 3a 42 3a 30 26 29 23 29 2a 1a 19 19 0f 11 1b 0c 07 09 05 0b 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0c 09 09 0a 0e 0e 11 14 12 20 1c 2b 2f 30 38 34 3b 42 40 46 44 4e 5d 6a 65 6e 7f 88 88 89 89 8b 97 91 9f a5 b0 b0 b8 ac 8d 78 63 54 51 49 56 4c 50 4f 48 4f 48 47 45 54 50 4b 4b 4d 52 58 53 5a 56 50 53 51 53 4d 4e 4d 4b 48 51 4a 3e 46 3c 44 32 44 43 39 39 3f 3f 43 3b 41 42 47 47 45 49 41 3e 42 42 51 4d 54 57 60 7c 9b ac 9b 8a 84 81 83 72 70 6e 60 6a 6b 6b 6d 61 59 4c 50 44 3e 32 2d 28 26 23 2c 1c 1a 11 05 07 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 04 06 06 0a 03 06 0e 11 20 1a 14 1f 1f 27 35 32 3a 4a 4b 5a 56 5e 65 6c 69 6b 75 7a 85 88 9b 9f a5 ae b5 b5 aa af ad ae b8 ba b7 ba a7 9f 89 74 78 69 59 55 59 56 54 54 4f 48 4d 4d 56 4d 50 52 52 59 5e 5a 5d 67 62 5e 5a 51 57 53 52 59 4a 4d 47 4d 4f 49 46 41 46 3e 44 41 43 45 45 49 45 41 45 4a 47 44 48 49 48 45 46 44 49 4c 52 51 5c 63 79 a0 b2 bb b9 b4 a9 a1 98 97 95 91 91 95 94 89 76 6a 62 66 60 51 4a 50 4d 45 3b 44 38 29 2c 1a 14 16 0f 13 11 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0b 0b 05 12 0a 0f 22 22 25 33 42 41 44 57 5e 72 80 88 8b 86 90 94 9a a1 a0 9b a5 ab b5 be c7 c3 c1 cf bf b7 b5 b4 ae aa ab a7 9e 96 7f 78 72 6c 63 67 62 59 5f 59 59 59 55 54 53 52 58 5b 5e 59 62 5d 58 60 60 67 67 60 5e 63 5a 53 52 5f 56 47 56 4f 54 4b 52 4d 44 45 49 44 41 43 4e 45 4b 50 48 44 4f 50 47 46 47 45 4c 3f 4e 4b 54 5d 5e 64 6c 75 89 a4 ba cd c4 c1 bd b7 b5 b1 b0 a7 a5 83 6f 5b 5e 59 60 5d 54 57 58 5d 6e 60 4f 41 35 32 20 26 29 27 20 1c 0d 09 07 06 05 06 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0b 06 07 12 03 0e 0c 17 20 26 30 44 4d 5e 6a 6c 79 85 9b a4 b5 c7 c9 ce d4 d2 cb d2 d0 cd d3 d5 d0 d5 c9 b6 af a5 98 97 90 91 86 83 85 7b 7a 6f 6f 69 6a 64 64 6e 5e 5f 66 66 60 56 60 4f 63 5c 5b 59 63 5d 5f 62 5a 5d 66 61 66 5f 60 5c 4f 57 53 51 59 4f 59 53 5e 51 54 4d 4f 46 48 4b 42 46 4a 48 4d 45 4c 42 44 4b 43 4b 46 46 4f 4c 53 52 50 57 5d 5c 66 5e 70 7a 89 a5 ad b7 be bc b8 ad 94 93 7d 69 5f 63 5a 61 5e 5b 5f 59 68 72 8c 7c 70 5b 4e 44 36 31 3b 36 2f 27 1b 0c 0b 06 0c 09 05 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 00 06 05 11 10 15 0b 17 1d 2b 35 42 47 45 58 5e 71 7d 81 85 85 8e 97 a1 af c0 c4 d5 d8 e9 df d2 d3 cb c9 c0 ab a2 99 90 92 8e 84 85 86 80 78 6e 74 71 73 6b 64 6c 60 62 66 6c 66 60 61 65 62 61 65 65 66 65 64 66 62 61 64 64 5e 65 66 62 67 5d 5a 62 5b 5d 5e 66 57 5a 5d 58 52 50 51 53 55 48 4e 50 43 43 4c 4d 50 52 4c 53 4d 4e 54 43 49 4a 4b 51 4e 5b 55 50 5e 64 62 67 67 6e 72 7b 81 80 89 94 83 88 79 6e 69 59 5d 61 62 62 5d 66 65 68 72 75 90 a0 87 7d 7a 61 51 47 53 5d 4a 32 24 12 19 0a 13 0f 0d 10 0c 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 09 05 08 11 0d 15 10 15 1a 25 37 3e 4e 58 58 58 5e 63 63 73 73 7f 85 7b 82 88 88 92 90 9b a9 ac b1 ad ae a8 a3 98 a3 a0 9a 96 91 8c 86 82 7a 74 7b 75 73 70 6e 69 65 67 68 66 68 6f 72 69 69 66 6d 6b 68 73 6b 6b 6c 69 70 6b 71 72 6f 71 6b 6c 69 68 5f 62 62 64 5e 63 66 5d 56 62 5c 5f 5d 58 57 5f 52 5a 4f 50 4e 58 53 54 52 4f 51 53 51 4b 4d 54 50 53 4d 56 4b 55 5a 5d 61 65 6b 69 6b 74 75 6b 67 62 6b 74 72 67 66 64 60 60 60 6d 62 64 65 70 69 65 6e 80 91 95 8f 82 64 58 5d 6b 80 6d 52 39 29 22 22 24 19 21 13 0d 05 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 02 06 05 03 0b 06 10 12 0b 1d 16 1c 2e 3c 3e 47 50 5d 62 63 59 6a 65 74 75 75 71 80 82 87 84 87 98 8c 9c 94 99 9e 9c 92 93 8e 96 9c 94 93 8c 84 86 83 7a 71 71 7b 6d 71 6f 6f 70 62 5f 72 63 6d 6c 6a 6a 6d 71 6e 6b 6b 71 6f 73 6c 74 6f 78 6e 6a 73 7a 6b 73 64 6b 67 61 65 67 60 66 65 64 5f 5f 58 61 63 60 54 5e 57 54 58 56 50 58 52 50 50 52 51 52 55 4a 46 4e 51 4e 4d 4b 4c 53 5c 62 5e 60 6e 68 62 6b 6e 68 68 69 5e 69 65 61 64 69 65 60 6b 65 64 6f 67 67 64 62 5d 6b 72 77 76 71 5b 5c 66 7e 9f 89 70 52 46 3f 30 36 2f 2d 24 15 0c 0c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0d 0a 05 0e 09 16 1a 1f 23 2f 40 47 47 56 56 64 67 5f 64 64 65 6e 70 76 7f 79 7d 80 85 8d 92 8d 8b 8a 98 90 91 a1 99 8c 8d 91 90 82 8d 8b 85 8f 85 79 74 75 71 66 67 6f 6d 70 66 68 69 67 6d 6f 70 78 76 79 6e 77 76 76 77 74 77 7c 78 72 78 7b 78 77 73 78 6e 6f 6c 6b 66 6b 68 6b 6b 65 5b 63 63 66 5b 61 63 62 62 5d 57 51 55 50 52 59 5c 54 51 58 51 51 55 50 4c 4a 50 4e 52 50 55 5e 69 65 6a 6c 66 63 68 69 6b 5f 60 67 6a 62 66 68 68 61 69 67 6a 68 66 64 63 61 64 64 63 64 66 63 5c 5d 60 76 9c a0 8d 74 63 54 49 5b 4d 44 29 1c 14 1c 12 0d 04 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 06 05 06 05 0a 07 0d 10 0c 17 18 1d 2f 33 48 54 51 52 5f 64 63 64 70 64 69 67 6f 71 78 75 7d 7d 7e 81 88 8e 8b 8f 8e 93 95 90 8f 9a 95 8e 8f 94 95 91 92 90 8d 89 8a 83 77 78 7a 7d 74 70 6d 67 6b 67 6c 68 73 71 74 75 6f 7c 7d 77 80 7c 83 84 77 84 79 7c 78 79 80 7c 7a 77 7a 6d 6a 7a 76 70 6a 62 69 66 64 63 69 65 60 65 6a 63 62 62 5f 5c 60 5f 59 60 55 53 59 5d 5f 55 54 54 4c 4f 4e 56 57 5c 59 5c 6c 66 65 69 6e 6e 6f 60 67 62 67 6a 6a 6e 6b 6b 61 68 6a 67 67 6f 70 6e 69 62 64 60 66 60 62 61 5a 62 5f 6c 83 a1 a7 99 88 8a 7b 7b 5f 55 44 2d 21 25 23 19 11 04 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 09 04 09 0a 0b 0a 17 1b 1e 2a 34 41 43 5e 5c 65 5d 5d 63 65 67 6f 71 6a 74 6b 6c 6c 73 6e 7d 7d 7d 7b 82 86 89 91 8b 98 99 97 96 a2 8e 95 91 92 9a 91 93 96 8c 90 85 7f 77 6f 76 73 76 75 74 74 6b 6b 68 70 68 73 7c 7d 7d 7f 85 82 7d 7b 85 84 7e 85 83 82 7a 83 79 7e 78 80 78 73 72 78 72 75 70 75 6d 6e 6a 65 62 6f 6d 66 60 6a 60 60 6a 5b 5a 61 65 63 5e 5e 5d 5e 60 54 52 4e 4d 4f 50 4f 54 5a 57 60 5d 66 6a 70 6f 6c 6a 69 66 66 6b 68 68 6a 6f 71 68 6f 6e 69 71 69 6d 6b 70 62 64 62 66 61 65 63 62 67 66 66 6f 87 a7 b4 a5 af a0 9a 7e 6c 5a 4b 33 41 3a 2c 1e 19 0c 08 03 01 0c 14 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 09 0e 16 16 1d 15 18 17 1e 27 40 51 58 75 6f 5a 5f 5a 60 62 68 6c 6e 6e 70 6a 71 6a 72 71 73 7b 79 78 78 78 77 82 86 90 90 94 99 9d 97 95 84 81 98 96 93 9c 94 91 93 8c 85 76 7e 7a 76 78 71 7a 76 6f 69 6f 71 6c 74 6e 82 81 7c 79 86 7c 84 88 86 87 8f 8e 8a 8c 80 86 84 87 84 81 7b 7d 79 78 7c 74 71 6f 6c 6f 69 6d 73 71 72 6c 6e 6a 68 66 6a 61 6a 64 58 5d 54 63 5a 55 60 5f 57 57 57 54 4d 54 52 58 60 59 63 5e 66 68 6c 6d 66 6e 64 67 67 6d 77 68 6f 74 6a 72 78 74 6f 6f 6e 6e 6c 6b 66 6c 63 67 6e 68 62 69 5b 64 69 6f 85 99 b0 bb bb ae a6 8e 70 65 59 5f 54 4c 33 1e 0b 07 09 04 08 16 17 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 02 16 25 23 23 25 26 2e 3e 47 55 62 75 7e 94 8b 6b 5a 64 5e 63 67 66 6c 6d 6d 6c 69 6e 70 77 70 70 7a 7b 83 7b 83 86 86 8c 9a 9a a0 a3 a2 a7 9f 9f 9a a1 a1 a0 9d a2 8c 8b 85 87 77 79 74 7a 70 74 71 64 76 6b 6e 76 72 77 82 81 84 85 85 87 8b 8f 89 88 97 85 8e 8a 8d 87 82 87 86 81 83 86 7e 7e 74 7c 77 7b 73 71 72 6a 79 6b 75 7b 74 6e 72 71 6c 6e 65 6a 5d 65 5f 66 63 5c 65 62 54 61 5a 5f 59 5b 53 56 5b 5b 62 6f 65 65 6e 69 6d 71 6e 6a 6c 6f 6a 79 71 6e 78 7f 7c 6d 71 71 76 6c 60 65 63 70 60 64 68 6d 69 6a 6a 69 69 67 69 74 80 9d bb c6 c3 af 96 87 72 69 67 65 50 30 1e 07 0e 06 06 05 17 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 09 00 06 16 0c 15 1d 1e
 2f 2c 32 40 56 61 71 80 91 9b 9d 95 7c 65 5f 64 65 63 70 76 63 70 6c 6b 71 6e 6e 76 74 78 7b 77 80 80 84 84 84 92 95 99 a1 9d a7 ad a3 a1 a3 99 a8 a2 9d 9a 9d 94 87 7d 78 7f 7e 7e 74 77 6c 74 6a 6f 77 6b 77 72 80 8c 87 87 91 8a 8e 8c 8f 90 98 9a 90 8b 8b 8d 91 85 8a 87 81 87 81 7e 82 7e 7c 7e 75 79 72 75 74 75 6d 75 72 74 6c 72 6d 75 70 6c 6f 72 67 64 68 61 64 64 59 5d 5c 5a 58 58 53 5d 5c 65 63 62 6c 6e 68 70 6d 6e 67 6f 72 79 7e 70 81 7f 7f 7f 84 7d 76 70 6b 70 6b 6b 66 74 6e 6e 6f 70 68 6b 72 6c 6a 69 69 6e 7c 7a 89 9c ab a6 98 89 72 70 68 73 6c 4b 30 1f 10 09 0e 13 16 11 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0c 0f 17 27 25 2b 36 48 55 68 7b 7d 95 a8 b8 a8 95 75 6b 63 5b 63 6b 67 65 72 73 67 72 71 6e 70 73 6f 78 7d 77 76 7e 80 7b 86 86 90 93 93 a4 98 aa ad af a9 a3 af 9e a1 a5 9e 97 91 8b 84 72 80 79 7b 75 72 71 72 73 6d 75 74 79 79 81 8a 78 90 8d 94 93 8d 94 8f 96 9a 94 91 8e 90 93 8f 8b 92 88 83 81 86 7e 81 7b 78 72 79 72 75 76 76 78 79 7c 7a 6c 70 72 6c 70 6a 6e 71 69 6d 6b 63 60 63 62 56 5c 53 53 52 60 5d 60 5b 64 68 64 68 6a 6f 6a 72 75 75 71 7b 77 7d 82 83 7b 82 81 78 7a 71 70 70 6c 6c 6f 66 71 71 6d 6f 6c 6b 67 6c 6f 71 6a 6b 75 7c 7e 78 7c 86 80 70 71 79 69 74 6f 51 35 32 1c 14 11 0b 15 11 09 07 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 09 0e 15 13 16 2b 27 32 3a 3b 57 71 7e 86 98 b4 bb c1 b2 86 74 65 69 6d 69 63 66 6a 72 69 6e 71 73 72 6c 6b 6e 76 70 78 7e 7e 7d 87 81 83 83 8c 8e 97 9d a4 a8 ab a6 b0 b0 af b2 a8 a3 a1 99 99 8e 86 86 7d 7e 79 74 74 76 77 7d 79 70 75 80 7c 81 8b 88 8e 90 8b 98 9c 8e 95 98 98 98 94 93 94 8d 92 90 87 87 91 87 89 85 79 80 7b 81 7c 73 77 7a 79 79 6d 76 78 77 7b 7e 6d 7b 70 69 64 6a 68 6b 64 64 6a 60 64 59 5f 56 55 52 5c 62 60 65 65 6d 70 6b 6e 6e 78 73 77 76 76 86 88 87 83 81 82 88 8a 81 71 6e 6a 72 6c 75 78 71 75 7a 7b 72 73 70 73 6d 72 71 74 72 75 6e 7d 77 82 76 80 6e 76 71 6f 6b 4f 42 47 40 30 1a 18 14 0e 08 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 09 05 09 0d 0a 17 1f 25 39 3b 41 5d 6b
 74 89 9c b3 c4 c1 b3 91 7f 75 69 6e 6a 78 5e 6a 71 71 76 74 78 79 73 79 7f 71 6f 7c 7a 80 7b 86 87 81 85 85 87 8f 97 8f a2 a5 ad b5 b7 b6 b4 aa af a5 ac 9c a5 99 97 8d 8b 83 83 81 79 7f 7c 75 76 70 79 7a 84 7c 80 83 85 8c 92 95 94 99 96 96 93 9d 95 97 90 94 92 95 97 8d 8d 87 88 8e 85 84 82 79 7c 7f 77 79 7e 7c 7a 86 7b 79 70 77 74 71 73 76 75 75 6f 6a 71 6b 6d 6a 64 62 61 5b 55 62 61 55 5c 5a 63 64 6a 6d 72 71 7c 75 7c 85 7f 87 89 88 87 86 8f 89 85 8d 83 77 7a 79 78 77 7a 7f 7e 81 79 79 77 77 77 78 73 73 76 70 76 74 7b 78 78 72 7c 78 7e 77 77 64 6a 50 4a 4f 52 4a 3e 25 1d 0d 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 08 06 09 09 12 11 1c 21 35 4d 52 6c 7a 84 97 ab c1 d6 d0 9d 8a 71 6d 71 73 65 6e 70 75 69 73 73 6b 70 76 80 80 7e 78 79 77 77 75 79 7b 88 87 79 84 81 8f 88 89 99 a3 9e aa b3 b4 b5 b7 b5 b5 b5 ad a4 a3 9d 8d 84 8f 81 7f 83 75 7c 74 75 7d 76 77 79 7b 7a 85 87 88 8b 8b 8a 92 8f 92 97 97 9b 98 9c 96 94 92 93 94 90 93 8b 8d 89 85 84 87 7f 7d 84 7e 7c 85 7d 84 7f 77 7d 75 7b 77 6e 76 7e 7b 75 72 74 72 69 6d 62 6a 68 64 65 60 64 5b 59 60 62 6c 65 6b 70 76 79 7e 77 79 78 85 8c 90 87 93 8a 8b 83 92 81 81 7a 72 79 70 6f 79 7f 83 7f 8a 7b 7d 7b 7a 80 7f 7b 7b 74 75 71 7b 76 7b 74 76 80 7b 7a 70 6f 60 4b 4a 5d 5e 4f 4e 40 2b 25 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 01 06 10 11 16 1f 27 2f 3e 50 75 85 8a a0 a1 b4 c9 dc d6 9d 7b 71 74 72 7e 74 70 70 70 71 73 75 72 7b 79 7b 7e 86 7f 83 7a 79 74 7f 79 83 8b 92 8a 87 8e 8c 86 8a 9c a0 ae b2 bb b7 b5 b7 ba b4 b1 ac a5 a6 a4 97 90 8f 85 8b 84 86 82 78 73 7c 71 74 76 7d 78 82 86 85 8a 82 8a 8c 98 8e 96 94 94 8d 93 92 92 95 8f 8e 8e 8f 84 86 84 85 8f 87 83 81 7c 7b 7d 7f 84 82 82 7d 8a 80 7b 74 7e 7a 7b 7b 7a 62 72 6d 73 75 69 6e 70 67 69 60 5d 64 66 64 60 66 66 6b 72 7d 7c 78 8e 85 81 90 91 92 89 94 8d 89 87 8d 82 7f 7b 7d 82 7d 7c 7e 86 7e 80 80 85 80 86 81 7a 7f 7c 75 7e 76 7a 76 7a 7d 7a 7c 83 79 7b 76 6e 5f 58 4b 6a 6c 5f 5a 56 4d 30 26 17 0a 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0d 11 0c 10 0a 15 12 1f 33 3c 4a 61 72 8f a1 ac b3 be
 c9 ce cf b2 80 76 78 76 73 76 6c 7b 77 71 7e 72 77 7a 7e 7f 83 8a 81 88 89 7f 7c 7b 83 7e 8b 93 89 94 90 9b 92 8f 99 9b aa aa b3 ba bb bb bc bc b9 b4 af ad ae a3 92 93 94 8a 84 84 83 7e 79 78 7b 7b 7c 7c 77 74 7f 87 84 8f 8b 8e 8f 8d 97 90 8c 98 94 94 95 8f 98 8b 96 97 90 8e 8f 86 92 88 88 88 84 87 7a 84 7f 84 88 82 7a 80 7a 81 82 7c 74 77 76 7a 7a 72 79 74 71 70 75 6a 71 62 61 6d 61 61 66 65 70 76 75 75 76 81 8a 89 91 8f 95 98 a1 96 97 9c 93 95 95 90 8e 78 83 8b 84 8b 8d 87 8c 8c 88 87 8d 89 85 8c 7f 82 78 74 74 82 76 7c 7f 81 81 81 72 82 7a 78 6e 5f 5d 5b 62 5f 67 71 65 4f 36 1e 1a 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0d 0b 0b 0c 16 1b 20 2f 4d 57 65 79 8d 9a 8c 9a 9c a4 b8 b8 a8 8e 74 73 75 78 73 78 75 77 71 73 70 78 81 76 7d 82 83 8b 84 84 88 89 85 81 7d 84 88 93 90 98 92 92 95 92 93 a3 a4 a7 b8 b5 ba c4 bd bf b9 b2 aa ae 9d 9f a1 98 94 90 8c 8d 80 85 7a 81 7c 6f 74 72 79 79 87 84 87 8b 8c 8f 8e 8b 92 8f 98 93 90 8e 8a 95 96 8f 8f 8f 8f 91 8d 90 86 91 84 87 8a 85 84 84 83 89 7e 80 81 83 7d 7d 7d 7c 7c 7f 81 80 7d 79 7a 78 79 6c 77 75 69 6d 69 68 62 69 6f 6d 77 73 7b 80 7d 8e 8a 88 93 97 95 95 9a 9c 9e a0 99 98 9a 92 92 7f 85 7e 84 8f 8f 92 8f 8c 90 89 83 8f 87 8a 7f 80 82 80 78 76 85 80 79 7c 76 78 7e 77 7c 7b 71 63 64 58 5b 65 72 7e 78 5b 37 27 15 10 11 07 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 00 09 06 03 02 0b 0c 11 1d 23 28 3d 54 66 7a 7a 92 8a 7e 70 70 78 83 8d 89 86 82 79 6f 7b 74 72 79 7a 75 77 7a 79 7c 81 7c 84 81 86 8c 8d 89 92 86 8d 85 8c 83 8f 95 91 99 97 a0 93 95 9f a5 aa b0 b4 bd bd bd c6 ba bc b5 b9 ab ab a4 a6 96 97 96 96 95 89 80 89 85 74 70 7d 77 7a 7f 7f 82 80 82 85 89 85 8d 8a 8c 87 8f 95 82 8c 8f 8a 8d 8b 91 86 92 84 8e 92 83 91 88 88 8e 81 80 90 7f 85 82 82 83 83 82 7e 86 81 7b 82 84 80 7f 7e 7b 77 75 78 76 74 76 6e 68 65 65 6a 68 70 77 7b 81 80 89 91 99 98 9a 9c a4 a5 a0 9e a7 8f 9b 97 96 94 91 86 8c 92 96 8f 96 94 8c 92 91 87 8f 90 8c 82 81 81 84 7a 7e 7a 78 82 78 7e 77 81 80 7e 7d 6b 65 62 5b 59 64 69 8b 94 75 4e 39 1c 1e 12 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 06 03 10 0a 1f 1a 24 36 41 55 70 80 97 9b 8e 66 74 73 6c 76 79
 6c 77 82 7a 7a 75 78 68 73 84 7d 7b 7f 78 7e 7d 85 8c 85 8d 86 8d 9d 98 8d 8a 8a 8d 8f 8e 96 94 a3 9c 9a 9d 9f a0 a6 9f b2 b2 ae bd b7 c6 c0 c0 b9 b9 b4 b0 ac a5 a6 a2 a0 9f 96 93 8e 92 7e 7e 7e 81 7d 7c 7f 7d 87 83 81 86 87 84 8d 84 86 8c 8b 8f 88 8a 8c 8f 8f 95 8d 95 91 8a 88 89 88 8d 89 88 90 8e 7f 83 89 83 7e 87 84 84 7d 7e 7e 81 7b 88 7b 84 88 7f 7c 7a 83 7b 7a 76 6a 71 6e 76 69 74 75 70 7b 80 85 87 8e 8d 92 97 a0 a1 a0 a2 a7 a2 99 a2 a1 9e 98 99 94 95 93 91 9a 98 99 9a 8f 93 9b 95 8f 92 93 84 8b 81 7f 78 7a 7f 80 7f 7e 7c 76 7c 7d 78 7a 73 64 63 60 5f 5c 64 6d 8c 9e 83 57 3c 30 1f 1c 0b 09 08 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 05 07 07 09 0d 14 1c 1e 33 3b 4e 6a 72 8a 95 a8 91 74 61 60 5e 69 6f 69 73 73 72 75 74 75 72 74 79 73 75 7e 80 80 81 7f 83 83 8e 8b 91 9f 93 96 9b 90 93 8e 92 8d 94 96 99 a0 9f a2 a5 ad a9 b5 b0 aa b7 bb bb bd b1 bd b7 b8 af b0 a7 a7 a1 9a a0 9f 93 95 92 8f 91 85 7e 86 76 7b 7d 74 80 80 86 7e 85 81 85 8d 8b 8c 85 87 8b 8c 8b 8b 8b 8a 85 92 8d 8e 90 90 8b 84 8a 8e 91 86 84 89 85 86 8a 84 84 7d 80 84 86 84 87 86 85 84 8a 84 8c 8a 81 7c 7f 7e 70 76 71 76 73 7b 79 7a 82 7f 84 8b 97 95 9c a5 a8 a2 a5 9f af a4 a1 a2 9e 9f a3 9a 9c 96 98 97 94 9b a3 9a 9a 9a 9b 9c 8f 90 8e 8e 88 84 89 7f 7d 7a 7e 7f 7c 7a 7e 75 7f 78 7d 75 70 65 60 59 61 67 6d 87 a8 91 6e 4f 36 20 19 1b 14 0d 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 05 08 0e 16 0f 14 23 25 34 47 5f 73 84 95 98 a2 96 7a 65 5d 65 62 67 73 6e 75 72 7a 6f 71 7a 76 70 6c 85 77 7a 7f 79 79 85 89 86 90 8f 93 9a a2 97 98 91 8a 8f 95 92 94 a2 9c a3 ae a7 b3 a8 aa ae b3 b5 ba be b8 b6 b6 b3 b3 b9 ab b1 a5 a3 a2 99 91 9f 99 9b 96 8f 8f 84 8a 82 83 7d 7a 78 85 7f 86 86 83 8a 84 8a 85 88 8e 91 87 85 89 8f 88 92 92 8e 97 90 94 90 91 9a 8b 8c 83 90 87 87 88 85 8c 84 81 89 80 89 88 83 7c 8a 88 8b 88 89 85 8e 87 82 82 7a 7b 7e 75 78 75 77 7e 75 7f 8e 8a 8f 91 99 a1 9e a4 ad ab b0 b0 ab a6 a3 a1 a5 a7 9f 9a 9a 96 a2 95 99 a0 9f a3 9a a6 a2 8b 93 89 92 8d 80 81 86 7d 79 82 80 80 80 79 79 7d 79 71 75 6d 6e 6e 68 65 6c 74 81 b4 a1 80 5e 3d 34 29 23 19 0e 07 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 10 12 18 18 20 22 38 42 54 5e 80 8f 94 92 85 7f 71 63 69 69 65 65 6b 66 6b
 77 6f 75 7a 73 78 74 70 77 74 79 7c 7b 87 87 83 90 85 89 9a 98 9b 9f a2 96 9d 97 a1 a0 98 9d a0 a3 ad b3 b0 97 ad b1 ae be b7 b7 c0 c1 b6 bf be bb b4 b0 a8 a3 a1 a4 a1 9e 9b a7 9d 97 9a 91 93 85 87 83 84 78 7d 7e 87 82 82 89 83 89 8f 8b 86 8e 8c 8b 8d 8f 8d 97 98 94 9c 9f 9a a2 9a 9d 9d 96 95 8e 86 83 8f 85 8d 81 87 86 88 8c 8a 8d 87 8b 8f 8b 8b 89 8b 90 84 81 85 91 8b 7f 86 71 76 83 82 7f 84 8f 8e 8d 97 9a a6 a5 aa aa ac b4 a9 aa ac a4 a5 a9 a1 a1 a5 ac a6 9d a5 9f a4 a9 af a7 a1 9b a3 98 97 95 8a 8a 84 8e 8f 8b 93 7d 82 7d 82 79 80 7d 77 7e 7d 7c 70 75 6a 71 78 73 84 ad b6 92 72 55 3a 2a 28 27 1b 11 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 0e 0b 17 1d 1c 25 34 43 4d 4f 51 5e 67 6f 68 67 65 61 66 67 62 60 67 69 6e 6b 74 73 72 71 75 7b 70 73 79 7b 7f 79 7e 7b 80 7f 85 8a 8a 8c 9b 95 a1 96 96 9a 9d a1 9a 98 a1 a0 99 a2 a1 a5 ac ae b6 b4 ad b5 b1 ba b8 be bc b5 ba b0 ae b5 a5 aa 9d 9a a5 a4 a0 a8 a1 98 9c 96 8e 95 94 8c 83 7e 7d 88 84 87 86 8b 8a 87 8f 8f 8b 96 94 8d 9a 96 93 9a 9a 9f 9f 9b ad a8 a9 a8 9f a0 9c 92 85 83 8d 85 89 8f 8b 81 8c 85 85 8c 8d 8c 96 8c 94 8b 8d 97 8b 9a 89 8e 8b 85 82 7b 84 83 8c 8c 88 8a 8f 95 a1 a4 a8 b0 b5 ab b3 b1 aa af a9 a9 a5 a9 a2 a7 a7 aa aa ab a0 a7 a8 a6 a8 a3 a2 a5 9d 97 91 93 8f 8e 8d 8b 8c 85 85 76 85 78 7d 79 80 7e 7a 79 82 77 72 7a 74 74 72 79 87 ab c4 a5 86 61 4b 37 38 2f 1f 17 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 18 1b 1c 1b 2a 3c 47 4a 56 51 54 5a 5b 60 58 57 5b 60 60 67 64 62 61 60 6b 6e 6f 75 6f 6e 73 72 70 77 78 76 75 70 7b 7a 7f 85 87 88 90 92 90 92 9b 9c 9b a2 a1 a2 99 9d 9f a2 9c a5 a5 a1 b1 ab a9 b4 b4 ba ae bb b5 bd b5 b4 b2 b5 ab b5 a7 a1 a1 a5 a4 a5 a7 9d a5 a3 9f 99 9c 95 8e 92 8c 8a 7e 84 84 8a 85 89 84 97 98 94 96 90 95 94 94 9d 9f 99 9f a5 a0 a4 a2 a5 ab aa 9e 9f 9e 95 92 85 8d 85 88 8b 8c 91 8f 91 95 88 93 87 95 96 9c 95 99 90 92 97 8f 90 91 8c 8d 88 88 87 87 84 8c 90 9e 9d a2 a1 ae aa b3 bb ac b1 af a9 a7 ad a7 a7 a6 a8 ad a1 ab ae a8 a7 ae aa b0 ae a1 a4 9e 9d 99 96 91 8a 94 8e 85 83 7d 7f 84 7c 82 75 71 7d 73 80 7c 83 74 71 6e 70 74 7c 7c 9b b9 af 95 69 55 51 3c 35 28 25 11 10 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 07 0b 1d 17 24 27 3b 47 52 51 57 54 59 56 5e 5f 5c 54 5d 5c 63 60 5c 63 66 60 66 69 72 68
 6e 76 77 76 7a 7d 77 7a 79 7e 78 7c 7f 84 86 84 87 82 8c 92 8e 94 93 9b 9c 9e 9f a6 a3 a3 a3 a3 ab a9 a5 a8 a4 a7 b6 b7 b4 b5 b4 b8 b9 b9 b8 bb b5 aa b1 a5 a0 a2 a8 a0 a3 a7 a2 ac a8 a0 9d 93 97 91 91 8e 8b 8d 8d 91 8b 8a 8d 95 9b 98 92 98 93 98 a1 95 9c 99 96 a0 a0 a4 a7 a3 a3 a3 aa a7 a7 a2 9c 88 85 88 87 8b 8e 92 8b 95 92 95 93 91 99 9a 98 9e 99 9d 97 96 9b 99 98 a2 9d 9e 95 95 8f 99 90 95 9d a0 a6 a5 a9 b1 b1 ae bb b5 b6 b1 b1 ad b1 ab ac ae ab af b4 b0 b3 b2 ac ad ac ad ab a4 a5 a8 99 9d 96 9a 8a 91 8f 84 81 80 83 7e 78 7c 6b 74 76 77 76 7b 75 6f 7a 75 79 75 76 75 92 bc c9 af 93 78 5e 50 40 30 1d 19 0e 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 19 13 22 29 28 37 52 62 59 57 55 58 58 5e 54 58 5a 64 59 5f 60 66 68 66 67 68 6b 6c 71 6f 72 79 75 7b 7d 7b 7b 79 79 7f 76 72 7e 82 84 7f 7b 87 8d 90 98 95 97 9c aa 9f a6 a6 a2 a3 9d a7 af a9 ab a9 ad b0 b0 ac b1 ac b0 ba b7 bb ae b4 ae ab a7 a5 a8 9e a5 a5 a3 a4 a8 a6 a5 a5 a2 a1 9c 92 92 8d 8b 8f 8e 86 93 90 8f 92 91 9a 95 9b 94 9c 96 95 98 96 96 96 93 9f 9e a1 a0 a0 a6 a0 97 9c 97 8d 8b 8e 88 8d 93 94 8a 9d 9a 92 9d 93 9d 9f 9e 9a 9b 9c 9e a3 a1 9f 9b a0 96 9c a4 94 9d 9e 95 a1 a4 9d a0 a8 b1 af bc b4 b3 aa b3 b8 b3 af a8 af b5 ae b5 b2 bc bd b7 bb b7 b1 b3 b5 ae ad ab a2 98 9f 96 97 98 8f 8b 80 7f 83 88 87 7d 79 74 7e 77 72 79 77 78 7a 7d 75 7a 75 78 79 89 b3 c7 b5 9e 85 71 66 54 44 34 24 15 16 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 08 12 11 16 24 29 3a 48 68 72 62 5e 52 55 5b 5b 5b 66 60 56 66 64 63 65 62 6f 69 6d 71 65 70 6e 7b 70 80 7d 81 7c 7a 76 7f 7e 7a 7d 7a 7e 81 86 85 86 8f 88 90 99 99 95 99 9d a3 a5 a2 aa a2 a5 a1 9f a6 a9 b1 af af ad b2 ad b7 b6 b6 af b7 ad a8 9f a5 95 a4 9e 9b a7 a8 a6 a2 a2 a0 a0 a8 9d 9c 9d 98 94 92 8c 8f 8d 89 91 92 90 91 8c 96 93 91 9e 96 94 95 97 96 94 95 99 94 96 8c 9f 97 8f 96 93 87 8e 7f 8e 93 91 97 94 92 99 96 a0 9e 97 9a 9a 99 a2 9f a1 a1 a4 a8 a6 a1 a6 a6 a3 9c a1 a5 a0 9e a2 a6 aa a8 ae b1 b8 b6 b6 b2 b0 b1 b3 b1 b0 aa ae a8 b7 b5 b7 b9 b3 bc b8 b3 b9 ae b5 b1 ab a9 a9 a2 9b 9e 9e 8f 93 8b 80 7a 7d 86 79 71 7a 77 75 71 73 6f 75 79 7c 79 77 6e 70 79 76 81 a0 bb c7 a6 a0 86 75 62 4f 42 2c 22 19 12 12 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 1d 22 32 39 45 61 7f 8c 6a 5b 5d 57 5e 5f 60 5d 64 57 5a 61 69 6e 6c 6f 6c 6e 68 6e 6f 70
 7b 7e 76 80 86 84 7d 7f 80 86 82 7f 86 7f 88 82 8a 81 8e 95 96 93 9b 9c 98 9b a0 a7 97 9c 9c 9f a3 a9 ac b1 ab a6 ac aa ae ac a3 b3 ae aa ad a6 aa a6 a9 9b 94 9a a0 a4 a0 a4 a2 9e a4 a3 a7 9f a5 a1 9a 96 9a 9d 96 99 8d 91 94 94 90 93 96 94 8d 89 93 92 91 98 90 92 92 96 93 90 94 91 94 8f 8e 93 89 94 88 96 93 a1 8e 96 88 9b 99 98 a3 a2 a2 a3 a3 a5 a1 a9 ab ad ab a4 a3 ad ac ad a6 af b0 ab b0 a8 b0 af a7 b1 b0 b8 b5 b8 b5 b1 b3 b8 bb b1 b3 b1 af b9 c0 be c1 b4 bc b5 bb b7 ba bd bb af a8 ac 9a 95 9c 9a 98 96 88 7f 7b 81 7f 76 7f 7b 7a 7d 74 75 72 6f 7b 80 74 74 78 6a 72 76 7a 91 bf c8 c2 ad 98 80 6f 5d 50 46 28 23 21 17 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 09 11 13 22 36 4a 51 63 7d 95 88 61 5b 57 5e 60 5f 5e 5f 5b 5f 61 63 70 6e 73 72 75 72 76 78 76 78 78 7f 78 7b 7f 86 84 84 81 85 88 83 84 8e 7f 8d 8a 85 8e 94 92 9c 95 9b 96 9a a4 a1 a3 9b a1 a1 9c 9d a0 a7 a8 a9 b1 ab ab a4 ac b1 b0 a9 a6 a5 a8 a1 a2 9d 9a 9c 99 94 9f a0 a6 ae a2 a0 ab a1 a5 9f 9f 9f 96 9c 97 93 9b 9a 96 95 90 8c 91 8d 8e 8e 92 92 93 8f 92 84 8b 90 8d 91 8c 91 8e 94 90 96 91 96 98 94 9a 94 9e 9f 9c 99 a1 9a a0 a8 a3 a7 b0 a8 b2 b2 ac b5 b5 af b4 b8 b3 ad b5 b0 b3 ae b2 ac b4 b5 b1 b3 b8 b8 be b2 b6 b3 be b5 b5 a6 b0 b7 b7 b8 ba bd bf bd b5 c0 c1 b7 c0 bf b4 b6 a6 a8 9d a1 9a 91 90 8d 8c 8d 80 81 85 76 77 80 74 7e 71 75 80 78 7c 74 77 7d 72 75 72 72 76 82 ab cc c7 bc 9f 90 80 6a 5d 4c 44 35 22 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 0c 14 17 2a 40 52 66 80 97 90 6e 59 56 5b 60 62 5e 5f 5e 5c 65 68 6e 6e 72 74 75 76 7e 80 74 6d 7b 7a 7d 7e 7a 7d 87 80 89 89 7c 86 80 7e 86 83 84 8d 87 92 8e 93 95 95 91 98 9f 9e a2 9b 9b a0 9b a1 a0 a3 a4 a4 b0 a6 a9 b0 a5 a4 a6 a7 a9 a7 a8 a5 a3 a1 9b 99 9a 97 95 9e 9a 9f a4 a0 a7 a5 9e a7 9f 9c 99 9a 97 96 96 93 92 8c 94 90 94 8e 8f 92 90 53 97 93 8f 94 93 88 92 89 8c 84 8f 87 98 94 8c 95 90 93 91 98 95 9a 9b 9a a5 99 a4 a0 aa a7 ad a9 b7 b2 b0 ad ad ba b8 b5 ba b8 b8 ba ae b2 ac af ac b4 b3 b4 b2 b5 af b5 b8 ae b5 ad b1 bb ae b4 b3 b9 b9 ba c2 bb bd be c0 bb be b1 bb ae b0 a4 9d 9b 99 96 90 8d 8e 8a 87 83 7e 7b 7a 77 81 75 7b 73 79 70 7d 76 7b 74 79 75 6f 6a 6c 75 76 94 c0 c2 b7 ab 9d 89 7e 6a 54 48 3d 2e 1c 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0d 0e 1a 25 37 4b 58 7e 91 a0 8d 63 64 61 55 5f 55 60 68 5d 6e 64 5c 6a 71 78 79 79 7f 7d 7c 7b 7b 7d
 7e 7d 7e 7b 8c 82 85 8a 83 8c 88 84 8a 8c 89 94 8d 8f 93 90 96 9b 96 8f 9d 96 97 9f 99 9a a1 a2 a3 a3 a2 a4 a3 a1 a4 a1 a6 a5 a8 a8 a7 a0 a3 a1 94 96 97 9b 94 8f 91 96 94 9a a5 9a a1 9d 9c a6 ab 9d a4 a6 a1 9f 99 9e 9d a0 9d 94 98 8f 9a 8f 8d 8f 79 90 8b 8b 8d 8c 8f 90 92 99 92 98 90 9a 97 9e 95 96 95 96 97 9c a3 9f ac a3 a1 a1 a9 ae aa ac b4 bc b1 b1 b4 bc bf be c2 c2 b6 b9 bf b9 b5 ba b7 b1 b3 b0 b5 b4 b8 b0 b7 b1 b4 b6 b5 bc bf af bc ba b6 bb ca c8 c1 c7 c6 c5 bd bb c0 c0 ad af aa a4 9b 9d 98 8a 8c 8d 8a 86 83 87 7b 82 75 78 6f 76 76 73 74 72 73 72 75 79 6c 6b 76 6c 75 76 89 ae be c9 be a6 9a 85 75 5b 4c 3e 2a 17 0b 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 0b 1c 28 2f 46 58 71 8b a8 99 76 65 57 61 5e 6b 5f 6c 63 68 6d 62 67 6e 74 73 74 79 7d 81 7b 80 74 88 84 80 7d 7e 86 81 88 7f 8a 89 8c 82 90 8d 8e 91 93 91 96 93 98 9c 9b 96 9b 9f 9b a3 a0 9a 92 a1 a1 9f 9e aa a3 a7 a3 a8 a8 a0 a2 9f 9d a6 9b 9a a0 95 9a 92 8e 95 96 96 95 99 9a 9a 9c a5 a5 a5 a0 a0 a0 a6 a4 9f a1 9e a0 9d a0 99 98 99 95 95 94 93 9b 91 99 9d 95 97 94 8e 93 95 99 96 97 90 96 97 a1 9f 98 9b 95 a7 a5 a5 a3 a9 a6 b0 ac b1 b4 b1 b7 b4 b5 bf c4 c3 c1 c8 c4 cb c0 b5 bb bc b9 b9 b9 b1 ad ab b0 b0 aa b1 b4 b5 ba bc b5 b5 c2 b6 ba c2 ba bb c6 c4 c9 cc bb bf c0 b7 b9 b1 b7 a7 a1 a3 9e 94 91 9a 8e 82 8a 85 83 85 7e 74 78 7e 7e 80 75 7c 76 75 75 77 6f 74 71 6d 6a 72 72 7e 7b 99 b8 b8 bd b5 9c 8e 7f 68 54 3b 29 15 0c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 12 11 27 3f 48 62 7f 9f a5 83 6f 6b 60 65 63 6a 63 62 6a 5f 67 64 6a 76 6e 79 77 75 7c 78 84 7c 7d 84 7e 7c 84 88 88 80 88 89 89 81 8b 8d 8a 8e 8b 99 93 8d 8d 90 9a 9c 96 93 95 9c 9f 94 98 96 94 9a a1 9e a0 9d 9d 9b 98 9a 9e 9b 9c a2 9d 99 96 93 97 97 98 8d 8b 8d 90 8e 97 97 97 9a 99 a7 95 a1 9c a4 a0 a7 a2 9e a6 a4 a8 a4 a1 9a 9e 9a 96 a5 9c 9d 96 9b 97 9f 92 91 99 9a 91 96 94 96 96 98 99 9c 95 9d a1 a1 a0 a5 ad a7 a3 a2 b0 ad b0 ba bc b8 be c3 c0 c9 c1 c2 c5 c8 c7 c1 c0 b6 b5 bd b8 b4 af ab af ae ae ae b0 b0 b1 bb b4 b1 be bc b7 b8 ba c5 b4 c6 c1 be be c3 c5 c1 bb be b7 b4 ae a6 a9 9e 92 8f 90 8a 97 86 84 84 7b 83 81 80 7b 7f 7a 75 7b 7a 7b 76 7b 6f 70 73 71 70 6b 7a 75 77 74 84 9d b9 bc b0 a1 94 83 72 55 47 25 23 09 00 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 16 14 18 33 45 56 70 83 9d 93 78 77 64 6b 66 5f 67 6d 63 63 66 70 6f 6c 6f 69 79 77 77 75 6f 7d 79 81 85
 89 86 83 84 8b 89 8b 84 8e 8f 87 9c 93 87 93 95 91 91 95 94 9c 9b 94 9a a4 9c 9f 9a 97 99 9d 9e 9d 9f 93 9c 9b 9f a0 a4 a0 9c 9e 9b a1 98 94 8d 96 8b 8b 8b 8b 8c 90 86 8c 90 97 95 99 9a 9f a1 9d ab a0 a5 a1 a9 a6 9e a3 a2 a8 a0 a4 a1 97 a4 9a 98 99 9c 98 9b 9a 95 9d 97 97 9c 9e 99 a0 99 99 9c 9f a6 9e ae a9 ae a5 af a4 ab b1 b2 b9 b8 bd c2 bd c6 bd c8 d0 cb c5 c7 c9 c0 bc b9 b0 b8 af ae ac b1 b1 ae b6 ac b3 b2 b1 ae bc b0 c1 b8 bd b7 be c1 bc c4 c3 bf ba bf b6 c2 b8 b5 ae b3 b3 a9 a4 a2 97 96 8b 86 8e 7e 88 79 75 81 81 83 76 83 7a 84 7d 78 79 7f 73 6e 74 6e 65 69 75 71 77 68 74 70 8b af b9 c1 ac 92 84 6d 59 4a 32 29 17 07 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 02 06 10 11 1d 1b 1f 33 46 60 7e 88 94 81 6e 72 6d 68 6d 63 64 68 67 65 6c 6d 71 75 75 70 7a 78 74 7f 81 7e 7c 86 79 80 87 7e 7b 8d 86 8a 93 97 85 95 92 94 8a 8e 8a 8d 92 8d a0 9e 9e a2 a4 a0 a3 a0 98 a2 9f a1 9b 98 99 a2 9e a0 a2 9a 99 a4 9a a1 98 9c 98 8a 91 92 86 8b 8d 85 89 8b 88 8f 8d 8d 9a 94 98 9f 9a a7 a0 a7 a1 a1 a7 a7 a8 a5 ae a8 a5 a8 a3 9f a7 a1 a0 a0 a1 9d a0 9f 9b 90 a3 90 a3 9e 99 a1 a2 9a a9 a4 a8 a6 ae b0 ad a7 b1 a7 b1 b5 b1 b2 ba c3 d0 cd ce c5 c5 c7 c2 c4 c1 bb b9 bd b0 ad b6 b7 b9 af b3 b0 b4 b1 ae b5 b7 b9 b7 b4 bb b9 b9 b9 b4 c0 bc bb c7 be c5 c6 b7 bf b4 b4 af b4 b2 a0 a6 9b 99 93 8d 91 93 8d 8c 85 84 78 81 7e 84 8c 78 80 82 79 7b 77 7a 73 74 72 7d 68 6e 75 6e 69 76 6b 76 71 88 b2 b0 a9 97 7a 6d 66 5e 4d 3d 25 0e 0a 05 0a 01 06 05 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 13 16 16 21 30 40 4c 63 6a 7d 7b 7a 70 73 70 6e 6a 6a 5c 63 61 6c 72 6c 65 6e 78 75 75 74 74 76 7c 77 84 83 7f 83 7f 82 81 8c 8c 8b 92 91 8c 8a 8f 92 93 90 8f 88 94 8e 93 9a 9b 99 9e a0 9d a0 a7 a6 9f 96 a1 9d 9b 9c 98 96 9d 95 95 99 9f a3 9b 99 98 8e 8e 91 8e 8e 84 85 8e 85 8b 81 85 8c 8e 92 94 92 96 94 98 a2 a7 a8 9a ae ac a9 ae a3 ab a6 a9 a8 a6 a1 a5 a4 a3 a2 a5 a2 a4 a4 a5 a0 9c a4 99 a4 a3 a5 a1 ad a6 a3 af af b4 aa b0 b1 b7 b6 c1 b9 b5 c4 be ce cc c3 cf c3 c0 c4 b9 b4 be b5 b0 b1 b9 ac af b9 af b2 b1 b8 a9 b5 b7 b3 b5 b3 bb b2 c2 c3 bb c7 c3 ba c4 c0 c5 bf b9 b8 b5 b4 af ad a4 a3 a4 9e 94 90 8d 89 85 88 88 84 89 83 83 7d 84 7b 82 81 79 74 70 6f 75 6d 75 6b 6b 6c 6e 77 76 6f 6d 6c 70 67 73 9b 9a 97 7b 6f 65 5d 62 53 40 30 21 12 0b 06 09 07 05 03 00 06 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 12 14 1f 22 22 2c 3c 4f 62 5f 6b 7e 80 7a 6c 71 70 6a 68 6c 60 63 6d 6f 70 6a 66 70 71 7b 78 7e 7c 7e 7c 7c 85 7c
 86 7f 84 89 85 89 86 8d 85 8f 90 92 97 94 9a 8e 9b 94 8a 9b 96 94 a1 9a a4 a4 a1 9e a3 9f a3 a9 9f 9f a2 9f a2 9e 99 9e 9b 96 99 94 92 90 8c 86 8d 8d 7f 88 7d 84 86 82 84 90 8e 84 93 90 93 99 9d a2 a0 9f a8 9f ae b2 ac a6 ac a7 ac ab ad ad b1 ad ae 9f 9d a8 9e a5 a3 9e a6 9f a7 a2 a5 ab ac a7 ab ad ab aa ab ae ae ae b7 b9 ba ba c7 c5 cd ca c9 ce c8 cb c2 c6 bf c5 b2 c5 bb b0 b1 ae b2 b1 ab ae ae af bd b1 b1 b5 b6 ba be c3 bb c7 ba be c6 c3 c0 c1 c6 c2 bb b5 bb b4 ad ad a7 9e 9f a1 94 98 91 8f 8b 90 8c 88 86 85 7b 83 81 7c 83 7c 75 7f 7c 73 73 75 6a 71 73 77 75 76 73 70 6e 61 66 68 6b 6d 75 87 7a 73 61 65 71 68 60 52 3a 23 17 0d 08 00 06 05 05 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 1b 1f 25 2c 33 35 3f 44 4b 53 5e 60 6d 77 83 84 78 6e 6e 68 6b 68 67 67 72 70 66 67 76 76 77 74 78 76 74 77 7d 85 86 7f 7e 82 8c 8f 87 87 8e 91 8f 88 8f 92 98 9d 91 99 99 9a 99 96 94 9b 96 9a a2 97 9e 9d a0 a6 a2 a3 a4 a3 a5 9f 9f a5 a5 a5 9b 91 98 98 8f 95 8a 86 85 84 7e 85 83 85 84 88 85 8b 8c 85 8c 8a 96 9d a2 a2 a4 a1 a7 ab af ae a6 a8 ab af af a0 b1 af a9 ae b2 ab a5 ac ab a6 ad ab a9 a3 ab ab af aa a5 b5 b6 ab af b8 ae b3 bb b5 c1 c0 c3 cc c6 ce d3 cc cf d4 c6 cb bf be be b0 ba b8 b0 b1 b1 b1 b5 ba af b9 af b6 b5 b6 b7 b9 c4 c1 b8 c7 c1 c9 c3 bd c3 bf c3 c1 c5 b4 ba b7 ac a3 a6 9d a1 98 92 8e 8e 96 8d 90 88 86 86 84 81 85 80 7d 82 83 83 79 81 78 79 75 75 71 74 76 71 6d 75 76 73 69 6b 64 6f 67 70 66 77 79 5c 5b 54 6d 7a 6b 60 4b 30 1e 15 0e 0f 06 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 11 1a 25 2e 39 45 4f 50 54 50 52 59 5e 69 73 83 85 81 75 67 69 69 6c 68 68 71 6c 71 6f 69 6d 78 6f 76 7d 7c 7c 78 78 76 88 7c 85 84 8e 80 8c 8d 8e 98 96 95 96 93 92 9e 98 9a 9a 94 99 96 9a 9b a4 a1 98 a2 9c 9e a2 a5 a6 a7 a6 aa a9 a9 a7 9b a0 9f a4 96 90 95 8e 87 8d 83 86 7c 7e 80 7f 7b 85 85 8a 88 8d 8f 94 95 9c 97 99 a1 a4 a3 a7 aa aa ab b3 ac b1 b3 b5 ae b6 b0 b2 ab ad b0 af ad ad a9 a7 a6 b3 b0 a6 a8 af af ad b3 b1 b0 b8 be bf c5 bf c1 c5 cb ce ce d9 de ce d1 d3 c9 be be b8 c0 bb ba b3 b6 ae b8 b0 b9 b1 b7 b9 b9 b7 ba b5 b6 b6 bd bf c6 c3 c2 c7 c2 c4 c4 b9 c2 bb bc b3 af ad ad a4 a6 99 a4 96 91 98 96 8e 8e 8c 89 85 89 87 8c 87 84 81 7e 7d 82 82 7e 76 79 73 75 76 70 76 75 73 70 63 67 6c 68 66 6a 60 67 60 73 61 5b 54 55 6e 7a 71 63 50 3b 2b 20 13 0e 09 05 0b 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 17 26 28 2b 31 30 42 56 5c 4e 52 55 59 65 6f 79 82 81 81 82 78 71 68 6b 69 67 68 67 69 73 70 7c 7a 7b 77 82 7c 76 7f 7f 78
 7b 7c 81 84 7e 90 82 8b 8f 92 8e 94 8f 98 97 96 95 95 96 9a a2 9f 99 99 9b 9e 9a 9d 9c 95 96 a3 a3 a1 9e a3 a8 a9 a6 a5 a5 a4 9e a1 97 9c 96 84 8c 86 88 80 7a 79 70 7c 87 7d 85 82 87 89 94 8b 91 92 9a a0 9f a1 ab a9 ab b0 a8 b4 b0 aa b1 ad b5 b0 b6 b4 b1 b2 b5 af b7 b0 af a8 b2 b0 ad ac b3 af ad b5 ae b8 c0 bb bf bd c1 cd cb d1 d6 d9 da d6 de d3 cd cd c8 c0 c3 c1 b0 b6 ba b3 b5 ba b2 bc b3 b8 b3 b5 b9 c1 bc bd b9 bc c4 c1 c1 bc c5 c4 c0 c4 c0 b9 b4 b5 b3 ab ab a4 a2 9a 9a 97 94 96 99 96 8d 89 92 85 8b 80 7c 80 7c 85 7d 7f 7d 85 81 7d 6e 71 74 78 7c 79 7a 78 73 72 75 69 6d 68 68 63 6a 67 6b 6b 5e 4f 55 4f 60 70 76 6d 59 41 2d 28 19 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 07 19 29 2e 39 2f 3a 39 4d 5e 55 5b 5b 56 5f 67 73 79 7e 7d 7f 7a 7a 70 68 68 67 6e 6d 70 68 70 72 7c 7a 79 7d 7c 7c 7d 81 7b 79 7a 84 7b 8b 81 86 8b 92 8c 91 8f 97 91 8d 9b 97 9b 97 9d 95 9d 9d a4 98 9b 9a a2 9f a0 9b a2 a1 9c a6 ab ae af 9f ab af a9 a6 a7 9e 9b 89 8e 8c 8b 83 84 7f 79 7f 84 7c 83 86 8a 88 8a 95 90 94 96 99 a3 a0 a0 a7 aa aa a9 ac ac b2 bf bd b0 b6 b2 b4 bf b7 b0 bc b6 af b0 b9 b6 b2 b3 b5 b6 b1 b1 b7 b5 b4 b6 bb c1 c7 c4 d1 ce d0 e1 dd e5 e4 e8 db da d2 cd c8 c1 c5 c0 ba be b9 b3 b9 b8 b5 c0 b5 be bc c3 be be c1 be b6 c3 b8 c1 c3 b9 c9 bd b9 c2 be b9 b4 b6 ac ad ab 9b a3 97 92 96 97 92 97 88 91 8c 91 84 8b 86 88 86 86 84 88 7c 7a 81 73 7e 77 7c 75 6a 7c 7a 7e 78 74 74 6d 6b 72 64 62 6b 6a 64 71 6f 5d 56 4f 4e 53 71 77 6d 62 4c 40 25 16 19 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 09 1b 28 33 32 3f 44 38 35 45 55 52 62 66 63 67 65 6d 6c 73 7f 7a 79 7a 79 71 67 64 61 65 72 6c 6f 7a 75 77 70 77 7c 72 74 80 7e 81 7b 80 85 8b 83 8c 89 8b 96 87 8d 94 96 96 99 9d a0 9c 9e 97 9e 98 a0 a3 9f 9d a2 a4 a0 a0 a6 ac a4 a3 a7 aa ad a3 a3 a4 a4 a4 a3 94 95 92 8c 91 87 82 84 7f 84 84 84 7e 81 85 80 88 8b 8a 87 92 92 99 96 a0 a2 aa a8 a5 ae b5 b2 b4 b4 b1 c0 b8 b2 bb b6 b2 b0 b4 b5 b3 ba ae b3 b2 ba b9 bd bd bd b7 b9 ae c0 bf ca d0 d2 cc d8 d8 e4 ea e4 e3 e0 da dc ce cd c5 c2 c4 be bd b9 b8 c4 ba bb bb c1 b6 b7 ba bd b7 b9 b8 c1 c3 be bd b8 b6 bd c8 b3 bc bd b3 b4 b5 ad a9 aa 9f a2 9d 97 95 93 9b 91 97 91 87 85 84 82 89 81 83 84 7a 86 79 7a 7f 7d 7c 7d 6e 7f 82 77 7b 75 77 74 71 74 6d 70 62 70 68 66 69 6e 69 62 5f 55 55 4a 55 6c 81 7f 62 5c 43 35 23 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 11 1e 1c 27 36 44 47 4e 47 4a 4a 50 5b 5b 64 60 64 6c 6c 6f 72 71 77 7d 78 6f 76 74 66 6c 6d 64 72 67 76 72 6f 75 70 78 7b 77 75 80
 7a 79 82 80 85 87 84 8a 8b 86 8c 8f 92 99 98 99 9b 95 a4 9d 9c a3 a2 a1 a3 a9 9f 98 a1 a2 9a a0 a3 9d a7 a3 a3 a7 a6 a2 a5 a1 a5 a1 99 93 8f 95 87 86 85 81 89 82 7e 74 7f 7d 86 82 8a 8c 8a 90 91 94 96 99 91 9e a7 a9 a6 ab b1 af b3 b6 af be b5 bd b9 bd be bb b3 b6 ac b2 b4 ba b9 bc bc c2 b9 ba b7 c1 b3 c1 c7 c8 cf da d9 e1 e8 ea ea e5 ea e5 e0 d4 d1 c7 c4 c9 bf c0 b5 b7 ba b9 c0 b9 b7 be b8 b3 b4 ba b2 bb b5 b8 b9 bc c0 bc bf b3 c0 b4 b6 bb ab b3 b0 a5 a8 a1 98 9e 9a 99 95 91 98 8a 8a 8d 8d 86 86 88 88 81 7e 7e 7b 80 85 79 83 7e 79 75 7e 79 75 73 75 70 6d 70 6f 64 6a 6d 68 64 66 66 6a 6b 66 61 59 59 4e 48 4e 67 77 7c 73 5c 45 2f 1b 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 17 25 25 2e 44 44 51 5e 55 4f 4e 56 5d 61 68 69 60 65 68 6d 6b 73 71 71 7a 77 74 74 74 71 71 73 73 72 77 6a 73 75 79 7a 79 74 7c 7b 7e 81 7a 82 87 84 86 89 88 8a 8e 8e 95 93 95 a2 9f 9e a5 a2 9e a9 a9 a4 a9 9e a6 9f a4 a3 9f a3 aa a3 a7 ab a2 aa aa a7 b1 a4 a4 a2 9a 99 8d 94 8e 83 7e 82 7e 86 7d 81 85 7a 83 86 85 85 8c 8d 92 8d 95 9c 9c 9f a6 a4 aa ae b6 b4 ba b7 c0 c5 c1 c2 b9 b8 bf bd b9 c3 b9 bc be c1 bd ba bc bf bc bb be c3 c8 c2 cd d3 d5 e1 e3 f2 ee f0 f8 f1 e7 e8 e2 da d1 d3 c9 bf bd c6 be bb bc c2 c4 b8 b4 c4 b9 ba b9 b9 c1 bb b4 b8 bc bc b6 b8 b8 b5 b4 bc b9 b6 b0 af a6 a4 ad a5 9d a1 99 97 92 90 95 8c 90 8e 8b 85 8e 81 88 83 85 87 7f 87 7c 7c 77 7d 7c 7d 7e 7d 7a 77 73 74 6d 72 6f 67 69 6d 6c 69 62 66 67 6d 6f 73 5c 5b 56 4e 51 65 7e 80 72 5e 50 37 1f 16 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 14 1c 26 25 3d 46 50 5d 62 5e 56 4b 62 59 5e 6d 67 63 69 6a 63 71 6f 68 70 6e 73 70 6f 70 6d 75 6c 71 71 6d 70 75 77 76 80 74 76 77 77 80 80 7f 80 80 85 85 7f 85 8b 87 8f 92 9d 98 a1 9d 95 a5 a4 9e 9f a2 a3 ab a9 a1 a6 a8 a3 aa a5 a5 ad a8 af a0 aa b1 a6 ac ad ad a9 a4 9f 9e 98 92 8b 8d 88 84 81 89 84 85 8b 88 8b 8c 8f 8c 94 93 9f 9e 9a a1 a2 ad ab ae aa ad b8 b4 be c2 c9 cc ca bf c4 c4 c6 c4 c2 c0 bd be bd c2 c3 bd c3 bd c0 c9 c3 ca cc d2 d9 e0 dd e7 f5 f4 f2 fe ec e8 e6 d9 d9 cf d0 cd c7 c3 ba bd c1 b6 b6 b3 b9 b4 b9 b7 b2 b7 b3 bb bd ba bc ba bb bb b7 b8 b9 bf b8 b4 b5 b0 b0 b0 a4 a9 9c 98 9c 96 92 95 92 95 8c 8f 98 86 83 87 88 8a 80 82 84 81 83 85 80 7e 79 7a 79 7a 79 7d 7d 6e 76 75 73 73 71 65 69 6d 69 64 6a 6d 71 70 67 67 5b 53 4a 58 5e 73 83 72 60 4f 41 28 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 14 15 26 2a 43 44 56 5d 6b 6b 54 53 51 5e 5e 5b 5e 64 6a 61 63 65 65 68 64 6e 6e 75 6f 68 6f 74 6f 75 6f 6c 77 77 72 75 77 78 79 7a 79
 83 79 81 7a 78 82 7f 87 8a 8c 90 91 9a 92 99 9f 9b 9e a2 a0 9d a5 a5 a5 a3 a4 ad a7 a2 af a9 a9 a8 a9 ad aa ab ab af ab b2 a4 a1 a8 a0 9f 97 9c 8f 91 90 8e 8c 88 8a 7a 8a 8b 81 8c 86 90 97 94 93 91 97 9d 9c 9f ab ae b1 af b1 ba c5 c5 c9 cc d5 d4 d1 ce ca cc ca d0 bb c1 c2 bb c1 c2 b8 bd c3 c3 c4 c9 c7 d3 d7 de e1 e7 ee f4 f4 f7 fc f6 ec df da cc ca c5 c0 c1 c3 bc b7 be b9 b4 b3 b8 ba b8 b9 b6 b7 b7 ba b5 b6 b1 b9 bb b7 b4 bc bb b6 b1 b2 af a6 ab a7 9f ac a0 94 99 95 94 90 91 93 8d 8b 8b 83 86 81 84 8c 88 85 81 77 7b 83 79 81 7a 7b 7e 75 7d 6f 75 77 76 72 64 70 6f 69 61 6a 65 61 62 6a 73 77 75 71 60 5a 54 4b 56 73 80 79 62 54 3c 23 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0f 0f 22 2f 30 43 4e 55 71 74 6b 58 53 54 5f 60 5e 64 66 67 60 63 65 65 6b 64 6c 6e 68 6e 68 68 6e 66 6d 71 6b 71 78 70 77 82 75 80 84 7d 7e 7b 82 81 7f 81 85 87 89 86 8d 94 91 96 94 9c a8 9d a3 9e 9e a3 a8 a5 a7 a5 a5 ad b4 ad ab a6 b0 b4 ac b3 aa a8 ab a5 ae a9 a2 ad a1 a5 9f 97 99 9d 95 95 87 89 85 89 83 88 8c 8b 93 93 87 8f 99 97 95 9e a5 a7 ac aa b3 bb c1 c4 ce c9 d4 d3 d3 d8 d7 d7 c9 dc d7 d6 d7 ce c3 c6 c6 ce cf c5 c5 c7 c3 cb d2 db e8 e5 eb ed f5 fa fa ff f8 f2 e8 e0 d5 d5 ca cc c6 c3 c4 be ba b7 b3 be b3 b7 b5 b6 b0 bd c0 b6 b9 b8 af b1 b9 b5 bb af a8 ba bb b0 bb ad ad a4 aa ac a0 a0 9b 91 96 94 92 8e 92 83 87 8d 82 87 88 7f 86 7e 84 83 7c 80 7d 7c 7d 7a 76 7a 76 73 79 71 77 6d 69 74 69 69 66 69 6d 5f 63 66 6f 7b 7d 71 77 65 5b 53 50 5a 70 7e 7b 6a 51 3d 25 1b 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 08 20 26 2b 3e 45 53 5a 73 73 6b 55 4e 57 55 5d 61 5a 62 62 61 61 68 6a 68 62 69 6c 6b 6b 6b 6c 6e 74 71 75 68 6b 69 6f 74 79 7e 7d 7e 7e 87 7f 83 80 83 80 85 88 8b 8d 8c 93 91 9c 99 95 9c 97 9f a1 9e a0 a6 a5 9f a6 ae 9f aa af a5 ba b5 b1 ad b6 b2 b0 b3 af b4 af b2 aa a1 a1 9d a8 9c 8f 94 8b 93 96 8e 85 8e 8b 8e 8c 93 93 91 91 99 9c 9a 98 97 a5 ad b4 bc c3 c7 c9 dc d6 e2 e2 de e8 e6 ea e9 e9 ea ee db de d3 d2 c9 cd cd cf cd d6 d7 e1 da df e8 ec f3 f9 ff ff ff fa fb e5 e1 e3 d8 ce c8 c7 ca bd be b8 b9 c1 bb bc bf c2 af bb b1 ab b2 b6 b4 bb b5 bb b7 b7 b5 b9 b9 b5 bb b0 b0 b0 ae aa ab a5 a0 a0 9c 9a 96 8f 95 8b 93 93 8e 97 89 82 85 8a 80 8d 83 83 7e 83 7c 81 78 7b 78 7f 76 76 76 68 6e 71 69 6e 73 68 65 64 63 5d 61 68 70 7a 76 6f 6a 6a 67 56 58 61 70 7e 7a 6e 5c 41 30 1b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 06 0f 1c 40 3a 48 5b 5d 70 74 63 55 4a 50 54 55 61 56 5d 5a 5a 64 66 65 64 65 62 67 6e 6c 6f 75 6b 6c 6f 72 70 6f 6c 74 76 77 76 71 7d 73
 81 80 7a 81 83 83 88 86 87 8d 89 86 8d 93 93 95 a0 9f 98 99 a3 9f a5 a4 ae ac a4 a9 a9 a8 a9 aa a8 a9 ad bd b6 b3 b8 b0 ac b0 aa b7 aa 9f a5 a3 9b 9e 9c 93 8f 91 91 8d 8f 93 90 94 8f 95 97 98 95 93 aa 9b a9 a6 ae b6 c9 c9 d5 e1 f7 fb f5 f2 ed f2 eb f1 f5 fd f9 f7 f1 e8 da d8 d5 c7 d0 ce db e1 e7 e2 eb e7 f3 f6 f9 fd ff ff ff f6 f2 ed df d6 ca c3 c6 bd c7 ba b9 c4 bc b8 bb bb b6 b9 b8 b8 b9 b1 b2 b8 b5 ba b9 b7 b3 b5 b4 b3 c1 b5 b9 af ad af ad aa ad a1 a1 9f 9c a0 9a 93 94 90 8b 90 85 86 84 84 89 76 80 7c 85 84 7b 7d 7d 74 78 7c 7e 7b 79 71 75 70 70 72 72 6c 62 61 66 5d 60 5e 5f 67 6b 6a 71 65 6e 6a 65 61 5e 64 6c 84 7b 71 5e 46 2f 20 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 0a 0f 20 38 3f 51 55 6b 6c 70 5a 55 51 59 56 51 56 5e 5c 60 60 5d 61 64 65 66 64 6e 6b 6e 66 71 68 6b 63 6c 6d 6f 6f 6f 73 75 73 7a 88 81 81 7c 7c 79 84 81 7f 82 85 83 85 93 8e 8e 93 98 9e a2 93 9f 95 9e a6 a2 aa a7 a2 a7 ae ab ae a9 b6 ad b4 b3 b7 b3 b6 b4 b0 ad af a6 ae ae a0 a7 9b 92 9b 96 92 99 9d 96 96 98 96 98 94 9b a1 9b 91 a0 a0 97 aa a1 b6 c4 c8 cd dd fa ff ff ff ff ff fb f6 f8 fe f9 f8 f5 fd f2 f1 de d7 df e3 e4 ee ec f4 f9 f9 fc fa fe ff ff ff ff ff f6 f9 e5 dd d2 ce c7 c2 c5 bc c4 c4 c1 c2 bb b7 bb b6 b4 b1 c1 b9 b9 b2 b3 b2 b3 bb bb b6 bf b6 b2 b2 af ba af ac ab ab a5 a2 9e a6 9d 9c a2 9b a1 95 99 92 8b 8b 85 85 86 85 86 8a 79 7f 7d 78 7c 77 7a 7e 7c 78 7a 80 76 6f 74 6d 6d 6e 6b 5e 66 62 6b 5e 5f 59 68 65 6d 6c 69 72 73 66 60 63 5f 73 84 80 71 5a 48 2e 1e 10 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 0d 14 16 36 45 53 5c 60 74 65 52 56 56 57 50 56 59 54 5a 60 59 61 61 64 63 5c 60 66 65 70 72 6f 71 71 6d 6e 78 72 6f 70 78 76 6f 80 7d 79 78 7c 82 80 81 82 87 8d 88 86 8f 8e 8c 8d 93 94 97 9f a0 a1 9e a2 a9 a2 a6 9f a7 a9 af aa aa b3 aa b4 b0 b4 b9 ac ac b0 ba b0 b2 b4 af ac a5 a1 a4 9b 98 9e 9e 9d 9a 9c a6 a0 a1 9f 99 a0 9f 9f a3 a0 9e a4 a3 ac b8 c4 cf e1 e1 fb ff ff ff ff ff ff ff ff ff ff f7 f8 ff fa fb f2 ed eb f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 f1 e0 d6 d3 cd c3 c7 c5 c2 c2 bf c2 bd c1 bb b9 b6 b8 c0 bb bc b3 b9 b1 b8 be b7 be b6 b7 bf b4 ae bb b8 b0 aa b2 aa a8 9f 9a 9b 9f 9e 9a 9a 9a 97 94 8e 90 91 8d 81 8f 81 81 82 84 85 7f 86 78 7a 7d 7d 78 7b 75 6e 72 76 6e 6b 6a 72 6a 68 63 65 61 5f 60 60 67 69 63 6a 6b 78 68 66 61 61 67 68 7f 83 74 61 48 33 1f 0e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 1a 29 3b 56 65 6a 68 5f 52 5b 4f 58 5d 5b 57 54 5c 57 59 54 59 5f 60 59 62 61 66 70 70 6b 73 71 65 66 75 6e 71 72 72 76 7a 76 7f 7e
 85 7f 7f 84 81 82 7e 86 85 8c 8f 95 8c 93 90 98 9a 95 96 9e a2 9d a1 a5 a4 9c a6 ac a9 ab b3 a9 ad af ab ba b3 ae ac b2 ae ab af a9 a4 a4 a4 a1 9b 9f 95 9a 9d a1 a4 a5 a9 a8 b1 b4 aa a6 9d 9e 98 a3 9c a9 a9 aa b9 c3 d6 e4 f0 fc ff ff ff ff ff ff ff ff ff f1 ef f9 f9 ff ff fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f2 e1 d3 cb c1 c9 c8 c9 c5 c0 c0 ba bc c5 bb bd b9 b3 bf c3 c6 b4 ba c4 b6 bf af b5 b6 b9 b6 bb b6 b7 b6 ac af a9 ac ac a2 a3 a4 a0 a0 98 96 98 94 93 8b 87 89 83 81 80 86 86 7c 82 81 7e 7f 74 7d 75 78 71 78 7b 6f 74 6a 6d 6f 70 68 6a 62 61 5e 5c 5e 5d 57 64 62 63 66 64 65 5f 71 5d 59 61 67 7e 86 72 64 4b 34 21 06 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 16 2e 39 4b 62 60 74 68 50 57 51 57 5d 55 57 5c 5a 61 60 5c 61 5c 5c 61 5f 60 66 67 70 71 71 73 75 70 72 70 72 70 76 87 73 7a 82 78 82 7e 81 83 85 81 8c 8e 8f 8a 90 8a 95 8d 96 97 97 96 97 9e a3 a0 9e 99 a7 a7 9d a5 a2 a6 a5 ae af ae ae b3 b0 ab a8 b4 b3 ae ae b0 a6 a6 a5 a2 9c 9e 96 9f 9e 9c a6 a8 b5 b1 c2 be b4 ac ad a1 a7 a7 a4 a9 b1 c2 ca d4 e7 f5 fb ff ff ff ff ff ff ff ff ff ff f8 ec f1 f3 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa f0 e3 d9 ce c8 be ca c7 c1 c7 be c9 bd c4 ba bb bc bf c1 b9 b9 bd ba bf bb c2 bd b7 bf bb b2 b4 b7 bb b7 ac b5 a1 a8 a9 9e 9f 9a a1 9e 9d 9b 9d 95 8d 8e 83 8b 8a 8b 8a 8c 87 7b 8d 7a 84 76 7c 7f 7c 83 75 76 75 74 72 6f 69 6d 60 68 68 60 5f 63 64 55 56 55 57 5b 60 5d 5d 5d 5f 5a 54 5d 5c 66 7f 7c 72 6a 4d 3d 27 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 0f 15 21 3f 4d 5b 6e 71 68 5d 54 54 59 5f 5a 5e 5c 5a 5c 5e 54 61 61 61 5e 5e 60 65 68 67 6e 6f 73 72 6a 70 70 72 72 72 7e 76 75 7b 7e 80 7e 88 89 7f 87 84 92 98 8e 8d 8b 8e 89 95 9a 9e 98 99 9d 9b 97 9d a0 9e a3 a4 a5 a7 a9 aa ad b0 af af b4 b6 ab b4 ae b1 ae b4 a1 a8 a0 9f a4 9f 9f 99 9c 9b a4 ac b0 b9 bc c6 c9 c5 c1 b5 b6 b8 b4 b6 bc c2 b9 da ea f5 ff ff ff ff ff ff ff ff ff ff ff ff f6 ea f3 f8 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 ef dc cf ce c5 d1 c1 c5 c7 bc c0 c2 c5 c4 c4 c0 c1 bd bd bd bb c4 c0 b6 b7 b9 b9 b3 b2 b8 a9 af b3 ad bb a9 a5 ac a8 a0 9e a4 9f 9a 9d 9a 92 9a 97 94 90 88 90 87 86 87 7e 82 85 80 86 8b 79 89 7b 79 7d 81 7f 77 6b 72 6f 72 70 65 67 68 65 5f 62 63 62 59 56 5b 52 63 5a 58 5c 53 5f 57 52 5e 65 7b 80 79 64 53 39 26 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 18 2b 36 3e 5d 6c 70 80 6b 59 54 51 54 5a 5f 5c 5c 60 5f 60 62 60 5c 5e 60 66 65 66 6d 69 6b 6e 6c 73 74 70 72 79 74 7b 71 78 7b 80
 7d 7c 84 84 83 8b 8d 86 8e 8c 8e 8d 92 8f 8e 92 91 8e 9d 9d 99 97 96 98 a1 a1 a7 a0 a6 a8 99 a6 ad ac a4 b1 a7 ac a7 ae b6 ab ad a5 a6 98 a8 a5 a3 a1 a5 9c a1 9e a2 b0 b5 c1 c9 d3 d5 d4 cf c4 c5 be bd cb d6 d7 ef ff ff ff ff ff ff ff ff ff ff ff ff fe f9 e6 e3 e5 f3 ff fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 f1 dd d2 ca d2 c8 c4 cc c5 bf c1 c1 b6 ba be bb ba b6 c0 be ba b6 bb b9 ba b6 ba b9 b7 b0 b3 b1 b1 b2 b1 ad ad b0 a6 9c a2 9c a0 a1 9d 95 a0 8d 98 8e 94 9a 8c 87 83 83 87 81 7d 84 81 82 82 81 7b 7d 79 77 75 7c 70 74 6d 6d 6b 70 68 64 6a 63 60 60 58 59 5b 5a 58 53 58 58 54 4a 52 52 4b 48 51 5b 82 7c 77 69 4d 38 20 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 08 14 16 28 34 4c 5a 67 70 7e 73 5c 5a 53 52 5b 59 5b 5c 5d 5b 5a 62 61 5b 60 61 5e 62 67 68 66 72 6e 68 70 72 74 71 6f 6e 73 7c 6e 78 7e 7d 79 84 84 84 87 8e 83 8a 85 90 90 89 93 93 90 93 92 96 99 9a 97 99 9b a1 91 9e a1 a5 9d a2 aa a1 a6 a4 b1 ab ac a8 ad ab 9f a2 9f ae a0 a2 9f aa a1 a2 9e 99 9f a1 a5 af bb cc e0 de ea e4 da d2 cf d8 d9 eb ef ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e9 de e1 e7 ec f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 e0 d5 d4 cb ce c7 c0 bd b5 c1 b7 b7 b8 b6 b8 bf af b5 b1 b1 b3 b8 b8 b3 b0 b0 ad b0 b7 ad b2 ad ad a9 af ae a3 a5 a7 9d 9d 9e 9a 91 92 9a 95 97 8e 8e 90 90 85 8d 8b 80 81 7f 7b 7d 7b 7d 76 7c 7c 77 75 73 77 72 75 71 6a 63 67 67 61 64 5e 53 5a 5a 64 59 49 56 51 55 57 4a 4a 50 41 53 50 4e 55 5c 7a 82 72 69 51 2a 28 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 08 09 14 28 2f 38 4b 52 66 7b 79 80 6a 59 59 4f 54 54 5d 5f 60 5c 61 57 66 63 64 67 67 64 66 6a 6b 6d 75 76 70 73 75 7a 75 71 74 78 78 7f 84 82 81 7e 85 8b 89 80 8b 89 8d 8f 92 8d 8f 8f 94 99 99 8b 92 95 9c 9a 99 a0 9e 9a 9f 9f 98 a3 a9 a5 a7 a9 b1 ab a4 ac aa b3 a9 a6 9d a8 ad a3 a7 ab 9f a4 a2 a3 a1 a3 b1 a7 b9 bf cb dc e8 e8 e5 ea e7 e8 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff fd de e0 db e2 e3 ee f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fc ee da d9 cd cd c2 c0 c7 bf b1 b3 b3 b4 b2 b1 ad ba a6 aa b3 b3 b0 a9 b2 a5 a9 ad ab af ac b0 a7 ac ac 9f a5 a3 a0 a3 a5 9f a4 96 93 99 9d 99 97 99 92 90 8e 8b 92 88 8a 7f 86 81 88 87 7a 80 79 7f 77 7e 7a 7c 78 77 62 6f 67 66 6c 65 62 64 62 61 5f 57 59 5a 54 51 55 5b 58 57 4c 49 51 52 4e 4b 48 4c 58 6f 74 74 67 52 41 23 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0d 0b 14 29 32 40 4c 5a 61 72 82 88 84 60 59 53 56 57 54 55 5f 5a 65 66 61 64 66 64 6a 65 6d 70 6a 74 6d 72 72 6d 77 7a 70 79 82 7a 7c 7d 81
 81 84 87 86 88 85 82 88 8f 92 90 8d 8e 8f 8e 8e 8c 92 91 95 96 97 9b 97 97 9e 99 95 9f 9a 9c a0 a4 a8 a8 aa a0 a6 a9 a2 af a6 a7 a8 a3 a5 a5 9c a8 9d a2 aa a2 a6 ab a9 b1 bb bc c8 d6 dc e2 e4 e7 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff dc ca cd df e0 e9 ec ef f2 fe ff ff ff ff ff ff ff ff ff ff ff ff ff f6 e4 d8 d6 cd cc c2 c1 c1 b4 ba b7 b0 b9 b0 ae aa ab ae a8 ab a4 ad 9e a8 a6 a6 aa aa a7 aa aa ac a7 9e a3 96 a2 a7 a3 9b a1 9c 9c 94 9f 93 94 92 94 8c 93 94 89 93 8b 86 8b 84 7b 82 7d 7c 7c 84 7c 76 78 7e 7b 7a 78 7b 74 73 67 6c 67 67 68 5f 63 64 61 63 5b 58 59 51 53 59 52 52 51 59 4d 48 4c 48 51 50 59 72 76 6f 67 54 37 2a 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 0c 15 21 29 3d 4d 5d 66 7f 82 88 7c 68 56 4d 58 59 54 59 50 55 59 67 61 64 70 61 63 66 66 6e 6a 68 71 6e 6e 77 75 76 72 6d 77 74 7b 7b 7f 79 77 7c 80 83 83 83 84 78 83 82 8d 80 8a 91 8b 8e 8d 8a 93 90 90 96 95 99 90 9b 99 9b 9e 9f 9e ac 9c 9d a0 a1 9f a7 ad a8 ae a5 a4 a4 ac 9f a7 a9 a7 9c a5 a2 aa a1 b2 b0 b0 b6 c2 c5 e0 db e5 ee f0 ff ff ff f8 f9 f6 ff ff ff ff ff ff fe ff fd dd cd c0 c1 d1 d2 e2 e8 f3 f0 f2 ff ff ff ff ff ff ff ff ff ff ff ff ed e2 db d7 d2 c4 c3 be b8 b8 b6 b7 ad ae a6 a7 aa a5 a7 a8 9e a1 a1 a2 a4 a1 9a a0 a0 a4 a5 9b a3 9f a8 a1 98 92 9a 99 9c 9c 97 9e 90 90 8c 97 97 8d 8b 84 89 8c 8b 8d 88 86 89 7a 7c 74 80 7e 7b 81 77 7f 79 70 77 6e 71 75 74 70 70 68 66 65 5f 59 64 5c 61 58 61 59 5d 50 54 4e 51 59 50 53 48 4a 4b 49 44 41 5e 69 7e 78 66 50 34 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 0f 1c 2f 3a 4d 50 61 6c 73 7f 85 8d 72 64 54 5a 5a 5a 51 54 58 5f 5f 6d 62 65 62 6d 69 72 6b 71 72 73 71 6f 6f 6d 7b 75 71 7b 75 7d 7c 7a 84 80 7a 7f 81 82 83 86 83 8b 83 86 87 87 8e 8a 92 8e 84 92 8e 8d 92 94 99 96 90 9e 9c 9f 9e 9e a4 9a a0 a4 a8 a0 a8 a6 a7 af 9f a4 a3 9e ac a9 a6 ac a5 a6 a0 a3 a5 aa a9 af b9 b0 bb c5 ce d7 e7 f8 ff ff ff fb f7 f9 ff ff ff ff ff ff fd ea cb 97 ba b4 b2 c1 d0 cf df eb f6 f5 f6 ff ff ff ff ff ff ff ff ff ff e3 e2 dc cf ce c3 c3 be bb ba ac ae a8 aa a4 ab aa a4 a8 a0 98 aa 9a a1 a2 a3 a5 95 9d a0 98 9a 9e a1 a0 9b a0 97 98 98 99 a6 9b 95 99 8d 90 92 95 8e 93 91 8b 8a 8a 8a 84 81 7b 80 80 7c 7b 7d 7b 77 76 77 76 7b 77 7a 71 70 6e 6e 70 6c 68 63 63 62 61 60 65 65 5f 65 5d 57 51 55 54 53 50 4c 50 4b 4e 50 48 4c 4c 53 65 77 75 61 51 2f 1f 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 12 14 25 2a 38 4d 54 5c 6b 77 86 89 95 75 5d 5e 52 53 54 50 5c 55 59 5b 5f 6d 63 62 6d 75 73 7a 74 75 7b 6f 70 71 74 77 71 79 7c 71 7b 80 78
 83 7f 80 7d 82 7e 81 82 7c 8b 7e 81 86 90 8b 8e 87 8e 85 8b 8a 90 92 94 98 90 92 9a 92 91 9d a4 95 9f a0 a5 a4 a4 a2 a4 af 9f a7 a5 a3 a7 a4 a4 aa aa 9e 9a a1 9c 99 a4 a2 a1 ab a6 b4 be c5 d8 df fd ff ff ff ff ff f3 ff ff ff ff ff ff e9 cb b6 7d aa aa b1 af ba c4 cb d6 e0 f6 fb ff ff ff ff ff ff ff ff ff f2 df cc c7 bf bc bc bc ba b4 aa b4 a9 af ad a9 a4 ad a3 ab a6 a2 9c a0 9a a0 a0 9a 95 94 9c 9b 97 95 99 98 99 98 93 98 94 99 9a 8f 95 94 86 8d 8f 8d 8f 8e 87 8d 8b 89 88 86 86 82 7f 7e 76 75 7e 72 72 72 77 84 75 6f 73 75 74 71 6b 6d 6a 60 5f 68 63 5f 63 60 5e 5f 5b 5b 5e 5c 56 52 56 53 53 47 52 40 50 44 47 48 54 5f 71 6d 67 54 35 21 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 06 11 1c 29 3a 4d 5d 63 6f 7b 84 8f 8a 81 5e 5b 4e 55 5a 50 58 53 54 60 5d 67 64 64 66 6a 77 7c 7a 7b 75 73 72 69 6e 69 70 74 70 74 6b 7a 72 7c 7e 85 7b 77 79 80 80 86 87 80 84 8a 82 87 87 83 87 85 84 80 8e 8b 93 92 8f 92 93 8c 91 9a 97 9f 9c 9a a4 a0 a0 a2 a2 9f a7 a1 a4 a3 a6 a5 a9 a6 a0 9a 9a 91 92 99 98 9b 8f a1 a5 a7 b2 b1 be d2 fc ff ff ff ff ff f7 fd ff ff ff ff e9 ca b5 a4 9d a1 a0 a3 a6 b1 bb c8 d5 d6 e8 ff ff ff ff ff ff ff ff ff f0 d6 ca c1 c1 b1 b6 ab b4 b5 b3 a8 aa a3 a5 a7 a4 9d 9c a7 9f a0 a3 98 98 9a 92 96 98 91 97 9e 98 93 93 91 8e 91 90 92 8e 92 94 8b 92 89 89 8c 8c 81 89 83 87 89 88 7d 79 76 88 7b 7d 82 72 73 72 73 78 77 78 79 78 68 6a 6d 67 73 6b 68 75 62 64 67 5e 5f 62 5e 61 65 5e 6a 5b 5f 5d 57 60 4c 4f 55 4c 44 43 4e 45 4f 4d 4f 61 78 66 65 58 3a 1b 08 07 03 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 15 1b 34 44 50 54 62 70 7b 82 8e 96 85 64 52 51 4e 54 5a 54 56 54 5e 5b 60 64 66 65 6d 6b 77 78 78 7d 6f 74 71 72 76 73 76 76 71 73 77 78 77 75 77 7b 77 82 7f 81 7a 78 7e 7b 7e 82 82 7b 80 81 89 8d 85 89 8f 86 98 8e 93 95 93 92 8e 98 94 98 a1 9b a2 9f 9b a2 a3 a1 a9 a5 a7 9f a2 a3 a0 94 96 93 8e 8c 8b 83 88 94 8f 93 94 9e ab b1 b5 ea ff ff ff ff ff ff ef ef f2 ff f0 d6 c1 b1 a1 9c a3 a6 b2 ae ad b6 c4 ca d0 e4 f5 ff ff ff ff ff ff ff fd df c3 bf b9 b8 ac b1 ae ab a7 a4 ad aa a2 a1 9f a2 a0 a7 a0 9c 92 a0 a2 94 97 98 93 90 8a 92 8a 94 92 90 91 8b 8d 8f 90 81 86 8f 89 84 8d 84 7f 85 8b 7e 89 8c 82 7e 79 7f 86 76 77 71 73 73 74 75 77 75 6c 71 76 77 75 6b 77 66 71 6b 71 69 64 67 66 6d 66 68 5a 5c 60 65 64 5c 5b 54 5e 54 51 56 4a 51 4e 49 4c 44 4d 51 52 60 69 67 68 53 35 22 09 05 0d 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 08 0f 10 21 2f 48 52 64 66 6d 7d 8e 8f 96 89 67 4d 57 54 57 59 58 5f 57 55 60 5e 60 60 65 71 78 7b 76 7d 7d 75 78 72 75 70 72 7b 74 7c 6f 75 79
 76 78 7a 79 81 71 7d 75 7b 7a 7d 7d 79 81 75 81 7f 82 8e 82 87 91 92 87 8e 8f 8d 8e 93 9b 8f 99 99 99 97 a3 9c 9e a3 a2 a5 a0 a5 a1 a1 a0 a2 9d 9f 8e 93 8b 87 8e 89 92 8e 8b 8d 8c 81 8a 96 9f a5 d3 ff ff ff ff ff ff f1 da d2 d4 cf be ab b1 ac a6 ac b4 b2 b2 b5 b5 b9 bb bd db ed f8 ff ff ff fe fe ff eb cb be c1 b6 b5 ab b3 b0 aa ad aa a9 a8 9f 9c a6 a7 a0 a2 9a 9d 9a 9c 9c 99 96 94 99 8f 95 8f 91 8f 91 8d 8c 8d 8c 87 88 89 87 8b 8b 8f 88 8b 84 7f 88 7e 85 7f 76 7b 76 84 80 7f 7c 75 76 73 73 6d 71 75 65 7b 6e 71 73 70 67 6f 6d 73 6a 6c 65 69 5e 5a 5c 62 61 62 5f 5a 66 57 59 55 54 54 53 4e 55 54 51 4a 40 4c 4e 4e 50 5b 6e 6a 64 4c 33 27 12 08 07 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 06 23 30 46 4e 5b 66 6b 7b 89 8f 92 88 5c 4e 54 4b 51 52 52 55 59 55 54 57 54 51 58 66 72 7e 76 78 76 75 77 74 74 73 6d 77 74 6b 77 71 72 75 78 7f 77 70 78 74 79 83 78 80 7d 77 75 77 82 79 81 7e 83 7d 8a 8d 86 8b 86 8e 8f 98 8f 8a 94 99 97 9a 97 9f 92 8f 9f 9b 9b a2 a1 9f 98 9e 99 8f 8f 89 88 7a 89 80 76 7f 7e 82 7b 87 89 8f 91 9f bf ff ff ff ff ff ff f6 d1 ba b7 ac ad aa a7 ae ae ae b1 ae a5 a9 ae b4 b4 c5 cc d3 e4 eb f5 f1 eb f2 f4 e0 ce ca c0 b8 b8 b3 b5 ae a8 a7 a5 9f a7 a3 9e 9f 96 9e a0 a2 9a 97 9b 98 94 96 96 96 93 93 87 8b 90 8e 89 7e 85 85 7b 7b 83 7c 83 83 7f 7a 83 77 7c 7e 78 7c 7b 7c 78 78 73 80 71 76 76 6d 6c 6e 71 6d 65 6e 6b 77 73 68 72 65 73 70 6b 74 64 60 61 61 64 61 60 66 65 62 5e 59 60 5b 58 53 54 51 4f 50 4b 4d 45 4f 49 44 49 47 57 6e 6c 5f 4e 37 28 1e 0e 03 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 08 16 2d 43 56 5e 6d 73 85 8b 96 97 8c 6b 52 56 4e 54 57 59 5a 55 57 59 54 62 56 5a 64 65 6e 6e 7b 78 74 7b 80 82 7e 77 7b 76 73 77 77 71 75 74 75 70 7b 7a 73 73 76 79 7a 79 73 77 76 7c 7b 7c 81 84 82 87 8e 8e 88 86 8b 90 87 8a 91 97 9a 99 9b 9d 96 97 92 9f 9a 9a 94 9a 93 99 96 91 93 83 83 86 80 7c 77 80 7b 80 82 83 80 7e 83 83 91 a1 de ff ff ff ff ff ee bf 9f a1 9e a0 a3 a8 a5 a1 9a 94 93 89 96 97 9c a9 aa b5 c3 d1 d2 d7 e0 de e6 e6 e1 cf c4 c4 bc bd b6 b7 ab b5 ae aa a4 a1 a1 a8 9d 9e 98 9c 99 9b 97 98 98 94 95 95 8d 91 89 85 88 86 85 89 7e 7e 86 7f 80 7f 82 84 88 78 7a 82 74 6f 77 77 7a 76 72 75 69 75 6d 75 71 6c 73 6d 68 6a 6d 6b 6d 6a 69 6d 6f 6f 71 6f 77 6f 6e 65 63 5f 5f 5e 61 66 60 64 5d 59 62 5f 5d 53 5e 4f 47 52 49 52 4b 4b 4d 54 51 4c 53 5a 6f 66 5a 54 3c 31 25 14 0f 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 13 14 28 44 58 66 6c 7a 79 84 9c 9a 84 69 5a 4c 58 51 56 5a 5b 57 5a 5c 55 56 5c 5e 63 69 68 66 77 72 72 6e 7b 80 81 81 80 80 75 6f 76 75
 71 79 75 71 78 6f 76 7e 73 7b 7b 75 78 7b 83 81 7f 78 85 83 86 80 81 86 86 86 8d 8a 83 90 87 94 95 8d 95 94 8e 91 8f 92 92 91 90 95 97 92 87 84 87 87 84 7d 79 75 78 72 7b 7b 7b 7f 79 83 80 86 8e 94 c4 ff ff ff ff ff e8 b2 97 98 95 9e 9e 8e 88 86 7c 75 79 75 7b 75 8a 86 95 9a a3 b2 b2 c2 ce d4 e1 e0 e2 d4 c0 c3 b9 bd b6 c2 b2 b9 b7 a6 b1 a7 a9 a2 a3 9f 98 9f 95 8f 94 98 8f 90 8a 8b 84 8a 89 82 7c 83 84 8a 7d 7e 77 7c 7a 79 81 7b 84 73 73 74 6c 78 6c 6d 6d 73 75 6e 6c 74 6e 71 6c 6d 6b 72 62 6d 6d 71 6b 6f 69 70 67 6e 74 71 68 67 6d 73 68 65 62 63 68 65 61 61 69 5f 65 58 55 53 54 5e 4f 51 49 56 53 4f 50 51 54 4c 5a 59 68 6e 61 4d 43 35 25 20 07 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 00 06 09 26 3a 5d 5e 6c 78 80 88 98 98 7f 65 54 5b 57 57 52 59 56 55 5b 58 50 59 59 5a 60 66 67 5f 68 6e 73 75 77 79 70 70 80 77 78 77 71 6d 74 6c 7c 6c 74 74 7b 76 6e 74 6f 73 7b 79 79 80 79 78 86 81 85 7f 86 7d 83 89 8e 84 89 89 8d 99 94 96 88 98 92 8c 87 8c 8d 90 8a 90 85 90 89 8e 87 81 83 81 77 71 78 79 76 77 77 7b 78 80 7b 7a 8a 8e a7 f4 ff ff ff ff d2 aa 90 8f 99 8c 85 7d 6e 63 62 60 62 6e 6d 70 75 65 7f 89 91 9a ad b3 c0 c6 ca dd dc cc cd c1 c1 ca bd c7 c0 b4 b6 ba b2 b4 a8 aa 9c 9f a2 9a 94 93 8c 94 8c 90 88 89 86 83 80 80 81 7d 76 75 7e 75 79 78 73 75 7c 72 71 71 73 77 6b 6f 75 70 6d 6f 6e 6a 6f 6b 66 6e 6c 70 6d 69 68 66 69 61 66 6a 69 72 68 6c 65 6d 63 67 6e 64 62 65 61 63 61 61 60 67 61 5a 5e 5c 58 53 55 53 53 50 50 52 4d 4c 50 46 50 4f 53 5e 67 68 5c 51 41 36 2b 1e 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 03 08 10 1d 32 4b 61 66 81 8c 91 96 8f 7e 61 55 50 4d 58 4d 56 5c 5a 5c 60 55 59 50 56 59 5d 61 62 64 69 6c 6c 73 6f 72 78 6f 79 74 74 72 72 6d 70 74 6f 74 80 79 79 77 7a 75 71 7b 7a 7d 7f 74 81 79 84 77 84 88 87 90 8a 80 84 84 8b 84 82 8e 92 8a 84 83 85 8c 84 91 8f 89 87 89 86 86 84 88 83 7b 72 75 74 74 77 74 72 75 78 78 75 81 83 7e 86 9b df ff ff ff ff c5 a0 8f 8a 80 72 5d 64 59 5b 5e 5d 69 66 69 6c 71 78 7d 81 88 91 9d a8 a8 b4 c4 ca d9 d5 d4 d4 cd ce c8 cb c8 c6 c1 c2 b9 b6 b8 b2 98 9f 9e 96 97 8f 8c 87 8b 80 82 84 81 7f 7d 7e 7f 7b 7a 76 75 7b 75 73 70 76 79 75 73 71 6c 67 66 6f 68 69 67 61 6b 6f 69 6c 6b 6d 65 66 62 6b 62 66 6f 6c 64 61 61 6c 6d 74 6c 6a 67 6a 67 67 63 5d 66 64 66 5e 65 63 5e 60 59 5c 4e 57 55 52 53 4e 56 4d 54 45 51 4d 4c 52 48 56 60 67 61 56 3f 39 31 23 12 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 08 0c 1a 31 4d 5d 67 72 85 90 96 94 88 6c 57 4e 57 55 56 5c 56 64 57 5d 5b 5a 5d 5e 5e 5b 60 65 67 6a 63 6a 69 72 73 79 7c 7f 79 76 6f 6f
 75 73 70 78 6c 72 7d 76 77 74 74 78 77 78 77 7b 80 7a 82 81 7e 82 8c 87 89 84 82 82 8e 84 85 87 8b 88 8a 91 8f 83 86 83 8e 86 88 84 83 85 7c 7f 88 77 7f 75 79 6d 79 7c 6c 6e 70 75 7c 81 76 7e 7b 88 93 c2 fd ff ff ef b2 96 85 6e 62 5a 55 5a 4f 4f 5d 5e 65 6f 69 73 74 78 7c 80 89 94 94 a3 ab b0 bf cb dd dd d8 dc dc e1 dd dd d6 dd d7 d1 cf b9 b6 b3 b5 a0 a6 9a 9c 94 88 8b 8e 88 82 8a 7c 82 84 7c 77 73 79 6f 71 6d 71 6b 73 71 73 6f 6c 70 74 71 6f 64 69 62 6b 67 5f 6c 69 69 5e 65 67 6b 6a 66 61 6c 67 61 66 69 6f 75 68 6e 71 6a 79 68 6d 67 62 69 68 63 6b 63 61 64 68 64 64 56 52 5b 5b 52 50 52 4f 4b 55 51 50 55 51 57 59 58 6b 6b 62 57 48 49 36 24 14 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 0a 06 08 12 30 45 53 6b 75 79 92 8b 95 85 62 55 59 59 54 5b 56 54 5d 5e 56 59 5b 51 5b 5e 61 60 63 62 67 66 71 6e 76 70 6a 75 76 73 73 6d 6f 74 74 76 72 6d 71 71 77 74 78 7c 76 71 7b 73 7a 80 7d 81 78 7f 7a 83 7b 87 82 80 88 7a 82 84 86 87 87 81 80 85 7e 87 8a 8c 8c 86 84 86 81 7f 81 7e 75 76 73 71 74 71 75 70 73 78 7c 73 76 75 7d 80 8c 95 b5 f3 fb ff db a4 85 6a 51 4d 51 4c 4e 53 59 60 66 67 66 6f 74 7a 74 84 84 90 95 a2 a5 9f aa b9 d1 d3 e9 e6 ea e9 f6 ed f2 eb e9 e2 d7 d6 d3 ca c3 b3 ab a6 9e 99 8a 89 86 80 81 75 85 79 7e 7d 75 7b 7b 76 76 6c 73 71 6e 67 69 6e 6e 6d 69 6e 6b 6b 65 69 62 5a 5f 62 6b 5d 61 5f 62 5e 5f 66 63 61 61 62 65 67 69 65 6a 6b 64 6d 6a 71 64 61 6c 5d 62 68 66 62 61 62 62 59 59 5b 59 59 51 57 4c 4d 53 50 4e 56 4e 55 4b 4f 52 52 57 5f 6a 5b 59 49 4d 3e 29 1f 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0b 14 19 27 36 52 69 75 7b 81 89 92 7e 62 60 58 5a 54 50 5d 5b 5e 5f 5a 63 51 59 60 5e 5f 5e 60 60 5e 5e 69 6f 77 73 76 7a 79 6e 78 72 74 72 6c 73 6f 6d 6d 65 76 77 71 6b 75 71 71 77 74 7a 77 79 7d 7b 80 7e 86 88 89 79 85 81 7f 86 84 7f 81 80 89 84 87 82 84 8d 81 89 82 7b 89 84 87 7b 78 74 75 77 73 6c 7b 71 75 71 80 7f 80 84 7a 89 89 88 af d1 f1 ef c8 89 6f 4d 48 47 4e 51 52 52 5a 56 60 6a 64 6f 77 76 81 88 8b 95 a2 a8 ac af bb c4 d0 e5 f4 fb ff fe ff fc ff f6 f8 e9 e3 e0 e3 d6 cc ba b3 ac a6 9e 8d 88 85 87 82 7f 7f 79 75 79 72 73 6c 6d 6c 6d 6a 63 70 6b 65 69 5c 6b 62 67 64 69 6a 68 5e 55 69 61 62 5c 61 65 62 66 5a 67 64 61 62 5f 64 62 64 67 64 62 6e 6b 67 6e 69 6f 66 69 66 6a 61 69 5f 63 5f 58 5c 54 50 4f 4f 52 56 54 50 4d 52 52 57 52 4f 4d 4e 51 59 6e 71 65 5d 47 46 36 25 18 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 05 11 10 15 26 35 50 5b 67 7e 84 8a 90 7e 64 56 51 63 59 57 5e 54 5d 5b 66 64 5f 5d 5a 53 5c 59 5f 61 5d 6c 68 70 74 7b 72 75 78 70 74 6b 72
 6e 6b 6b 71 6e 72 79 70 6d 75 75 74 74 70 73 78 71 6b 74 7e 77 7d 85 75 81 7d 84 7e 82 78 7e 85 80 82 86 80 7e 83 82 8e 8c 84 87 89 84 95 87 8a 86 77 76 78 6c 72 6e 70 6b 78 7a 76 7a 7c 79 7d 7d 88 93 98 c9 ee e3 af 7f 57 49 45 46 4f 4e 4d 54 5f 5f 65 6c 77 79 7c 7e 80 96 a8 aa b4 b8 b9 bf c3 d5 db ed fe ff ff ff ff ff ff ff ff fe f4 eb ea e1 da c2 b6 a8 a5 99 95 91 7c 84 84 7d 81 75 75 6c 70 74 76 70 6c 66 67 6d 67 67 66 6b 6b 71 5f 6a 6e 63 67 64 68 62 62 65 66 5e 64 61 63 66 60 66 5f 5a 5f 69 69 63 65 5f 6b 6a 6b 6c 69 6f 67 67 70 65 64 63 61 67 5f 5e 56 58 4e 5e 53 58 51 5a 50 4e 56 58 4e 55 51 4f 53 4f 57 58 5c 6a 6d 75 62 59 4d 34 30 1b 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 10 0a 1b 14 26 33 45 58 5d 74 88 7d 8b 85 6a 58 54 55 5d 59 5c 5d 56 5b 5d 5a 54 58 5d 57 62 55 55 63 5e 5d 6b 71 79 80 7a 76 74 70 68 6d 76 72 75 72 69 6f 73 76 6a 7f 73 68 72 73 70 75 79 6c 71 75 7a 78 7b 7f 7d 81 7a 78 7e 7d 80 84 84 86 83 7c 86 84 87 82 83 8a 90 85 8d 94 93 88 8a 84 79 7b 73 74 76 6b 74 75 6f 77 77 7d 7d 82 85 8a 85 81 94 ad dd d8 9e 60 4f 42 46 43 4f 44 55 5a 5b 66 6c 70 70 77 7f 8d 98 a8 b7 c0 bf cc d1 d6 d8 dd f2 fc ff ff ff ff ff ff ff ff ff ff ff fa f9 ea d7 cb bc a5 a5 9a 97 8c 8a 7d 77 84 7d 7d 79 73 73 72 68 6a 60 65 5f 60 67 64 6a 6b 63 68 62 6d 66 5a 5d 68 65 64 62 5a 64 67 5a 60 6a 68 67 63 62 61 65 63 68 6a 5f 6a 6a 6a 6f 71 6c 6c 6c 6f 6a 6a 6e 6d 5e 62 67 5a 64 60 54 5e 5d 53 56 4b 58 50 56 56 56 5b 56 54 50 47 50 51 5b 68 73 6d 65 5a 50 38 34 18 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 11 13 10 16 24 2e 35 40 5f 72 79 8b 89 81 66 52 4f 4e 5a 58 61 57 5e 5e 50 5f 5e 59 5f 51 62 56 59 57 63 68 6b 77 77 6d 6f 6a 6c 64 65 6b 65 6b 6f 66 6f 73 6d 69 6a 6c 6f 69 6d 6b 6c 6a 69 68 74 6d 75 75 79 80 7d 80 7a 7a 7d 7b 80 87 85 87 81 81 84 74 7f 82 80 80 80 78 86 89 8f 89 8c 85 80 79 77 6b 6b 74 75 7f 75 77 73 7c 7e 7b 74 77 7a 7b 84 9c d3 cc 84 52 3d 3c 3a 3f 41 47 51 59 5c 65 70 78 7d 89 8e a0 b4 b9 d4 cd d1 dd e1 ef f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f0 e8 d4 c4 b9 a5 95 93 90 88 7f 81 7c 7e 7a 7b 77 76 6e 70 6a 65 69 61 5f 65 63 60 62 64 6e 5e 69 67 60 5e 63 63 61 63 5a 5c 61 60 67 6b 62 61 67 6a 68 66 69 63 61 65 65 67 63 6b 6b 69 6e 5e 67 70 6b 65 63 60 6a 5b 61 66 59 59 56 56 4b 57 50 4b 56 51 54 50 4f 5b 51 58 4b 50 52 5a 77 70 6e 66 54 50 3e 26 1d 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 09 0d 18 1a 22 29 29 32 40 46 5a 6c 77 84 7a 62 58 5f 56 57 51 63 5b 68 5b 5e 61 53 5a 56 58 5b 5a 5c 5e 63 63 6b 79 71 70 70 69 60 69 61 6c 68
 69 6d 69 69 72 74 6a 74 6a 65 6e 6c 69 69 68 68 62 6a 72 66 71 7b 7a 78 76 7c 80 85 8b 8d 8a 89 80 85 7e 79 77 78 77 77 7b 80 7a 82 88 85 7e 87 87 7d 7a 7b 6b 73 74 6d 71 69 76 76 79 75 73 72 75 71 76 90 8f b1 b9 71 4d 3f 3c 43 3f 47 49 4d 5c 5e 69 74 86 8e 9b a3 bb d1 d6 e0 df ef f4 f5 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 ee d8 d0 b6 a9 9c 93 8b 89 7e 80 7a 7c 7c 7c 77 74 72 6a 72 65 6c 62 5d 63 62 61 69 64 6c 61 5f 6e 68 60 5d 5f 63 5d 6a 65 5b 5f 64 72 65 6d 6d 65 66 6b 6b 64 68 6d 6f 6a 69 65 6c 71 69 76 67 6f 6c 62 67 5d 69 65 67 5f 59 58 5e 4f 57 53 5b 55 4d 59 5a 4f 53 51 4e 55 50 51 57 5a 67 73 6f 61 53 56 42 30 16 06 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 0f 14 11 16 28 28 2b 32 33 38 47 60 6e 73 66 5b 4f 51 60 59 5d 5a 56 60 63 5f 61 4f 50 5d 55 5b 58 56 61 63 6a 71 6e 6b 72 62 69 62 59 60 66 65 64 6c 6b 6c 6f 64 66 6e 75 6e 6a 6b 68 60 65 65 61 6a 66 74 6c 6f 76 71 7c 77 85 84 82 90 8b 87 85 77 76 7b 76 7e 7a 7a 7e 78 76 82 79 85 83 7c 79 76 76 7f 72 73 76 6f 6d 6f 74 74 74 71 6c 76 70 70 79 83 82 9b 99 6c 4e 38 3c 3e 3e 48 51 59 5a 66 74 85 8e 9e aa c0 d4 e6 f4 f1 fa f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 e2 d1 c4 ac a0 94 8b 8d 7d 83 82 7b 74 7b 74 6b 72 6a 6e 67 62 64 66 65 6a 64 69 61 67 64 64 65 5e 60 64 64 5d 5f 61 62 63 65 68 67 62 60 66 66 66 64 61 69 66 6f 6a 6c 69 75 67 72 6d 69 6e 6d 6b 67 67 63 63 64 5a 61 5c 57 5f 4d 51 52 50 54 57 55 58 58 54 54 4d 53 55 55 52 6a 79 7b 74 6b 57 55 44 2f 18 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 16 1c 21 1d 2f 2c 29 33 3a 4a 4c 52 5b 59 5a 57 56 54 5c 53 5a 5c 53 66 5f 56 58 52 5b 5d 5e 5e 5c 67 64 62 64 6f 75 5f 66 63 61 53 5c 69 65 63 6b 6d 66 68 6c 6d 62 6e 6b 65 64 65 65 65 5f 62 5f 68 68 68 70 67 74 78 81 84 84 7c 79 80 7f 7f 78 72 7b 72 6f 7d 77 74 77 72 75 7d 71 7f 83 80 7c 7b 7a 76 77 73 72 6b 71 75 77 75 70 6c 65 6d 71 77 77 7a 8a 80 57 3d 35 2d 3a 42 42 53 5f 65 6b 7a 8c 9b ab c1 d6 e3 f0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e8 d9 bc aa 9f 90 8b 84 81 82 7c 81 72 75 6e 6b 68 6f 61 63 63 60 5b 58 5d 5d 5c 68 5c 62 61 68 5d 61 64 57 5a 5f 59 61 5d 5e 61 5f 5d 5d 60 57 57 61 61 67 70 68 6c 6f 6a 72 68 6d 6d 74 6d 6c 65 66 68 65 65 68 65 57 59 5c 58 59 5b 59 54 56 53 57 5e 55 52 50 56 4d 50 56 56 61 6f 7e 74 6a 5c 58 3c 2c 12 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 17 25 28 25 2f 2a 29 31 32 3a 42 47 4f 52 58 5b 52 56 53 47 50 53 57 60 5a 59 58 55 57 55 5b 5f 5e 66 5f 5d 61 65 65 5d 5f 54 64 5f 60 6d 5b
 60 65 64 5f 70 61 6d 6c 6c 78 61 65 6e 67 65 5a 5e 63 62 64 64 61 6c 65 71 7a 82 86 7e 85 7f 78 7d 74 76 76 72 72 77 6f 7c 79 79 7b 7d 79 75 75 79 80 7d 7a 77 6f 70 75 73 70 81 6e 6f 6c 68 6c 7a 74 75 74 86 81 78 4d 40 2e 35 39 43 50 56 5e 6a 73 90 a6 b3 c4 d6 ea ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f5 d7 c0 b3 a0 9e 8d 88 89 78 76 79 78 6c 72 6e 6a 67 64 66 69 63 62 5d 63 61 5a 63 5f 61 69 64 63 5c 5f 66 61 5a 5c 5d 5d 5e 64 56 64 5a 55 58 53 5c 5c 65 63 68 64 64 65 64 70 68 72 6e 70 7b 6e 6f 6a 5d 69 61 65 5f 5e 60 58 5c 57 52 5a 59 57 58 58 56 54 51 50 52 4d 51 61 65 7b 80 77 65 58 59 3e 21 11 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 1d 25 2b 26 26 2b 36 32 30 3e 40 48 49 53 50 54 52 56 50 53 54 55 4c 59 55 5f 5e 52 58 57 58 5e 58 54 5d 62 5c 69 64 67 5f 5b 62 5b 5a 61 5f 62 65 63 63 60 67 60 64 6a 69 6e 69 65 63 60 5c 60 63 67 5e 5f 61 5d 69 6c 72 7a 79 7b 76 7b 77 76 74 75 74 6d 70 76 75 79 6f 7e 79 72 78 78 74 7c 6c 7e 74 84 78 74 72 76 73 71 6d 70 71 6f 75 74 7b 78 7a 7b 7d 67 3b 2f 31 30 3c 46 4c 5b 64 77 83 98 ae c9 cd ef f8 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f4 df ca ae a6 9d 89 88 7e 84 7b 7b 75 70 76 70 69 6b 67 66 60 5e 64 5e 66 60 5c 63 64 5f 62 68 58 56 62 5c 59 5f 5a 5b 61 5e 5b 66 62 5d 5e 5c 5b 54 5e 61 5d 67 64 60 6b 74 67 71 6f 78 6b 6e 6b 70 73 66 64 62 6c 65 5b 59 59 59 5c 57 59 4e 52 59 54 57 58 61 52 59 57 56 60 6d 7d 78 7c 6b 5c 56 3e 27 14 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 17 20 2d 30 27 33 28 32 3d 3d 42 4f 44 47 46 4d 51 4b 46 52 50 52 56 56 55 53 5d 51 4a 57 56 54 5e 5a 57 5a 5d 5b 5d 5c 5e 5f 63 61 55 5b 64 5f 5d 5e 61 5d 64 60 69 62 66 6d 6c 67 63 65 5c 62 5c 59 5e 5d 66 61 5d 6a 6a 6a 6d 6c 78 79 78 70 69 6a 6b 71 6f 6b 6d 78 69 73 74 6c 75 73 76 7d 79 75 7b 72 6f 74 72 71 6d 72 6a 6a 66 67 68 68 71 74 77 7b 7a 62 42 35 2d 32 37 46 44 61 69 7c 87 9e b9 d3 df fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa e0 c6 b9 a1 91 86 7e 80 7f 78 7a 71 6d 6c 6b 65 61 66 64 5d 56 5f 62 5b 5f 64 59 61 5b 57 63 5b 63 62 5f 5d 5b 5c 61 55 65 5a 59 5d 59 5b 56 50 5a 56 62 5a 5f 64 6a 67 6b 67 69 70 73 75 70 70 72 6a 61 60 61 62 64 5b 5c 59 5a 54 59 57 51 53 54 55 54 53 5c 4e 53 50 4f 67 72 7d 7d 7a 6f 57 4a 3c 21 10 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 18 2d 2e 33 35 2d 2e 2c 30 3b 45 49 42 41 4a 50 4e 5c 51 52 55 4e 52 5f 53 57 54 50 4d 54 51 62 5c 56 58 59 5f 5a 62 59 5d 55 5b 57 63 63 5b
 5c 61 62 60 66 5a 65 5d 60 66 64 69 6e 61 5b 63 5f 5e 66 5f 6a 66 63 64 68 6a 67 6f 69 74 79 75 6c 6b 6c 6f 71 6e 6f 73 72 72 6f 71 72 6e 6f 6e 75 7f 78 72 6c 72 6b 6b 6a 6a 75 69 65 6d 62 60 60 6c 6b 6e 82 6f 66 40 2b 2b 35 46 45 4f 69 79 88 98 a9 c2 d5 e9 fe ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fa db c6 ab a2 9c 8c 87 83 7b 75 78 77 6c 73 6e 62 66 66 57 61 5f 63 56 5c 57 5b 5a 5e 5a 60 62 5f 5b 5d 5e 5b 5d 55 60 62 61 59 60 5c 62 5a 55 54 5b 58 54 5b 5f 5f 61 5e 6b 68 6e 72 74 73 76 70 6f 6a 6a 67 5e 66 65 61 5f 5d 56 5a 52 56 50 53 59 55 5a 58 53 53 52 52 56 61 7b 7c 79 75 65 57 4a 34 18 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 19 26 38 3c 3d 36 3b 30 36 44 4f 42 4b 43 4c 52 54 4e 4f 47 50 4d 51 59 53 55 59 57 4d 4d 56 57 56 52 57 52 59 67 5d 5a 64 62 64 5e 60 64 62 5a 5e 61 57 62 61 5b 5f 5c 5f 69 67 6f 66 66 64 69 60 5f 5e 55 61 65 61 65 64 61 66 66 60 65 69 64 5f 6c 70 6a 68 6f 6f 74 76 6d 74 70 79 6b 6f 76 74 7a 71 6c 6f 69 6d 73 65 6d 68 6a 66 65 65 71 6b 63 71 70 6d 5a 43 27 30 37 3e 4e 55 68 80 86 97 ac d0 e8 f4 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe de c6 b8 a3 96 87 81 81 80 82 74 73 72 6c 6e 5e 66 5f 61 62 5d 60 5f 57 58 5b 61 5e 5c 63 64 5e 61 61 64 5b 5b 66 5a 5f 59 5e 5a 62 62 5b 5d 5c 5b 63 5b 58 5f 63 5d 5f 65 65 6d 75 74 75 77 72 72 6e 6c 6b 67 69 6b 62 61 5f 58 57 57 58 5a 4e 54 58 50 51 4e 4a 48 55 5a 60 7c 80 70 70 63 53 49 2e 13 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 07 15 20 3b 46 3e 45 2d 30 3c 41 4e 4f 4b 4e 49 51 53 4b 53 4b 59 51 55 59 54 56 59 53 4e 54 51 52 58 57 50 52 55 5c 61 5d 60 61 62 5a 5f 63 5d 55 66 5c 55 5e 63 59 5f 64 63 5d 64 70 6e 62 5d 61 54 51 5c 5c 5c 5c 61 5f 5a 5d 62 60 63 63 5f 63 6b 65 6f 6d 6b 6b 71 6e 68 65 6c 71 69 72 6e 76 70 6c 5f 67 6e 65 68 6a 64 67 67 5c 65 6b 6e 5f 64 69 65 79 6a 59 3f 2f 34 35 39 51 57 6d 7d 8c a5 b7 d8 f2 fb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 e4 c9 b5 ae 9e 8a 84 7b 7d 7c 75 75 74 6c 64 6a 64 62 5d 57 60 53 58 58 53 5d 58 57 52 59 64 5e 60 61 52 55 59 5c 62 52 57 58 5c 52 64 53 59 52 54 60 5b 59 59 60 60 5d 61 5b 6c 6f 78 75 74 72 6e 6f 6c 66 61 66 67 61 60 59 59 57 59 54 59 4a 4d 51 4e 51 4a 51 4c 4f 59 66 84 81 7e 6e 62 4f 40 24 13 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 29 35 46 54 4c 45 45 44 4c 57 45 47 47 4f 4c 51 54 50 51 52 53 56 58 55 53 4c 52 59 5a 53 55 50 52 51 5b 5a 5c 5d 60 5f 63 5f 60 60 57 5e
 5b 57 5c 5b 57 5c 57 5b 5c 5e 65 66 6d 6b 61 60 5b 4f 52 5d 53 5c 59 4e 5e 50 5e 53 5e 5f 5c 5d 68 66 66 6b 61 67 74 69 68 73 6d 79 6b 70 6c 63 70 6a 6b 6d 6e 6e 6c 65 62 66 62 64 6a 5f 69 68 68 6a 69 6a 6f 6a 61 3f 30 2f 31 3d 4f 5c 72 88 9e 9f c3 d7 ef ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f7 d5 c8 b7 a3 92 91 93 81 83 6e 79 70 70 6a 65 6c 5b 5b 5a 59 5e 59 5d 56 55 51 5f 57 5d 5d 5d 5e 54 5a 5b 5b 62 54 5e 59 5f 5a 60 5c 53 5d 5a 55 5a 5f 59 5d 59 56 5e 57 66 68 6f 76 76 7c 6e 78 5f 62 6c 64 5b 68 5f 51 5f 62 51 56 55 54 53 4a 57 52 4f 4c 4e 47 4d 54 5f 6b 7f 82 7e 6e 64 4c 39 17 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 22 3a 45 58 57 54 5c 4d 5c 61 53 45 44 4d 49 56 4a 4f 52 4e 56 54 4f 54 54 55 4c 52 59 53 53 54 54 55 53 5a 5b 5b 5a 5e 60 5d 59 60 5f 5b 5c 5e 5d 56 60 61 65 59 5e 60 6a 6f 69 63 52 51 52 5f 5a 56 50 54 52 60 55 5a 60 56 59 61 5f 64 5f 66 6e 6c 6d 6f 70 6b 6e 6d 75 70 70 70 66 68 6e 63 66 65 69 6f 65 65 66 69 67 66 66 62 64 66 62 64 67 66 66 66 62 3e 37 33 33 42 4a 60 72 87 98 ac be e2 fd ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ea d5 bd af a5 96 8e 87 82 7f 78 80 72 6e 6d 61 64 65 5f 57 55 55 4f 55 54 5a 56 5d 5f 5a 5e 5b 59 5d 5d 54 5e 55 65 5a 59 60 59 5c 55 5a 5e 5c 5d 55 5e 5c 61 64 61 61 54 66 68 71 70 77 74 73 6c 66 66 68 64 66 62 62 60 62 64 59 59 51 57 51 4e 4d 47 4f 56 4f 56 55 4f 60 70 84 81 75 68 58 48 34 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 04 1f 3a 4b 55 68 69 6c 69 66 66 57 54 47 4b 45 55 52 59 49 53 51 56 5b 59 56 52 4f 52 56 57 58 53 55 59 59 52 59 57 5b 63 5d 61 5e 55 5a 58 56 55 5c 56 56 5e 54 5a 60 6a 6d 69 61 5c 5a 53 56 51 55 53 4d 55 55 5c 52 4b 56 54 56 50 5e 63 67 69 64 6b 69 75 61 72 6e 6a 69 6a 6a 6c 6c 6c 6e 68 6a 61 62 60 63 66 62 60 66 61 62 6c 62 5e 60 65 69 65 65 67 57 41 2f 39 3d 37 4d 56 6d 87 98 af c2 db fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e6 c9 b6 ac a1 96 92 8f 89 87 77 7f 70 76 71 5b 65 5e 5d 5c 59 54 50 55 52 52 56 4d 5d 59 60 5a 5b 5b 5a 5a 60 58 58 4f 53 5c 59 5b 57 5a 5a 56 52 53 56 5e 57 56 59 5a 60 5f 70 70 75 74 75 77 66 6b 69 62 62 61 5f 5d 61 5b 5c 53 52 4f 4f 52 52 50 4e 51 53 50 54 4b 54 62 77 82 7a 71 68 50 39 1f 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0b 13 34 4c 59 6f 67 6d 76 78 74 61 5b 47 4b 52 56 60 53 54 5a 49 52 5c 5d 56 5b 5b 57 4e 57 52 4e 61 53 56 50 54 58 5a 60 5b 60 62 5a 56 57
 54 60 5b 58 4e 58 55 51 5d 60 6a 6d 61 4c 59 53 4f 55 55 5b 52 52 57 53 53 5d 50 50 59 5b 59 5d 62 60 6b 6e 68 6f 6c 66 6d 68 6c 70 62 6e 66 6d 62 5d 68 69 5d 64 67 5d 63 64 69 67 5f 62 5e 5d 63 5f 61 64 5c 64 60 45 32 31 35 3c 48 55 6d 85 96 ad ca db f7 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fb e2 d2 b4 ad 9b 9d 89 8e 7f 89 7b 7c 6f 73 72 64 6b 60 59 5e 4b 56 58 52 59 4d 5a 56 57 59 61 5a 5a 58 5b 5d 5b 5b 52 57 55 59 59 65 56 4e 52 56 56 5a 52 54 5b 5b 5d 5c 5b 66 69 6b 76 77 6b 69 62 63 61 62 5d 66 5b 58 5b 56 53 54 51 4f 44 50 49 53 4d 50 52 4f 4c 4e 52 6b 75 84 7d 6e 5c 44 2d 1c 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 11 28 42 5d 69 6b 72 74 80 87 76 6b 53 54 61 6e 60 56 52 4a 50 5d 68 6b 6c 59 62 56 54 55 58 61 64 60 5d 59 4b 5c 56 52 60 5c 5a 59 5c 61 56 60 59 54 59 5a 5e 5a 57 5f 68 62 59 60 53 54 4d 54 55 52 51 4e 54 4d 58 56 50 5c 58 58 5e 64 64 6c 64 66 64 6c 6a 71 74 6c 71 75 61 66 67 5c 65 66 69 61 62 5d 5e 63 66 5e 65 5a 68 5d 63 5e 61 65 64 68 67 64 5e 40 2d 31 35 46 4a 5c 6c 84 90 a7 cc e1 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 d7 c1 a9 a1 9d 94 8b 93 83 8d 81 7a 7a 74 6d 68 5c 61 58 58 4d 51 56 4e 50 58 4d 5d 61 59 5a 5f 59 5d 5e 56 57 5e 58 5a 5d 5b 55 54 57 5c 56 5a 51 54 56 5e 60 5d 61 5a 5e 65 6e 6f 70 76 64 70 63 60 66 5c 62 60 58 60 5a 5e 56 59 58 4f 4e 4d 50 50 4f 55 52 4f 51 57 55 6a 85 7f 78 69 53 2f 16 15 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 0f 22 39 54 58 65 7b 79 85 89 7d 78 5e 64 6a 6e 67 66 57 52 56 5c 67 79 7a 61 5a 57 53 65 67 65 69 67 66 5f 54 57 5a 4e 52 55 5e 5b 60 59 57 5a 5a 5d 55 55 57 5d 5b 65 65 62 5f 55 54 53 4f 56 52 51 50 4e 59 49 53 54 50 57 58 52 60 64 61 6a 6c 6a 63 6a 70 6e 6e 66 71 6f 73 6b 69 68 62 61 63 6d 64 69 64 67 62 5b 69 59 59 61 68 65 60 5d 60 5a 5e 65 60 45 31 36 37 41 4c 56 6f 87 8f a6 b8 d8 ee ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e9 d8 c5 b2 a6 93 90 88 86 87 7d 7c 7b 77 76 6e 63 62 59 54 53 5f 54 56 53 52 4f 51 4b 5b 56 54 64 4c 5d 57 54 5b 58 56 58 54 52 58 58 57 5a 5d 54 53 58 5f 59 56 5a 60 58 5e 6d 6a 67 6a 6f 65 60 5c 5e 64 58 60 5e 58 5c 54 59 53 55 58 4d 54 4f 46 55 50 5d 4f 50 4d 56 57 6d 85 83 74 5c 42 26 0e 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 0f 1b 35 4f 58 6a 68 6f 7d 84 79 77 69 62 5b 60 6a 59 4e 55 50 55 57 66 69 5e 5d 51 55 5c 5b 64 5e 6c 72 62 5d 53 54 58 54 55 5e 5b 5a 58
 5d 56 53 53 51 54 56 5a 55 60 5a 64 5a 52 51 55 4c 4c 51 50 52 4e 53 55 5b 56 4c 54 56 5c 5e 61 61 5e 5a 6e 6c 66 67 71 7e 63 78 68 60 69 62 6a 61 5e 65 63 5b 63 5f 5c 62 5b 5f 5b 59 58 50 59 5b 5d 56 5a 57 5f 56 45 36 32 32 3d 43 50 63 7b 8f 9e b2 c9 eb ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e4 c7 bf a9 a0 98 96 85 89 84 82 73 72 74 72 6a 63 5f 61 61 5c 52 4d 52 4e 4b 51 50 54 52 4f 53 57 52 56 5a 58 53 55 59 53 4e 57 57 53 58 51 52 5d 4c 4d 58 5a 60 59 50 5d 5b 65 64 6b 63 66 59 65 4f 5c 59 59 5a 5f 54 5c 51 55 57 54 50 4a 52 58 49 4e 4d 54 54 52 4c 54 5f 73 7f 7b 6d 50 34 1d 0c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 02 08 15 21 47 5b 68 66 71 78 82 7d 84 69 5b 58 60 56 59 4c 55 4d 58 54 56 5d 5d 4e 53 55 59 5e 58 56 58 67 6d 65 5f 52 50 4e 54 57 5a 5b 5c 57 5e 4c 57 5a 4f 5c 56 5a 5a 5c 5f 57 55 5c 55 4b 51 4e 4e 4c 4c 4d 52 51 54 5c 56 58 56 51 5d 61 63 6b 6a 67 66 6a 68 76 75 6d 69 63 6f 6e 69 68 66 5f 6a 66 59 61 61 57 58 58 57 4d 56 54 5b 52 51 58 57 57 5f 5b 46 2f 37 31 42 4b 4b 5a 73 84 90 ab c2 d9 f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 df c6 b1 a1 98 90 86 83 82 83 83 79 7b 6c 70 64 6b 60 5b 55 5a 57 52 51 45 4b 57 51 51 56 53 56 56 4a 50 51 57 58 57 50 55 57 56 55 58 54 53 54 54 5c 55 5e 59 5a 5b 5f 66 65 62 6d 68 5e 5b 65 5a 52 55 59 5c 5d 56 5a 58 4f 4f 52 4d 4e 4c 56 50 56 56 55 4f 52 4f 56 56 5a 6a 78 73 63 41 25 16 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 06 01 06 16 23 36 53 63 5b 6c 78 7a 7a 7f 6a 5b 4d 54 58 54 54 51 4f 4d 55 4b 50 50 4b 50 4f 53 56 57 58 57 53 64 67 5f 5b 57 50 52 55 50 55 53 59 5a 5b 51 4e 54 56 4f 51 5f 5d 5b 5a 5d 55 52 56 54 51 51 51 4f 54 4f 4f 53 53 50 4e 54 60 5e 66 60 66 64 67 69 6e 71 75 71 71 6a 65 6a 64 64 69 64 66 61 5e 62 5f 60 57 57 56 52 4c 57 51 4d 4b 4e 50 4b 4d 53 52 41 2b 31 31 3a 40 50 5c 6a 6f 8c 9d b3 c9 e0 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f1 d4 b5 a4 9f 97 89 8c 84 85 7d 7e 79 76 6b 6e 63 67 65 5d 51 58 5b 55 56 50 4c 4b 51 4f 54 50 56 4e 5c 56 52 55 52 54 55 4b 55 5a 58 55 53 52 55 55 55 5e 60 53 52 5c 5e 6f 64 6a 61 5e 55 61 5f 64 5c 50 54 4e 55 57 53 5c 54 59 55 53 58 4c 50 57 54 52 51 53 4f 49 4d 52 5b 6b 74 66 4d 2e 20 0d 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 08 14 0f 2d 3c 5b 5c 6c 79 76 7d 7b 7a 58 55 56 4d 49 46 4c 51 51 53 4e 56 47 50 47 50 4b 50 5c 56 58 54 54 5c 5c 53 53 5a 5d 57 57 5e 56
 56 51 50 50 52 4b 52 56 54 58 5d 58 53 5a 50 57 5b 54 4b 53 4c 50 53 54 59 52 52 4a 51 59 59 59 5c 5b 5c 64 62 6b 5f 6a 6d 69 65 6a 65 69 60 65 69 66 64 63 5a 62 5a 5a 53 4f 57 51 56 4a 4e 4e 45 47 54 4c 45 4f 50 4b 2d 2c 2e 38 48 4f 51 64 68 77 8a a5 ba d1 f1 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ec cd b7 9c 94 8b 8e 90 8a 84 85 76 78 79 67 73 66 67 62 5b 5a 59 52 52 54 56 4b 4f 4c 4f 52 4e 56 50 54 52 55 54 52 52 4f 53 59 54 4d 58 57 54 5e 57 57 58 55 54 5a 5f 59 5f 60 5f 57 5a 5d 55 56 54 50 53 5a 4d 54 51 5b 4a 5c 5d 50 54 4f 51 56 51 4e 49 52 52 51 49 40 51 53 69 6b 5d 44 29 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 06 06 18 24 39 4e 5c 62 71 73 79 7e 7a 6d 57 51 51 4a 4f 4c 4d 4f 4a 53 49 4c 4d 52 5a 4f 54 54 56 5c 53 53 5c 56 55 56 55 56 5a 5a 55 57 5a 58 5a 53 58 52 56 5d 51 5c 58 5a 60 5f 4f 54 5a 51 5e 54 4b 4f 4f 50 55 5b 4c 59 52 56 5d 5c 61 69 65 64 59 60 63 64 65 68 67 6a 63 63 68 6a 6d 67 67 69 60 5f 58 50 59 51 47 51 4c 48 47 44 46 3e 4b 52 48 46 4f 3b 2d 2c 38 39 3d 46 55 5e 64 74 89 98 ab ba db f6 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e3 cc ab 9f 96 88 8d 7e 80 7e 7d 7f 75 75 6c 66 64 62 57 56 4a 4b 47 48 56 55 55 59 54 5b 52 57 5c 4d 4e 50 4e 4e 57 53 56 53 5a 56 55 54 58 54 5b 52 52 55 58 54 61 5f 60 64 5b 5f 5d 5b 60 59 51 53 55 4f 57 53 59 59 58 4e 52 50 55 5d 52 56 57 5c 4f 52 4f 4e 4d 4c 4b 51 4d 63 64 4d 3f 30 19 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 09 10 18 19 2d 36 4f 58 6d 71 7a 80 75 69 60 52 4b 4b 4e 51 53 53 56 51 51 44 55 49 54 46 4c 55 5b 54 53 55 50 5a 5f 5c 5a 51 51 53 4f 56 53 58 58 52 56 50 56 4f 5e 58 52 5b 5b 5f 56 5f 59 5b 57 5c 53 59 53 52 4a 50 58 58 59 55 58 5f 59 5a 63 5f 65 69 5f 63 6d 64 6c 66 66 65 6b 6d 63 66 5d 62 64 63 5c 59 5b 5a 5f 4f 4a 4d 43 44 45 3d 3e 43 3d 36 42 37 28 2e 35 42 3f 47 4f 58 5d 72 7e 8f 9b aa c1 dd f3 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f8 dd bb a4 95 90 8b 7d 84 83 82 78 7e 73 73 68 67 62 62 54 54 57 49 48 4e 4c 44 51 50 51 54 55 56 51 5f 5b 52 56 57 52 54 5e 50 55 59 5b 5d 5b 5e 57 4f 4e 57 5d 59 5c 5f 61 56 5a 59 5a 51 50 5d 57 5c 55 5c 55 57 5a 57 52 54 52 54 55 57 55 54 4e 59 5b 53 54 4d 52 47 54 4b 55 58 56 46 2a 20 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 12 24 31 3d 52 59 73 70 74 7e 74 63 57 52 45 48 4d 4f 50 50 4a 51 40 3d 46 46 4d 50 45 52 50 52 4f 50 5c 66 66 65 66 4f 4b 4c 53
 4c 58 4f 53 56 5b 58 61 5e 60 58 66 5f 57 67 63 5f 5c 59 5a 5a 4b 55 51 56 4e 51 52 4f 55 5d 59 5a 5b 5b 64 5a 60 60 5f 6e 5e 62 66 6a 6a 68 6b 6a 60 65 63 5e 62 5e 58 58 4b 4e 4b 42 46 46 40 41 3d 40 3d 3d 36 40 35 27 2c 2c 35 44 3f 3e 51 5b 60 67 7e 8e 9b b6 c4 e2 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ef c7 b7 a2 8e 86 7f 86 82 7e 80 7d 72 70 6d 60 67 5b 5c 55 50 4e 4c 48 4e 44 47 48 4f 49 52 4b 57 59 53 52 50 59 5e 55 59 52 55 49 57 53 52 54 4f 51 5d 50 52 5e 54 5e 5d 5e 5a 5c 55 5e 54 50 59 54 4e 55 4f 4f 54 5a 53 56 4d 54 54 52 58 54 4d 5b 53 57 50 4c 49 4a 47 4d 4b 4d 55 4c 36 2f 0e 13 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 07 09 0f 09 1b 19 2b 2f 42 51 5e 71 70 7e 79 64 50 44 46 50 47 51 4c 4e 44 4a 4c 4a 4b 48 50 55 4f 47 4e 5e 52 51 5a 5c 72 75 6e 62 5b 5a 55 55 50 53 59 50 5c 5c 61 67 65 63 64 62 67 58 67 6a 5c 63 5a 56 5c 4d 56 52 59 55 56 52 59 59 57 55 5b 5a 5f 59 5a 61 64 60 67 6f 66 62 64 61 65 69 61 66 65 61 5b 59 55 58 59 56 4e 44 45 3a 45 45 45 41 31 38 39 39 3a 23 28 33 35 3c 38 3f 4c 53 64 6e 73 77 8b a7 ba cc e4 fc ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff e3 c5 ac 92 86 85 82 83 7f 76 77 71 76 66 69 68 66 57 5e 4f 51 49 45 3c 4a 43 49 4a 50 4f 53 56 4e 54 4e 4b 4d 53 51 58 59 56 52 59 5a 55 5a 51 4d 55 50 51 58 5a 5b 62 60 5a 52 59 4d 50 5b 4e 53 53 4e 5a 53 4e 4d 51 55 50 4f 4b 4e 57 54 59 4d 54 57 51 4f 4d 4a 44 43 43 49 59 52 47 32 19 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 06 0e 12 1a 1d 24 2b 32 42 57 68 6f 7e 7b 63 5d 4a 49 4b 4f 49 50 4d 4f 49 4f 4f 4f 4c 48 48 54 56 4a 53 49 4e 56 5d 67 73 78 61 5b 56 57 58 5f 5f 5f 63 61 69 64 5d 69 65 5f 5c 5f 5b 59 5f 69 64 68 5f 60 63 5c 62 52 54 56 5f 56 5b 5c 57 60 55 64 61 62 5e 66 62 69 65 6a 69 63 69 6c 5f 6d 6b 5c 5c 5e 5b 59 52 52 56 51 46 49 42 41 40 3d 3a 3c 3a 3c 38 32 23 26 30 35 3b 3a 43 53 55 63 63 7b 78 81 99 a9 b5 d1 e2 fa ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ee d8 bf a4 91 8b 89 81 7f 84 7b 76 78 71 6b 6b 65 58 65 5d 50 51 51 4f 44 49 48 48 49 49 4b 4e 51 55 55 5e 56 4f 5d 54 5c 5a 55 50 4b 56 53 54 58 51 51 56 50 57 5e 60 62 60 5f 5c 5d 5b 62 5f 4f 52 48 5a 57 55 58 5a 4d 55 56 54 5a 4d 56 53 4e 50 4f 53 51 4a 55 4b 4c 53 4b 52 56 56 3d 2d 12 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0c 07 0d 13 0b 26 24 2b 3d 44 55 70 79 74 66 4f 4e 47 47 4f 45 46 4f 4c 42 4f 4a 4d 4c 4c 50 4d 4a 4f 4e 4d 51 4c 4f 56 61 6f 5e 57 51 5a
 60 63 5b 5f 67 5f 61 5e 5a 5b 50 5c 5e 57 5a 5c 52 5f 59 64 59 62 5e 5b 5b 52 59 5c 50 52 57 5d 57 57 52 53 5f 61 55 64 5f 66 68 65 67 67 62 56 6a 60 65 68 62 5f 5c 5b 57 54 41 40 40 3d 3e 42 45 38 36 2f 35 39 33 35 24 1f 23 2d 3b 33 3b 44 4a 5c 60 6f 74 7d 89 9d a5 be d0 e2 f2 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff f9 e6 c6 ae 9a 89 7c 7c 6e 7a 79 77 77 72 6a 62 68 5a 60 59 59 56 50 4b 48 48 41 48 47 51 50 4c 4a 50 4b 55 54 4f 51 55 55 53 51 4f 4e 51 4a 54 52 52 50 52 55 55 51 53 5a 66 61 63 56 57 51 53 57 55 53 54 54 4e 4f 58 48 4f 51 55 55 58 4f 54 54 5a 4d 51 4d 4e 49 49 4a 4c 46 52 4c 53 4e 27 22 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 09 0b 14 13 12 15 1d 15 27 2f 3b 4c 5d 70 75 72 5c 4c 4c 43 4f 4c 4a 4b 42 4b 45 4a 4f 4a 52 4f 4f 4d 59 4c 51 53 53 4b 55 51 5b 5b 5e 64 59 56 5f 55 60 5e 5d 57 57 5a 5c 54 52 52 54 58 5b 5a 55 5b 59 5c 54 58 55 5d 55 5b 5a 59 59 56 54 59 5e 59 66 60 5d 5a 64 63 66 68 59 61 63 5f 67 61 5c 5e 66 60 60 57 56 4f 56 51 45 41 42 47 3b 3a 3a 3d 31 30 2b 34 31 1b 1b 24 25 2e 38 40 41 4b 5b 56 67 6b 70 80 8b 9b a4 b9 cd d5 e9 ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff ff fe f1 d0 b3 9e 8c 8a 7c 7a 77 77 74 76 70 72 66 66 62 59 58 61 54 52 51 4d 4d 49 48 53 4e 4b 4b 51 52 50 4f 59 4d 4d 50 56 51 54 50 53 58 54 56 54 52 4f 4e 59 51 55 5b 64 54 55 56 5d 55 53 5a 53 50 53 50 50 56 51 55 50 4d 54 49 51 4f 53 51 51 54 4b 52 49 4a 43 49 4b 4e 4c 4a 55 50 4a 44 29 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 08 05 0e 13 16 13 19 20 32 3f 49 5b 6f 74 73 5f 46 4b 44 4c 44 50 48 51 43 49 45 46 4e 48 49 50 4d 4a 4b 51 54 55 60 58 53 55 4c 58 61 55 5c 5f 5c 56 4f 4d 4e 53 4c 5d 51 55 5c 55 5c 52 55 5b 60 5c 58 59 59 61 5b 5d 67 62 67 65 55 5f 5d 58 5c 61 59 5f 64 62 65 5c 5e 60 65 5c 62 64 66 67 66 5a 61 65 65 54 58 58 4d 4d 49 49 40 43 33 3a 38 2f 2b 38 2e 2b 20 12 18 23 34 33 39 37 4d 4a 61 5b 5e 66 7c 7d 8a 9a 9f b0 c0 d4 f1 f9 ff ff ff ff ff ff ff ff ff ff ff ff ff fb ef db c4 b1 91 83 80 80 7c 78 79 74 6f 72 65 65 5e 66 61 5c 50 55 50 4c 56 46 47 4a 47 45 4b 50 53 48 50 4f 54 4e 4f 56 4d 5a 56 59 53 52 4b 52 53 55 5d 53 52 54 54 58 5e 5a 5b 62 5f 61 52 58 55 53 57 60 54 57 4d 52 4c 53 50 55 52 4f 53 4e 5a 54 50 46 54 51 3f 4b 4b 4a 53 4d 50 55 4f 3d 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0f 0f 11 0b 0f 19 28 29 34 3f 50 6c 75 75 69 52 48 46 4c 41 4c 47 4e 4a 41 43 4c 45 50 4d 51 53 4d 4e 53 5a 5b 5b 50 50 4d 4e 52 53 54
 51 59 53 4f 55 54 53 52 59 4d 53 4f 57 5d 54 54 5f 56 57 54 5b 5c 57 63 65 60 5f 63 6b 65 60 64 64 60 59 5d 4e 5d 63 5d 65 5a 61 60 67 5b 5c 60 65 67 61 68 5f 5d 5d 4e 59 51 46 41 40 4e 40 3c 3b 3e 33 34 29 2e 30 2d 1b 14 18 23 25 2e 34 3e 41 4b 53 59 5e 65 70 7c 84 83 98 a3 a5 b9 d6 de f0 ff ff ff ff ff ff ff ff ff ff ff ec ef e0 bd b9 9e 98 84 7c 79 6d 74 6c 63 67 62 61 5f 5d 5e 51 58 51 57 50 4f 4a 42 45 49 47 4d 4b 4e 4e 4f 52 53 50 4f 4a 4a 53 57 50 55 4d 50 56 53 58 53 56 53 54 60 56 5f 5e 62 58 5e 5c 51 52 54 59 50 55 5c 52 52 4d 51 4c 4f 50 50 50 4f 4c 59 4f 52 4b 4e 4d 4e 41 46 50 4d 4d 4b 57 49 3f 2e 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 07 10 12 16 16 1f 1f 27 37 39 49 5e 72 73 71 55 4d 3e 40 49 4b 49 50 4c 46 4b 4c 4c 4b 4c 4f 4f 53 4c 57 53 54 5e 52 56 55 53 56 53 47 4d 51 4d 45 50 4f 4d 48 4e 52 57 4a 4f 50 4e 58 57 57 55 54 58 54 60 51 5d 5c 62 64 6a 69 69 6c 64 5e 62 55 61 60 62 5c 64 5c 63 64 57 5b 5f 64 62 64 5a 53 5c 58 59 56 52 53 47 46 39 44 41 44 3a 32 2c 29 29 2c 28 28 16 0e 13 14 1a 26 2e 3f 3e 4b 4d 54 5e 5f 64 62 71 79 81 8c 91 a7 b9 d0 e4 ed f6 fc ff f2 ff ff ff fb f8 ed e0 dd c4 b7 9d 96 83 80 76 76 71 6a 6d 72 6a 6c 65 68 5b 5c 53 4f 53 4c 45 47 4d 4c 48 4c 48 46 43 51 4b 54 4e 4d 55 55 51 4e 53 55 50 4c 4d 4d 52 57 54 5b 53 59 53 5a 59 60 55 52 57 58 52 58 54 5a 62 63 63 59 59 53 55 54 56 4f 51 52 4c 52 52 4c 51 48 46 43 47 49 49 45 50 43 46 4c 51 51 34 22 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 08 0f 11 12 0d 17 1b 2c 31 3e 42 56 72 7c 76 5b 4e 49 3f 3b 43 49 49 45 43 42 47 4d 4d 4b 51 4e 4e 48 43 54 56 5c 5d 55 51 53 55 4f 4d 53 52 4e 50 4e 53 4c 58 50 52 4e 50 54 54 4f 50 5b 55 5a 54 54 5b 55 5d 58 5b 5c 57 59 69 60 64 61 57 56 64 60 61 65 54 5e 64 64 64 5f 65 58 62 5f 58 5e 65 5a 59 5f 51 52 49 51 48 3e 41 39 39 34 38 33 37 31 28 2f 2c 19 09 16 08 1c 1d 26 35 3d 3f 47 56 53 5f 6a 67 6d 72 77 84 8c 93 a0 bb cb ce df e4 e8 e0 e5 ef f6 ec ed e2 d6 cb b8 aa 90 8f 81 7a 75 6b 6b 6c 67 6b 62 5e 65 5c 56 5d 52 51 4a 57 44 51 4f 4a 4d 4b 4b 4d 43 4a 4a 54 50 55 56 52 50 56 5a 56 50 57 54 5a 5c 59 55 54 57 54 57 5c 56 5f 56 5a 5a 5d 56 58 5c 5c 5f 5b 63 60 55 5f 57 55 52 53 55 4e 52 52 47 56 46 4d 4c 44 4a 4a 3c 47 4e 4d 4c 4c 4d 37 24 18 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 13 12 19 21 1b 28 2e 37 4c 5a 64 73 79 6a 5b 48 42 48 42 49 50 44 46 4b 46 48 4f 51 4f 4c 44 4e 49 51 5b 5f 5b 5c 54 4e 4c 4b 4f
 4e 52 54 50 51 50 51 53 4e 52 51 58 59 56 55 4c 5b 54 50 5a 52 53 4c 53 52 57 54 5e 55 59 59 5a 5e 5c 55 5c 5b 59 56 59 64 5b 60 68 65 55 63 62 5e 61 60 64 5a 5e 64 57 4b 52 4e 4b 43 43 3b 3d 39 3f 37 29 31 2b 33 2e 1b 0a 0c 0f 15 15 25 31 32 3b 45 47 4d 5c 5b 5f 69 69 68 78 7a 8a 95 a4 b1 bd c3 cc ce d4 dc df e2 df d9 cd ba b2 aa 9d 8d 82 74 71 6f 66 6d 67 68 69 69 65 5d 59 5c 5d 4a 50 59 49 4f 45 43 4c 41 44 4d 44 52 52 53 54 58 58 5c 5e 57 4e 60 5a 53 5a 53 5e 5f 5a 51 5e 5e 59 61 58 57 58 5a 5c 60 5f 55 57 57 62 5c 5d 60 63 5f 5a 62 52 4d 4b 53 55 50 53 48 4b 4b 4a 51 4e 46 49 44 4e 45 44 4d 4c 4b 33 19 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 08 1b 1a 20 22 22 2c 2c 3d 54 64 78 84 76 59 44 44 3b 44 3f 45 3e 4a 41 4a 53 4f 4e 4e 47 45 4a 44 50 52 52 44 47 52 51 4b 49 54 51 53 4c 4a 4d 52 4b 4b 4e 51 54 48 56 50 60 54 4f 4f 5e 4f 55 54 52 58 5b 5b 50 58 4c 53 58 57 54 58 58 5b 5d 5f 60 59 60 5c 63 5d 5a 61 63 5b 5b 64 64 57 5e 5f 61 5a 4f 4c 49 4b 40 42 3d 3a 37 2f 32 30 34 27 2c 28 1b 05 0f 0d 12 12 19 1d 2a 36 3a 42 4d 5b 56 54 5a 69 6d 6c 6f 79 84 8b 95 9e aa b2 b8 bf be d0 ca d3 bd b3 ac a3 9c 90 87 7c 72 70 72 65 6d 6a 5e 69 66 64 5e 5d 58 5a 5c 4f 52 49 4a 46 4b 4d 49 4c 4d 44 4b 4d 4c 53 52 59 57 5a 5d 5d 58 59 54 54 5a 5e 5e 56 53 5c 5c 60 5f 58 58 5b 57 60 63 5e 4e 4e 51 5a 59 54 51 5d 60 5e 59 4f 48 4c 51 49 4b 4b 45 4e 4f 45 45 44 3e 47 3a 43 47 49 51 42 3e 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0b 06 15 19 1e 20 1f 27 29 35 42 4e 56 7f 82 7e 65 4b 40 3e 45 42 41 45 44 46 45 49 49 48 49 4b 4c 45 47 4a 4f 52 4f 54 54 44 4d 4a 4f 5a 50 4d 4b 4e 53 51 4d 55 55 4d 56 46 5e 54 52 56 51 4f 59 50 4b 58 50 53 52 59 55 52 56 54 54 56 5a 5c 5a 54 54 59 5f 61 60 5b 5c 5c 5f 61 56 60 58 60 5c 5d 55 57 50 49 52 4d 46 46 48 43 3b 36 35 32 28 2a 2c 2c 26 1c 0a 09 0b 0c 0f 15 2a 2a 2f 37 39 46 51 4d 54 5b 5f 5e 66 6c 70 77 75 89 89 97 9b 9b aa b3 be c4 b8 b7 a8 9c 9a 8a 84 82 7a 74 70 71 69 6a 64 6a 62 5d 61 65 5e 5d 5e 59 5b 54 58 59 4b 4d 46 47 46 47 48 52 50 52 59 60 61 67 5e 64 68 60 5c 5a 58 57 62 60 54 62 5e 5c 5b 5b 61 56 54 51 57 5c 5f 67 55 51 50 4d 49 52 68 58 58 54 5b 54 4c 50 4d 4f 48 46 45 4c 43 50 40 3d 48 44 4a 4f 53 4f 40 2e 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 05 03 0f 14 1a 18 20 21 30 39 3b 4c 5c 70 85 80 70 4e 46 3d 40 48 46 45 45 39 44 47 54 48 51 50 4e 48 44 51 4e 4d 4d 4e 4e 4e 49 42 4e
 51 43 4a 47 4a 4f 45 48 52 50 55 5a 51 4e 56 4d 54 52 4e 5a 52 51 57 49 56 51 4e 52 4e 5a 5d 56 5b 58 5e 5b 57 5b 5a 5d 5d 5a 57 5b 5d 55 5e 5a 5c 5f 5f 5a 5e 60 53 57 4f 57 52 51 43 49 40 3c 3e 3a 31 25 2b 2c 2b 2d 13 04 06 05 0a 0a 16 1b 1c 28 29 3e 3a 45 41 4d 53 58 54 5d 5c 5f 6b 67 78 78 7f 80 92 91 99 a5 aa b3 9d 9b 81 82 7e 76 74 71 74 6e 69 69 68 64 62 66 68 5e 60 5c 5e 63 5c 56 4f 51 52 4e 52 51 4c 51 58 56 5b 54 5d 5c 63 5e 62 62 59 64 5e 69 5c 5e 62 5d 65 5d 61 61 5c 5b 5a 55 59 59 50 50 55 5f 5a 5c 51 52 48 4a 58 5d 63 5e 58 5b 4c 4c 48 45 48 53 49 45 4c 45 44 41 3a 4b 47 4b 44 50 4a 38 22 0a 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 15 1a 19 19 1f 2a 2e 2f 39 46 58 6a 78 7d 6f 52 44 43 42 44 47 49 48 48 44 44 44 40 4b 48 47 47 3f 3f 51 45 46 4a 45 46 44 49 4a 47 4c 47 44 41 46 46 4b 47 4b 41 55 50 4b 4c 52 4b 53 4d 54 48 50 54 5c 57 53 55 4e 4b 47 54 52 53 5a 52 50 56 51 4f 52 56 52 57 57 54 62 63 5d 5c 59 5c 5d 5b 56 59 51 4f 4f 51 53 4c 4f 41 41 38 37 36 2c 2d 24 34 2a 18 05 06 05 09 01 09 05 14 1c 27 28 2f 3d 48 48 4f 49 53 54 58 5e 59 67 5f 66 7b 7b 7a 83 81 8b 96 93 95 90 85 7a 7d 6c 72 6f 6b 68 62 62 5e 5f 66 5e 61 5c 59 61 59 5f 5d 53 51 5a 4d 56 50 4a 52 4f 53 53 53 5a 5f 63 60 56 58 66 5e 60 5d 66 61 59 67 64 57 5f 57 55 59 5c 56 54 58 57 56 55 54 4b 4b 54 4a 4e 50 50 51 55 4d 5b 55 59 55 4e 52 4c 50 54 49 4d 4a 42 40 3e 44 4e 49 45 43 4a 3f 30 14 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 15 16 21 20 20 27 34 33 3f 3d 46 6a 70 76 70 52 44 42 48 47 44 3a 44 40 41 45 44 47 42 51 45 48 4b 47 45 44 4f 4d 4a 4e 3f 4c 49 4a 49 49 46 46 49 45 47 4e 4a 53 4a 4a 4d 55 4c 48 4f 52 54 4c 50 52 53 4e 4b 4d 49 50 50 55 54 58 57 4d 52 4e 54 59 55 5c 51 55 55 52 5a 5d 5d 54 56 5a 5d 53 62 58 53 59 4f 4c 45 54 4a 4e 41 33 2f 31 34 2a 30 2a 2c 21 06 06 05 03 06 06 0c 09 11 16 1a 29 30 36 41 3c 4a 57 49 54 54 58 60 5d 5c 66 69 6e 62 77 7e 8b 86 85 82 6e 76 74 6d 61 62 65 66 62 5d 61 56 5e 63 5c 5d 52 60 58 57 56 54 4d 50 53 50 4f 48 4c 50 55 50 45 5c 58 5a 60 5b 57 69 60 5c 61 61 57 58 60 59 58 5f 51 53 57 57 56 58 5f 55 52 4f 49 4f 4a 42 51 55 4c 4f 52 59 58 56 56 52 51 4d 51 49 53 45 4b 46 4b 44 45 44 49 4c 47 43 4a 45 3c 28 0c 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 0f 20 19 21 23 30 2a 30 39 49 54 73 76 65 57 4a 3e 3b 42 40 40 41 3c 3f 3e 3b 4c 49 49 48 3b 41 49 46 4f 4a 4c 4a 43 4c 4f 4f
 4f 4a 47 4a 50 49 45 4d 4d 50 4a 48 51 52 51 5d 52 51 4d 53 54 50 4a 4c 52 50 48 4a 4c 51 53 4a 4e 4c 49 59 4b 57 4d 51 55 55 56 56 57 57 5b 56 62 5d 5b 59 5c 5a 51 53 55 4f 55 53 45 54 4c 43 40 37 37 30 2a 2a 2d 31 1a 02 06 05 04 05 06 08 05 10 1a 1b 19 21 2b 32 47 42 42 3d 45 4b 4f 52 51 51 59 55 58 61 65 74 7c 82 7a 78 67 6c 6a 65 68 64 5e 64 64 59 5b 5e 58 5b 55 58 59 5e 4b 60 4b 59 4e 55 4f 4f 51 52 4e 45 4c 51 4c 4e 4f 52 57 5e 5b 5b 5b 59 5e 53 5b 56 54 5b 57 5c 4b 51 60 53 5c 5c 62 5b 4d 45 4a 48 50 4d 46 4b 4e 46 52 5d 4d 56 58 50 53 44 4e 4f 51 46 49 45 4d 4b 44 41 4c 44 46 4a 49 45 34 21 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 13 1f 19 1c 28 23 35 33 37 40 4d 5b 5e 5a 4e 44 3c 3e 43 41 3c 39 42 44 3e 38 3c 44 48 47 46 42 48 4b 44 46 4b 3e 41 40 3e 48 47 4e 45 45 42 41 40 4d 51 42 51 4a 49 53 4f 52 55 4f 56 50 45 56 50 4f 45 49 4f 47 46 46 49 46 50 4e 52 53 4c 55 51 4c 58 52 53 5c 5e 58 5b 5b 5e 58 63 5a 56 5d 60 57 59 4f 53 4b 56 4c 52 4b 42 30 26 33 33 2e 2f 27 14 00 06 05 03 00 06 05 04 0c 0a 12 1f 1f 2b 31 2f 41 3e 3c 39 45 41 44 40 4a 4b 4d 54 4e 53 64 74 70 74 74 62 69 66 65 5d 64 64 66 5b 56 5a 54 5c 5f 5c 63 52 57 52 59 54 51 51 4b 4c 4b 4d 49 42 4c 46 49 4d 4c 4b 55 64 5a 5b 5e 50 50 4e 47 46 4d 56 57 52 4f 4f 4f 53 55 53 5c 52 4f 47 45 4b 47 50 4b 46 47 4d 51 52 48 56 51 49 55 55 4c 51 4c 4e 47 47 49 48 3b 4e 41 48 4a 44 4c 3f 40 2a 15 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 14 16 20 16 1e 29 25 36 3e 43 48 4a 59 50 46 3d 42 3f 46 46 3b 41 38 44 3d 3c 40 4b 45 47 47 48 4b 46 42 44 45 47 42 44 44 48 44 4a 44 3f 41 45 4c 47 41 4d 3e 4a 4a 4c 59 55 53 50 52 4c 45 4a 4e 4a 49 4b 4a 47 43 47 4e 54 58 54 4d 4d 4c 4f 57 53 51 55 55 5a 5c 5a 50 5d 61 55 5e 5c 5d 55 55 58 59 59 56 5a 53 5e 4a 48 36 38 33 2f 2f 32 3a 2f 1e 09 06 05 03 00 06 05 03 0a 06 0e 11 17 27 2a 2e 33 2f 36 34 3d 3d 42 3d 45 41 45 40 4d 4f 59 6a 6a 6a 61 5e 68 68 5e 5c 55 63 5d 56 5c 51 57 54 5c 5e 5e 57 53 53 61 4e 51 4b 55 4a 4a 48 57 4e 4a 51 41 4c 51 55 5e 60 5f 59 57 53 4c 4d 4c 45 4d 47 4c 4a 4f 54 54 55 4d 54 57 4b 4f 45 45 4a 40 4a 43 49 48 54 4b 4c 4f 55 4d 5a 5a 53 54 45 4b 44 47 46 44 46 46 44 42 4d 48 45 3e 3d 33 2b 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 06 14 1c 1b 2e 26 27 33 39 3b 45 47 4e 45 47 43 3e 40 43 3f 37 3e 45 41 3e 45 3e 3b 44 45 47 44 4b 43 44 47 46 41 45 44 47 48
 4b 40 43 3f 4a 42 3b 48 42 48 4e 4d 4a 53 4c 45 50 4f 4e 4e 50 4c 50 44 4e 4e 52 45 47 4b 45 51 48 4b 49 4c 49 50 51 4d 4f 4e 55 55 5a 5a 5d 5b 5c 5d 61 57 62 58 5b 5c 56 59 58 51 4f 57 53 49 38 3a 2e 38 2e 3e 31 2e 23 09 06 05 03 00 06 05 08 09 06 09 0a 10 15 1b 1f 2e 2a 34 34 31 37 3c 3f 3a 42 44 39 46 41 45 64 6f 62 5d 5b 5e 5e 56 5c 5a 60 5e 5b 5b 5c 5c 5e 5c 58 5c 5a 54 55 54 53 56 51 49 51 4f 4c 4f 4f 46 41 4e 4e 59 5b 58 5c 58 51 4e 4e 50 4e 48 42 4a 4c 4b 4d 54 4a 50 5b 59 56 48 46 4c 49 44 48 44 4a 48 4c 5b 49 45 48 51 52 59 4b 59 51 48 52 46 4d 40 47 3b 46 44 42 47 48 4e 45 41 39 31 20 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 07 12 19 21 1a 29 29 33 38 3a 41 41 4a 44 3c 49 40 3b 44 40 3d 3b 39 42 39 3b 3e 49 42 44 42 43 48 45 40 44 3e 43 38 3e 3d 4a 40 40 42 3e 42 43 3c 49 45 47 4e 4c 48 3e 51 4a 48 49 4a 50 4f 44 4a 49 47 4b 44 47 3e 4a 53 4e 51 4e 45 46 5a 51 53 4b 4f 56 5d 5c 57 53 59 5a 5e 5e 5c 5f 5b 57 5a 5a 57 54 55 4b 51 54 52 4b 41 2f 34 2f 2e 2a 34 31 16 0b 06 05 03 00 06 05 03 00 08 06 03 12 17 16 17 25 1f 27 36 2c 2f 30 33 37 36 36 35 3d 3a 4b 58 62 5b 59 58 5d 5e 53 5c 55 56 5e 57 58 5a 54 51 5c 5a 58 49 5d 4b 56 4b 4f 49 46 41 49 4c 46 48 4a 4a 4a 4b 5d 52 50 5d 4a 47 4d 48 49 48 4b 50 44 49 45 4a 4e 4f 4b 4c 54 51 4f 45 46 44 47 48 4c 48 47 4a 3e 4b 45 49 53 52 4d 50 50 55 48 45 4a 47 47 44 42 4c 41 40 49 47 4c 44 3d 33 1e 11 07 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 10 13 1e 1e 1a 24 2d 2e 32 31 39 3a 49 43 3d 46 35 40 3c 3d 3a 38 3a 38 41 47 38 41 40 42 49 3e 44 40 3a 40 45 40 44 45 48 41 47 3e 39 40 3a 3e 43 40 4d 43 45 4a 45 4a 4c 4c 52 4e 50 42 4e 43 46 4c 49 47 45 41 4d 46 4d 4b 42 50 51 4c 4c 53 48 49 4c 50 55 5f 4f 55 55 59 54 59 5a 55 58 57 5e 56 4c 55 51 53 5b 4e 45 3e 36 3d 2e 2a 32 34 2a 1f 01 06 05 03 00 06 05 03 00 06 05 04 0b 06 11 10 1c 1e 25 24 21 28 2d 33 30 38 32 30 35 2e 3d 54 5a 52 54 59 5a 54 54 4f 5e 54 58 53 57 57 57 57 5a 5d 54 53 54 4d 4a 4c 4a 43 48 3e 4f 45 46 46 43 48 4d 53 4b 4c 4f 4d 4e 42 47 44 4b 47 42 51 41 4c 51 43 4c 46 4d 4a 4e 4a 46 47 4c 45 44 47 51 4b 4c 44 43 44 47 4b 4f 52 54 45 49 42 43 46 42 49 40 42 44 45 43 46 41 45 45 43 3f 2b 15 07 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 12 23 20 2a 24 2f 33 34 3a 3d 3f 46 45 40 40 3e 3e 38 3e 3d 3a 3d 44 40 36 41 44 3f 47 48 47 4c 41 42 43 45 3a 40 41 43
 3c 42 41 48 45 43 41 43 45 46 44 48 4c 45 48 49 50 52 4b 4d 49 4d 53 45 53 48 4c 47 41 46 47 4e 4e 43 49 4d 4d 54 4c 4a 52 50 4e 5a 59 50 55 55 5b 58 5c 57 59 55 60 57 56 56 5a 55 56 57 52 3f 47 40 3a 3a 32 34 2f 2f 1f 08 06 05 03 00 06 05 03 01 06 05 03 09 06 05 0b 0f 1b 19 20 1f 2f 27 31 2b 30 28 31 2d 32 37 4f 50 53 54 53 54 53 48 58 52 5d 5d 55 5b 5e 59 5b 5c 52 5b 52 4e 51 49 49 47 45 47 41 43 42 44 44 4b 4b 50 4c 44 4f 42 46 4f 49 47 45 4d 4c 4f 49 4e 4c 43 4a 4e 42 4e 49 48 4e 4b 4e 47 47 50 4c 52 4e 48 46 49 3f 4b 4e 47 54 4e 48 50 4e 4e 4a 41 4d 46 41 4b 42 49 4a 43 49 46 3b 39 29 15 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 11 21 25 2a 25 31 33 40 3f 42 3f 3e 3f 41 3f 40 3e 39 34 37 41 3a 35 3c 3d 44 46 44 41 3e 41 40 42 40 45 3e 44 42 42 40 44 35 41 3e 42 3c 40 40 3e 3c 3e 41 4c 45 4c 49 48 4a 4b 4a 49 49 49 4a 4c 52 48 3d 3b 48 4a 42 46 4a 48 4d 49 55 4d 52 52 50 53 50 56 5b 56 5a 53 55 56 55 5c 56 55 52 5b 5b 56 51 62 55 4c 41 3d 33 35 2f 30 2b 2f 20 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 10 0b 14 12 14 1c 25 24 2f 27 2c 2c 27 2a 28 48 4c 53 58 50 54 56 55 55 54 53 52 53 5e 52 54 5c 5a 54 50 4b 52 46 4d 49 3e 45 40 3d 43 44 3e 41 43 48 4d 4d 4c 43 44 4a 49 44 45 48 48 4d 4e 45 4f 40 43 43 4a 43 4f 42 49 4d 4b 4c 49 4d 4e 4f 4f 4c 49 46 42 49 4e 49 4b 4e 53 4e 4a 49 45 4d 4a 42 42 3e 3e 48 43 47 44 45 3e 3d 36 1d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 11 1f 17 1a 2b 28 30 36 33 44 3d 40 39 37 3c 41 41 3b 41 36 36 44 38 38 44 3f 43 3e 3f 38 35 44 42 39 47 3e 40 3e 44 41 3e 36 3d 3f 40 32 41 3b 51 3d 41 48 51 45 44 41 47 43 4b 4d 44 48 45 4b 4b 52 37 46 42 4b 4e 43 44 45 51 46 48 4a 4e 56 51 4f 56 52 5a 4f 5a 5a 53 54 58 4e 5a 53 56 5b 56 55 56 56 58 5e 50 44 3d 35 34 30 2d 36 2f 1a 08 06 05 03 00 06 05 03 00 06 05 03 03 06 05 05 04 06 08 06 10 15 17 1c 21 22 25 1c 26 22 2d 3d 49 50 4e 40 54 4b 4a 53 55 51 54 4a 50 55 55 58 50 55 56 4d 45 3f 48 40 47 4c 46 47 45 49 41 52 45 4a 4d 49 4a 46 46 46 46 4b 4b 3b 3e 45 3e 4a 3e 4b 48 45 49 4d 4a 43 45 49 5b 52 4d 49 44 4b 48 45 47 3e 41 43 41 4a 4b 4a 52 42 49 47 47 49 3f 49 49 3d 47 40 47 48 46 42 44 41 28 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 12 13 24 2a 2b 2c 34 39 42 36 3b 3a 41 3a 3f 40 3f 3e 3c 39 44 45 40 3c 41 3b 44 44 3d 40 3f 3d 3d 3f 45 37 37 38 42
 3d 41 3e 3e 3e 41 3d 4b 3f 41 4c 49 3f 44 48 4c 49 4b 41 54 4a 50 48 40 4b 49 47 4b 47 48 4b 4e 4c 47 3f 4a 41 4c 50 4a 50 4c 52 51 4f 56 51 57 54 58 59 5c 51 5f 56 54 55 50 5d 52 57 52 60 54 47 3f 41 38 41 36 2f 34 26 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 06 09 04 04 12 0e 13 17 1c 1b 1e 1f 1b 26 44 53 44 47 45 4e 4f 49 4d 4e 51 58 4d 4f 51 54 55 4e 47 50 49 51 42 45 45 43 43 4a 48 45 46 45 49 49 46 48 45 45 45 4d 45 46 4a 4e 46 46 4d 45 44 3b 48 44 3e 40 40 48 4b 4b 58 5b 52 4d 48 41 42 4b 4a 4a 41 44 44 47 41 46 49 47 47 4b 41 46 48 41 3e 45 43 49 3d 43 49 42 42 42 38 1d 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 11 1b 1e 2b 2f 2c 36 3d 30 3b 3e 3b 34 3d 46 41 3a 3e 3c 3a 3c 44 45 3a 42 42 39 38 37 3f 3c 44 3a 3e 3a 37 40 3a 3b 43 3e 3d 3d 35 36 44 3c 44 40 47 44 49 4d 45 4b 46 41 45 43 4c 4a 47 4b 44 42 4e 4c 49 4f 46 4c 4d 49 4b 4d 43 47 4a 53 4f 53 54 48 53 50 4e 5a 54 55 54 47 57 57 5a 4b 55 5b 54 57 58 5d 5b 46 47 3e 38 34 35 3a 37 23 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 06 0e 0c 16 10 17 13 17 19 1c 37 40 40 47 44 4d 4b 46 47 51 47 52 51 52 4f 50 56 50 4d 50 4d 47 41 47 47 4c 49 47 45 49 48 45 44 47 48 49 46 45 44 45 45 49 47 47 44 40 4d 48 47 44 49 40 3f 43 41 40 4b 46 49 49 4b 49 3e 46 47 42 44 40 47 43 45 45 43 4f 4a 4d 3f 3e 47 46 40 46 45 48 39 4b 4e 44 46 44 40 35 21 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 15 23 27 28 3a 36 3d 35 39 3d 37 42 3a 35 3c 3c 3a 44 3a 43 32 34 3d 35 45 3d 3c 35 39 37 37 3c 35 3a 38 40 35 44 36 3f 35 31 37 39 38 3a 41 3b 41 42 3b 4e 43 46 47 4c 3f 48 47 49 49 49 3e 50 41 44 44 49 45 46 4e 4a 52 43 47 4e 4a 4f 49 46 48 4d 51 4e 57 4f 54 51 4c 55 50 4e 52 53 5a 59 53 4f 5b 5e 53 49 40 3b 38 35 40 2b 25 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 07 0e 13 17 16 14 29 42 37 4d 3c 45 41 41 49 47 4c 4f 4f 49 4f 48 49 49 43 52 49 49 47 44 4d 42 47 46 46 48 4a 43 45 41 44 51 49 44 4c 50 41 45 4a 4c 45 45 47 42 43 3f 4a 44 3e 41 3f 45 42 44 4c 4a 44 46 51 45 49 47 44 44 38 41 40 3f 45 43 39 49 39 3e 48 45 44 41 40 47 44 4a 47 3d 4c 35 35 32 1a 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 16 23 27 27 34 40 3e 3c 3b 3f 36 3c 40 36 40 3b 3c 44 3f 46 33 3c 39 38 3f 3f 37 32 40 37 35 39 34 45 3e 44
 33 39 39 3c 3f 3c 34 3e 43 3c 45 3e 3f 45 47 45 47 42 45 4a 4b 48 43 52 4f 48 49 43 49 4a 4d 42 4b 4c 45 4e 42 48 4b 4f 51 48 4a 44 4f 4e 4a 51 57 52 55 53 50 59 58 4f 52 5a 56 54 52 5e 64 62 51 49 44 40 40 3d 3c 3a 2b 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 00 06 0f 08 11 07 18 2d 41 3f 40 3f 46 4c 49 49 49 50 4f 52 4f 49 52 45 49 49 48 44 47 45 4f 45 45 42 42 4d 4c 43 49 46 40 48 4c 47 41 48 4a 54 4f 4a 46 46 42 4c 50 46 44 3b 44 42 40 3e 47 43 42 47 3e 3e 4a 4a 3d 42 4b 3a 47 45 4a 45 46 46 4b 3f 48 43 43 4a 43 45 46 44 48 43 45 4e 44 49 3f 38 25 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 0c 21 34 33 32 32 3f 3a 42 40 38 3c 39 3a 3f 41 3e 31 33 39 3b 38 3a 30 39 36 3e 35 43 3a 40 3e 3e 3f 36 3c 3d 38 3b 40 38 33 3c 38 38 38 40 40 38 41 43 43 44 52 46 48 4d 4d 4a 49 4a 49 48 45 43 4c 4a 52 4a 43 43 48 4a 52 4b 4d 4a 4f 4d 4c 4f 4d 4d 54 4c 53 5a 52 52 54 55 52 54 59 60 55 5b 61 5b 5a 49 42 3f 3f 38 38 3d 25 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 06 05 03 0f 09 09 1d 38 3b 42 42 43 4d 40 46 49 41 55 4c 48 45 50 4a 49 45 46 48 48 41 46 45 4b 45 43 4e 4f 48 4b 44 48 47 51 49 4b 42 50 4c 42 45 49 46 3a 41 44 3f 3d 4b 48 44 3e 3f 45 3e 3f 4a 42 39 3c 49 45 47 3f 43 49 38 45 40 43 44 4d 47 4c 3f 45 3b 3c 4a 3a 3d 41 42 45 41 41 45 36 2f 1a 08 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 0f 18 26 31 34 40 3d 2f 38 38 3e 36 33 38 40 3f 35 3f 3b 3b 32 3f 3a 33 34 3b 41 38 36 41 44 37 39 37 34 37 37 37 3a 33 35 3e 36 41 3e 39 39 3f 3e 3b 42 44 45 47 46 42 54 55 4e 55 50 46 45 48 4b 4d 54 50 40 45 4b 4c 42 46 47 45 4e 4e 49 4c 4d 42 51 54 50 4f 4f 54 55 52 58 50 56 51 54 56 5a 5c 60 51 50 4b 44 43 42 3c 3c 24 0e 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 0a 21 34 3a 37 3f 41 42 44 45 44 4d 42 4c 4d 49 46 48 45 47 41 4b 42 47 4f 4b 4f 47 4b 4d 41 4d 47 3d 44 45 44 41 49 44 45 46 45 44 44 44 49 44 39 45 46 47 3d 43 4a 3a 4c 48 46 45 4b 45 43 45 40 48 41 44 43 3d 44 46 47 42 41 41 44 48 3e 47 3f 40 41 42 46 41 41 43 42 49 3a 22 12 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 13 1a 22 32 3a 38 35 41 39 3b 3c 30 33 3a 35 3b 37 38 3b 33 34 2b 33 33 36 3c 3f 3a 3b 3e 42 39 3d 3e
 35 3a 3f 2f 38 33 3a 3c 3d 36 3f 40 41 3d 39 3e 3d 41 42 46 42 4c 55 4f 52 4a 47 44 47 46 53 3c 27 34 51 4d 48 44 41 47 49 4e 49 45 40 45 45 4b 54 4e 55 4e 4b 4e 52 4d 5a 52 53 54 5a 62 58 58 5c 50 4e 48 41 49 37 42 2f 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 1d 2f 3f 43 3f 3b 45 41 3f 44 3f 48 41 49 4d 4b 3c 4b 4e 44 45 4b 48 48 41 4a 50 47 49 4c 42 42 48 42 4d 45 40 3a 3d 48 4b 41 3e 4c 41 42 48 46 47 48 44 44 42 40 42 4c 3e 44 45 46 49 41 42 40 3d 3d 49 44 46 45 47 4d 43 3a 44 44 44 45 46 41 43 40 42 49 49 44 49 44 3d 2d 1a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 13 27 2a 35 40 33 39 3a 39 3b 3d 36 3b 33 35 3a 38 39 39 32 39 36 3a 3a 39 39 3b 37 39 3e 39 3d 37 35 37 38 3b 3a 3b 3a 3e 39 3c 42 3a 44 3c 34 3e 3f 36 40 3f 47 4b 4c 4b 5b 4c 44 4d 43 4c 47 45 4a 4d 4f 46 43 49 48 47 4d 45 45 49 45 48 4a 44 47 47 48 52 58 59 55 5d 54 5a 59 59 50 5c 60 5e 56 51 52 4f 44 44 43 3a 37 14 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 12 33 36 3d 38 3f 44 34 43 42 3f 46 43 4e 4b 43 45 40 41 3f 42 49 4d 46 4a 4e 4c 45 49 4e 52 48 3e 46 4c 47 47 46 4d 4f 48 47 46 40 3b 49 49 44 3f 43 3b 4d 3e 3e 47 50 3e 45 47 45 4a 43 47 45 3d 41 3d 4f 3d 49 37 48 40 44 4d 47 48 49 4c 3d 41 41 48 41 3e 4e 42 3c 38 26 17 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 06 05 16 2b 2f 35 33 3c 39 3a 41 40 36 3d 38 2f 36 36 39 37 3b 39 38 32 3b 34 3b 2d 3a 3b 37 3d 35 39 36 32 36 33 37 41 34 3a 3b 37 36 34 3f 44 38 3c 40 3f 3f 3a 40 46 43 4d 53 54 47 4c 46 42 52 49 45 40 43 4b 3d 44 47 3f 4c 4c 49 49 41 4c 47 4c 52 4d 4b 49 51 51 4d 56 4f 52 55 52 5a 62 54 5d 59 51 55 48 40 49 3d 3c 30 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 16 29 38 46 39 40 39 3f 3b 42 3f 49 3e 48 42 43 44 45 48 45 44 4f 40 4a 4a 4a 4b 4b 41 48 44 48 46 44 4d 42 46 42 42 41 48 4c 3f 45 38 43 47 48 43 44 43 45 3f 3e 3f 48 3d 45 3f 42 3e 49 3b 46 39 42 45 40 42 46 42 44 41 46 47 47 3e 43 43 43 43 3a 45 45 3f 48 3d 3d 2f 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 12 30 28 30 30 3c 36 3b 3e 39 3c 36 34 2f 37 31 38 32 36 30 2b 35 38 3e 38 3c 37 35 38 30 3e 3b
 33 35 42 34 3c 35 39 36 37 3b 37 38 33 41 3f 41 39 3a 3c 47 36 3e 38 40 4a 51 48 41 49 42 47 49 4a 43 45 4b 42 41 41 44 40 47 50 4e 47 45 3e 45 4b 50 4d 50 4c 53 4b 54 56 51 56 5f 5c 5d 61 55 52 4e 46 50 4e 42 55 40 38 24 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 31 39 3d 35 40 3e 43 3e 41 3a 3e 45 47 46 43 46 4b 49 45 45 48 43 45 48 47 41 4a 48 4c 49 47 46 4a 48 44 3f 43 45 43 3b 47 47 47 3f 44 3f 3e 45 4b 40 43 4b 46 4d 42 45 47 46 45 3f 3a 43 46 41 41 48 47 3c 49 44 44 45 4a 49 4a 48 40 42 3f 48 44 47 46 45 44 3a 36 21 10 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 28 35 3a 3e 3c 38 3f 39 3b 33 38 3b 31 2e 36 33 32 31 2e 3a 35 3c 31 3a 37 37 3c 35 3b 3d 3a 35 3d 36 37 35 38 42 3a 37 3b 41 3b 3b 39 41 3d 43 39 3f 3f 3d 41 44 45 3d 4d 52 49 49 4b 4b 50 4d 55 4c 43 4c 47 51 54 46 4a 49 45 44 51 44 41 41 4f 51 55 55 55 53 57 53 56 5e 52 58 5e 57 54 59 4b 52 50 4c 4b 4b 39 21 08 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 13 2e 30 3f 3c 44 37 47 3e 3f 41 54 42 40 46 49 40 48 46 49 4c 50 4f 53 46 4b 4f 47 4a 47 44 46 49 4a 46 44 45 3d 47 42 41 4c 42 3f 40 47 3c 44 49 45 51 45 40 48 45 45 3b 41 43 45 41 46 47 42 49 4a 4c 49 41 4a 40 4b 45 49 43 43 45 4a 48 4b 4c 46 44 44 43 47 3a 2b 18 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0f 25 39 38 3a 3b 3b 35 2b 37 2b 33 3b 34 3a 33 3a 2f 39 31 37 33 38 35 3b 3c 39 3b 34 41 3d 32 35 39 36 3a 3b 3c 33 3b 3f 39 3a 3a 38 39 40 38 45 41 3e 42 41 3f 40 48 4d 57 45 3c 47 4a 57 57 52 4d 48 47 48 49 54 45 40 43 45 4d 49 4b 45 4c 50 4a 48 49 4b 47 4f 54 5c 64 5d 5e 52 59 56 56 49 55 53 4f 55 4a 3c 21 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 29 30 3d 3e 46 3b 3b 3d 3c 3e 43 44 44 43 52 47 48 49 4c 47 4f 4b 4c 42 4b 3e 49 50 4b 4f 4a 40 4d 45 40 47 46 48 48 48 46 40 47 47 43 4b 47 3e 44 45 4d 3f 40 3e 47 42 41 42 42 3f 44 40 44 42 44 44 50 45 47 49 42 4e 4a 43 4d 40 47 45 49 4e 49 43 4e 44 3f 2e 17 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 1f 2b 33 3a 3e 3a 34 39 40 33 3a 2e 31 35 32 34 36 35 2b 39 32 41 31 36 3a 38 34 33 32
 34 36 3a 2e 3a 35 36 36 3a 36 39 3c 34 3a 38 3b 4a 3c 37 44 3d 3e 46 40 4d 3e 3f 44 47 46 45 47 59 50 54 55 54 48 4c 54 4f 42 4c 40 40 4a 3f 4b 46 43 4c 51 54 4f 51 52 58 52 52 59 5b 5a 51 58 56 5c 57 50 4a 43 47 45 3f 23 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 28 37 44 38 47 47 44 3c 41 44 46 52 4d 53 4e 4a 51 42 46 44 45 46 48 48 46 48 41 4d 46 3f 44 45 4c 4f 4a 3a 42 50 42 45 44 3a 47 43 3a 49 3c 47 44 45 49 3e 4a 45 47 46 45 4b 42 3f 41 3e 41 45 4c 3d 46 45 44 44 42 42 46 53 4c 49 40 49 44 49 49 4d 44 3d 35 26 19 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 08 0b 1e 37 2c 37 3b 3f 32 35 37 40 30 36 33 3e 2d 2f 37 2e 37 37 3f 3c 3d 3b 39 39 36 33 3a 3d 37 3e 3a 39 39 39 34 37 3c 36 37 40 39 3d 3a 39 41 45 3f 49 4d 43 44 40 44 45 4c 43 46 45 4b 4b 4c 4f 50 50 53 5c 5a 4b 4b 4c 45 46 47 50 48 4f 49 4f 4b 5a 52 51 4e 59 58 5b 5b 5b 57 5a 53 4f 53 54 57 4d 4b 48 37 26 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 10 2f 39 41 3c 3a 3c 3e 45 49 4e 4c 52 58 4e 4e 42 4f 4a 52 40 3f 4b 47 44 4c 4a 4f 4a 44 4c 4a 48 4d 47 4e 43 4e 41 49 4b 46 48 43 4c 44 41 44 4b 43 49 42 40 49 3b 49 45 42 51 44 38 3f 40 4f 4d 4c 45 44 3e 48 45 45 4b 46 49 4a 46 46 50 4b 46 44 45 48 3f 2e 1e 0d 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0a 15 2d 32 34 3d 36 34 3c 39 38 35 2e 3b 38 36 36 31 3a 38 3c 3c 35 3e 3b 38 39 40 32 33 43 3a 3c 3d 3b 38 3b 3e 3a 3a 41 42 3f 39 42 3b 36 3a 3a 36 42 41 47 41 41 49 45 43 46 41 48 4f 50 52 55 59 4f 50 59 5e 53 55 46 49 43 47 47 45 4d 4f 4e 4c 53 4b 54 53 53 54 57 59 56 59 59 57 55 55 4e 4d 4e 55 4e 42 2d 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 27 3b 48 42 3f 42 41 4a 43 50 54 4e 52 4c 4c 41 4b 48 4c 48 3c 4a 47 45 44 45 4d 41 51 49 51 4a 4e 4c 48 4a 47 3c 44 45 48 45 47 3e 3b 4a 47 48 4a 45 3f 44 46 44 42 44 3b 39 45 42 50 3f 48 46 45 40 4b 41 3d 3e 44 54 47 4e 55 49 41 45 3f 40 3e 3d 3e 36 26 16 11 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 1c 32 2f 39 3b 30 38 35 38 38 39 2f 3c 30 35 33 3b 39 35 3d 38 3f 3f 3e 3b 34 39
 43 3b 37 3a 37 3f 39 3b 36 34 3d 42 34 36 3c 45 3a 40 3d 45 38 42 40 40 44 40 41 46 45 42 41 47 47 4e 4d 51 4b 4d 50 54 56 55 51 48 42 44 45 4b 4b 45 4c 4d 4b 4f 58 51 53 53 59 5d 58 5e 4c 55 4e 56 58 50 49 51 45 49 46 24 0d 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 29 3e 43 42 3f 3f 42 42 52 4a 57 3e 47 46 45 46 41 42 42 41 4a 44 42 47 4a 45 42 40 43 4d 45 46 45 47 42 49 40 41 46 41 3f 41 41 44 3f 44 45 43 3f 3b 3c 3a 46 42 44 4c 45 47 48 3d 3e 3b 41 44 48 44 45 46 43 40 4c 4e 47 4e 46 47 4a 44 45 46 47 44 3b 2f 1f 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 12 23 2f 37 38 36 35 3c 3a 39 3c 38 38 32 35 39 3a 38 3b 37 34 3d 3c 3b 3b 3c 44 38 35 39 35 33 3a 38 38 3a 40 3e 35 32 3f 42 40 40 36 3e 47 3f 3b 46 3d 3f 44 43 48 44 46 43 50 4c 4d 48 48 50 4f 4d 53 54 52 50 47 43 4e 3e 4d 4a 46 46 50 52 53 56 4e 4b 55 50 5b 57 58 5b 57 58 5a 53 55 4f 51 4f 46 3e 2f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 40 4b 40 3e 42 42 49 4d 49 44 3f 45 3e 45 45 46 4c 3f 44 4b 49 4d 48 58 40 45 47 49 4d 4e 46 44 47 3e 42 47 48 49 47 4a 3c 46 41 46 4c 47 44 4a 47 4c 44 43 42 4a 48 3e 43 43 3e 46 40 45 4a 4a 44 4e 43 42 4a 42 40 50 4d 51 46 4d 4f 46 4a 4b 37 3b 1e 17 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 11 1d 35 32 32 38 2e 39 34 3b 33 2f 3a 3b 33 33 3a 3e 35 3e 3d 3b 3f 36 37 41 42 45 34 37 3c 3e 38 38 3b 40 37 41 3f 40 41 42 43 3f 3e 44 39 42 43 3e 43 40 40 47 45 4d 4d 4b 49 4b 4e 46 4b 4b 4b 52 53 4f 50 4f 49 4f 41 4c 4b 49 48 4d 43 55 4e 54 4d 57 56 56 5d 55 51 49 50 4f 53 51 50 50 4a 4e 46 35 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 26 3d 47 44 42 4a 4c 44 45 3c 43 3f 44 48 44 43 42 48 4e 44 46 4d 48 46 50 48 4a 45 4f 46 4e 3f 4b 49 3f 43 40 3e 47 42 49 4b 43 45 43 49 47 3d 43 44 44 45 44 41 3e 48 44 44 42 3c 4d 47 40 49 46 3b 46 44 47 45 4d 4a 49 50 4f 48 4d 44 44 4c 41 3d 2a 11 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0a 21 26 2e 39 3b 37 34 39 38 38 37 33 38 2c 31 33 3b 37 36 3a 41 40 3b 3c 37
 32 3d 34 37 36 38 39 3e 3d 46 3b 3b 3e 3e 3d 3d 3a 39 46 45 3e 42 43 3c 3b 3e 38 41 3d 46 41 45 46 45 46 49 48 50 4c 54 4f 4f 4d 4a 45 49 47 4a 49 43 4b 46 4d 4c 4a 4d 50 53 59 51 54 58 59 4d 54 4b 5a 47 4a 4e 4d 43 3d 33 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 08 20 35 49 41 4b 47 4b 45 41 43 43 48 46 41 49 4a 46 45 44 41 47 47 45 4c 4b 3f 4e 49 46 42 48 48 46 44 45 40 40 47 3f 43 42 47 46 44 40 3c 51 40 3e 45 47 3e 41 42 48 4b 46 40 3a 3e 3b 45 44 42 43 3f 43 3a 43 47 47 47 43 49 54 4c 4c 46 41 3d 3e 26 1f 0c 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 20 2a 34 2f 37 32 3b 30 34 39 39 36 3e 33 35 3b 39 39 41 42 36 36 39 30 3a 3b 34 34 34 38 3d 35 40 37 3a 39 38 3d 3d 39 3d 3c 44 42 43 3f 41 3d 3f 3d 45 44 42 45 4a 40 4a 4c 4b 4e 40 4a 4d 4f 51 4f 54 4d 43 49 52 4b 55 49 4e 4f 50 4d 4b 44 4c 5b 57 58 5a 53 52 54 4d 4a 55 4e 51 55 4f 4a 3d 36 15 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 2a 4d 51 4a 49 53 46 47 48 47 44 46 40 41 4a 44 43 45 45 44 47 40 45 42 43 4b 3f 49 44 4f 4c 3d 44 3e 4a 3c 3c 45 3f 45 41 4a 4a 4c 49 43 44 44 42 3f 42 41 4e 45 49 42 3b 45 3e 3e 46 42 40 49 4d 44 46 40 44 4a 47 47 4f 49 55 4a 4a 43 44 3b 3c 1d 1d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 16 24 2b 2c 35 37 36 45 3a 3e 3b 33 31 38 35 40 37 35 44 39 40 41 36 39 37 3f 33 41 38 38 39 3b 3f 48 36 3c 39 3d 41 44 42 3f 42 3b 3b 45 3d 3f 43 41 49 41 40 3c 40 4d 44 47 51 45 4d 47 46 45 4c 56 4a 52 44 46 4d 48 4d 52 4a 4d 4e 56 4e 4d 4c 47 55 4d 4f 55 4e 56 52 51 51 4d 4c 50 48 4b 3b 35 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 31 59 56 49 49 3e 44 45 47 42 3e 37 48 3e 47 45 4d 49 4c 44 49 43 48 42 4b 45 44 49 48 46 43 47 49 3e 44 44 45 4e 43 3f 47 43 43 41 3e 42 44 44 3e 3d 44 3a 41 45 42 3e 3c 43 41 44 4d 45 42 41 52 4b 47 45 45 43 45 47 49 47 4b 4e 4a 43 43 3e 30 16 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 20 29 38 3b 44 3b 34 35 33 3a 32 38 30 33 3a 35 39 34 3a 34 31 38 38
 3f 38 3f 39 3d 3d 36 3a 37 33 3e 42 3b 3b 3a 3d 4a 39 45 40 41 39 3d 44 3f 44 45 3f 3d 3d 3e 3f 45 3e 45 46 44 45 47 48 4b 53 52 49 47 42 44 47 45 43 4b 48 4b 53 47 46 47 4b 43 58 52 50 47 4d 50 52 51 4e 53 4d 45 4b 49 3a 10 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 26 56 57 50 49 3f 44 43 41 38 44 44 3a 45 42 48 49 3f 43 3d 49 4a 43 4a 4a 45 40 42 46 43 49 3b 39 44 43 42 3e 46 46 47 39 44 43 3c 42 43 3e 40 48 3c 40 3f 41 37 45 3b 46 43 3f 48 47 42 44 38 42 47 42 43 4b 4c 4f 4b 4d 40 4e 4c 3d 48 3d 30 1e 12 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 09 10 22 2d 34 36 3b 34 3b 43 3a 39 31 38 3a 3b 35 39 40 3a 41 3e 38 35 3c 36 3f 3b 37 3a 3c 37 36 42 3d 35 3f 41 3e 3f 41 43 45 3f 3a 47 41 44 46 3d 45 49 3b 41 4a 41 48 42 46 47 47 45 51 50 47 49 4c 44 4d 4c 46 50 48 4e 4e 47 4e 52 49 4d 4f 50 4e 54 50 51 55 4c 53 50 4d 48 47 4f 56 4a 44 32 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 21 44 45 3f 48 41 3e 40 3d 40 44 48 4c 40 49 48 43 46 44 45 4d 44 4a 49 4d 46 45 46 4e 48 42 3a 46 41 3c 45 40 4d 48 47 49 3b 3f 43 3c 41 46 41 41 41 3c 41 48 41 48 3f 39 4a 4a 47 40 3e 41 51 46 43 43 48 49 4c 50 49 4f 4d 4d 44 3d 3b 3c 26 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 0a 15 2c 32 36 38 34 37 3b 32 33 32 36 36 35 3c 3d 36 38 38 3a 3a 39 3c 3e 37 3f 37 3f 36 3d 35 3f 40 3a 3f 43 3b 49 3d 3b 40 4b 36 39 4a 42 45 4f 3d 4b 44 40 3c 42 4c 41 4d 48 41 46 44 49 4e 49 4b 48 43 47 44 51 48 4b 50 43 4e 50 4a 47 4d 4d 4f 58 4c 5b 54 4c 4c 4d 4c 45 48 44 52 49 4a 32 11 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 20 3c 44 40 41 48 41 43 3f 40 41 40 45 46 49 46 42 40 48 40 4c 46 4a 49 49 49 44 4f 4e 49 4a 42 40 48 44 3e 39 43 40 3d 40 3e 3b 49 45 43 44 3e 3a 42 44 32 4a 41 44 46 3c 3f 46 41 41 42 45 49 45 48 44 49 45 4a 49 4b 50 53 4b 46 42 3c 27 1c 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 22 24 2d 31 3b 43 31 40 39 3c 36 31 3a 34 36 32 30 31 38 3d 38
 40 35 35 35 3f 40 3a 34 3b 3b 3e 3e 3d 41 44 43 41 3f 3f 41 36 49 41 41 3f 43 48 44 41 40 48 43 3a 44 43 43 4b 45 43 4a 46 4b 48 4e 46 43 4b 4c 4c 44 48 4b 45 4a 4a 4b 4b 48 4c 4e 4d 52 4b 4a 4b 48 4a 4c 50 4a 51 46 41 39 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 17 37 44 3f 3e 4b 3b 3d 47 3c 42 47 44 4b 45 43 47 48 49 39 42 4a 4f 40 4e 46 43 47 43 42 43 3d 3d 40 44 44 3e 41 46 3f 4a 45 43 3c 45 49 45 48 3d 3f 43 3e 3e 46 44 44 3e 45 3d 3d 47 47 42 44 44 4d 45 41 45 49 43 4d 4f 49 50 43 31 2b 24 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0e 15 24 26 2f 39 3b 42 3a 3d 34 36 36 38 38 3a 3a 3c 3b 36 33 39 3e 3f 3b 30 34 39 39 3b 3a 3a 3e 36 3e 3b 44 44 3f 40 37 46 3b 49 3f 3a 3a 3c 39 40 3d 41 3a 44 41 3d 44 41 47 47 48 48 47 3c 4e 41 4b 4f 4c 49 4a 4a 43 47 48 40 47 46 4f 4d 4e 4e 4a 4b 4c 48 49 45 54 53 4d 4a 4c 46 47 33 15 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 1d 35 44 35 3b 3c 40 42 3f 3f 4a 41 42 3e 44 46 48 3e 48 48 4d 45 4b 45 48 46 4a 48 4a 44 49 3e 3d 49 45 44 3c 44 40 3d 3f 40 44 3d 3b 42 3f 47 3e 3e 45 3e 3a 3e 41 41 3d 47 3f 3f 45 45 44 4f 4b 47 45 47 47 4c 42 45 4b 44 49 3b 38 23 1c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 19 27 35 3a 39 39 3c 3b 39 37 3a 37 39 3b 3f 39 37 39 41 3c 3a 38 42 3e 38 36 38 3a 3b 3c 3b 3e 43 3a 3e 44 47 3e 40 3e 43 40 41 3e 3c 43 39 44 3d 3b 41 43 46 3e 40 47 46 40 42 45 4a 4c 46 44 4e 44 3e 49 49 4c 44 47 4b 48 42 45 4d 4b 4e 4e 47 4e 48 43 49 4d 48 45 45 4b 45 48 48 3b 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 19 2c 43 38 3c 36 38 3f 46 3d 45 3e 3c 47 48 50 44 4e 4d 44 46 43 4f 4e 4e 49 44 44 45 46 47 3f 3e 4a 44 3a 42 3c 44 45 42 46 40 3b 44 3d 49 42 44 3b 40 3d 40 47 45 48 4c 3f 43 41 4a 49 49 40 47 44 46 46 4f 45 4b 49 49 43 41 37 29 16 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0b 20 2d 35 3e 32 39 3f 38 3c 37 35 39 44 3f 37 42 39 38 3f
 42 39 3e 40 36 3b 3e 39 40 41 40 3e 40 3b 3c 44 48 42 3d 44 42 44 3b 37 48 40 41 3e 38 44 3e 3e 41 43 3d 43 3e 44 3f 44 4c 3d 3d 40 3d 40 41 49 3f 4b 47 44 4f 41 4b 52 4a 4d 49 48 51 4e 4a 48 48 4e 4c 4c 4c 43 4e 48 41 3b 19 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 2d 3c 41 3f 45 43 3c 46 40 46 3c 42 44 46 4c 46 50 47 4a 4f 48 49 48 4f 4b 44 4a 42 43 43 3c 3a 38 3d 44 46 3c 44 3f 3d 41 3d 43 43 41 45 3d 45 3d 3d 3c 44 3a 45 40 3b 41 3c 42 43 48 44 43 41 3e 3d 40 3d 4b 43 45 47 41 3a 2c 12 0f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 0c 21 31 30 39 3e 3a 37 36 36 3c 41 3c 35 43 31 31 40 32 3e 3b 37 38 3e 34 3c 3d 39 3e 3b 45 36 43 43 45 3d 44 47 3f 40 42 45 3f 40 3d 35 3d 37 3d 3f 40 40 3c 41 42 3f 40 40 41 43 3c 49 44 41 4c 42 45 3d 41 3d 43 47 49 48 46 4c 46 4d 4d 46 45 4a 45 4d 42 49 42 46 46 44 44 38 3d 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0d 28 34 3c 3d 41 42 3d 3e 46 40 46 47 50 48 46 49 44 4a 50 50 46 45 48 49 44 42 44 4c 42 3c 3f 3c 46 40 3f 38 41 45 40 41 4a 46 43 39 3e 3c 3a 46 45 44 44 42 40 4b 3b 41 3d 40 40 47 43 41 45 49 42 45 39 4a 3e 3f 3a 48 3d 30 1e 12 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 09 15 22 34 33 3d 3b 3b 38 3f 3a 39 3f 3b 41 3e 3e 37 3c 3b 40 3f 3e 3d 3e 3e 3c 3c 40 42 44 39 49 40 47 44 3c 4a 44 3b 43 41 3d 45 3b 3d 47 34 3e 42 3d 44 45 42 3a 3c 36 46 41 40 42 43 3f 38 49 48 42 49 46 41 48 3a 47 4a 40 44 4d 52 47 47 4f 4c 49 4c 4f 4d 4d 4a 42 47 48 40 40 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0f 32 3d 35 41 41 3e 44 3d 50 4d 49 48 3f 41 4c 45 4d 4f 46 49 41 43 48 4c 4d 44 43 43 42 42 40 3d 3c 39 3b 3e 49 45 49 3f 3c 41 40 41 45 41 3f 43 45 3a 43 3e 40 40 3e 3e 40 45 40 47 45 42 43 4c 4a 4a 44 4d 4a 42 41 37 2a 20 0d 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 13 2a 34 3c 39 37 36 3a 35 47 37 36 3c 36 30 35 42
 39 41 32 36 38 3d 33 3f 3f 3a 40 3d 42 46 45 3b 3e 44 3c 3e 44 41 42 3e 3d 3a 36 3e 3e 3e 40 42 37 42 41 41 38 3e 42 3c 40 38 42 3b 3e 44 3f 3e 44 41 3f 45 43 46 45 40 48 42 4b 44 41 4a 49 48 4a 46 42 4a 46 42 49 45 41 37 1f 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 29 44 3f 45 3e 40 48 44 48 3e 49 46 42 49 4a 50 48 45 45 4a 45 4a 51 3b 44 43 4b 42 3e 44 37 41 3e 36 3b 46 40 45 40 3d 40 49 3f 3e 3e 44 40 44 3c 44 3d 39 3f 3f 46 3f 44 39 41 47 42 3e 4a 42 45 46 52 4f 47 50 36 2f 1d 12 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 11 1d 2f 34 39 34 3b 33 3a 44 3a 36 39 36 41 3a 32 3e 3d 3e 3d 38 43 37 3b 3f 3b 3b 3c 3f 43 3d 39 3a 3a 3a 44 42 40 43 32 3d 3c 3c 3a 3b 3b 3a 41 3e 3c 43 40 3a 3e 44 3d 40 44 4a 44 3e 3e 43 43 3b 3f 40 46 45 4a 47 40 47 43 47 49 4b 41 46 46 47 45 46 3d 46 3d 42 46 48 3c 20 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0e 2c 42 44 4a 48 43 3b 45 4e 46 4c 47 44 4d 46 55 47 4c 45 44 4c 49 47 4a 39 3e 40 3c 36 43 43 41 3b 3d 42 41 40 3b 3e 41 3c 44 40 3b 3f 3c 41 3e 42 45 3b 3b 37 42 41 44 44 42 3d 3a 47 42 45 4f 45 4c 4f 52 57 3b 37 29 0e 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 2a 34 35 2d 36 3c 35 3b 42 3b 42 39 38 3d 3a 45 41 3d 3b 3a 41 40 40 3b 3e 3a 3e 3d 46 41 3a 41 3b 44 41 3b 40 3e 3c 40 48 35 3f 41 38 3f 3d 39 38 39 42 3a 37 3c 3f 41 3f 39 39 49 3f 44 47 4a 42 41 41 45 48 47 3f 44 3e 51 49 4b 44 41 46 40 46 45 44 3c 44 47 40 3e 3b 1e 07 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 29 3f 3f 44 43 3a 40 46 42 4b 48 4d 56 4b 50 50 46 4b 46 44 4d 44 4a 46 3e 43 49 46 4a 48 46 3b 44 44 41 3b 3e 3c 41 43 3c 41 41 3d 46 3f 42 3e 43 3e 40 38 3b 43 45 3e 43 41 41 46 45 47 52 52 51 47 4d 4e 3a 34 24 11 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 0e 19 24 35 34 38 3e 40 3f 3d 3f 39 3e 41 37 45
 3e 47 36 38 36 45 3d 45 3d 45 34 3c 37 41 43 39 40 41 3f 49 43 39 3d 3f 40 38 3d 3d 37 40 3e 46 49 3d 42 43 39 4a 40 41 43 42 3a 45 4a 42 39 3d 42 40 43 44 41 45 44 39 4a 3d 41 44 47 4f 48 44 3c 46 45 44 45 42 3f 3d 43 3d 1e 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 29 45 3e 49 45 48 4a 45 4d 50 4a 4e 4d 4e 51 52 4c 54 44 4d 42 41 3c 48 3a 3a 40 3d 42 3f 40 41 48 44 41 3f 40 43 37 3b 44 2d 49 43 39 44 39 39 3b 45 3d 40 40 40 3d 40 43 43 3c 41 40 45 52 52 45 4b 4b 41 38 25 13 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 1b 2a 30 34 36 38 32 3c 3d 3f 3d 38 38 3a 42 38 34 3d 38 3e 3b 38 3f 3e 3e 44 3c 3a 3f 3d 45 44 3e 41 45 3e 3e 33 3c 3a 40 40 3a 3b 3d 3c 3e 3c 3e 45 42 3a 38 3f 41 44 3c 40 44 3e 3d 45 48 46 39 44 3e 42 41 39 42 4b 4a 4c 46 3f 43 43 42 3e 44 44 45 3d 3c 3c 3d 3d 22 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 2a 38 3c 44 45 3b 44 44 4d 50 4e 51 52 54 52 4a 49 3f 3f 44 43 3e 42 43 40 44 36 42 41 46 3b 3f 45 3a 3e 49 3e 3d 43 3c 43 46 37 3b 3d 3c 33 3d 37 3c 41 3d 3b 44 43 3f 45 4b 41 44 45 46 47 4c 3e 49 3a 32 27 14 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 07 0d 1a 2d 29 38 36 44 42 3a 3a 3f 39 3e 3b 37 3b 3f 39 38 47 3c 42 3a 42 3f 3e 38 3e 39 41 44 46 3e 3d 3e 45 41 3e 39 3c 3d 35 3d 41 44 3c 3c 3e 40 45 40 3f 45 3e 3d 40 36 47 46 3e 3c 40 45 3e 42 44 45 46 42 45 3e 45 44 44 3f 49 46 46 40 3d 3e 48 3d 3e 49 49 44 39 26 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 27 41 41 3d 4a 3e 4f 47 44 52 4d 51 51 4d 4b 44 4a 47 41 4a 3e 46 3c 44 39 3c 3b 43 3e 45 48 45 49 42 3d 42 43 3d 3e 36 42 3d 38 3f 3b 44 44 39 43 3d 3e 47 3e 40 3e 39 3b 41 44 3e 3e 45 4f 45 42 3b 2e 20 1a 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 13 22 2e 37 43 3d 42 3e 44 45 3b 41 39
 39 3f 3d 37 37 41 38 3b 3b 41 3d 43 41 3b 39 3c 40 3d 3c 43 37 3c 41 3c 45 38 3a 3c 3d 44 48 47 40 42 40 48 3c 3b 37 40 3b 39 3e 44 47 47 39 43 43 43 3e 48 4b 41 45 48 42 40 4e 44 49 4b 4a 42 45 45 3b 41 39 49 42 45 35 41 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1f 48 44 42 48 3e 44 4b 49 4a 4e 4f 47 46 44 43 45 47 41 43 3d 43 3e 3e 43 33 41 48 45 43 40 42 43 3d 47 42 3d 3c 39 3e 3b 46 40 44 40 38 40 40 3c 3d 3d 41 3d 3c 44 38 3b 3d 3d 47 4a 46 41 3d 37 2e 1d 13 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 15 1e 22 31 3b 36 44 3b 3a 3b 36 35 3c 37 40 36 3e 38 32 3f 44 3e 38 43 36 35 3b 3a 39 39 3d 47 35 3c 41 33 3c 38 3c 36 3a 35 3a 43 47 3a 38 41 3a 36 3d 3b 3c 34 43 3b 3d 44 38 44 42 42 3a 3f 43 44 43 43 4a 44 47 49 4b 4a 47 51 47 49 3e 44 44 42 43 46 3e 3a 2b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 20 3d 3e 47 49 44 3c 48 44 46 47 46 43 3e 48 42 3e 44 46 43 40 42 40 3d 37 3f 39 3b 3e 37 43 41 40 41 38 39 42 42 40 3c 3a 3f 40 38 3d 38 42 3b 3b 39 3c 38 31 3a 3d 3f 48 45 3e 46 3d 44 47 3b 25 20 0d 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0e 16 28 2d 3f 3c 42 48 36 43 3e 41 3d 40 3e 3b 45 38 3e 33 34 4c 43 42 3f 3c 3e 3e 3d 3a 42 3d 42 31 3b 3b 40 38 44 47 43 37 3c 3b 3d 3a 3c 44 32 3b 36 34 35 3e 3a 42 3a 44 3b 44 3c 3d 4a 42 40 49 48 45 43 41 4d 4e 53 4b 43 46 44 43 48 49 40 45 4b 43 45 47 25 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 40 3f 4c 44 4b 41 47 49 4e 42 4d 3c 43 49 3e 47 3d 42 3d 39 46 44 4a 3a 41 43 39 3f 45 3d 47 39 45 3e 3e 42 44 45 31 3f 3a 40 41 43 3c 3b 45 3e 44 3e 3c 37 43 3e 41 3c 43 3c 3d 3b 43 32 2f 22 0e 04 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 15 26 35 3a 38 3f 3e 37 3a 3f
 40 3a 41 3b 3b 40 37 40 36 35 3d 3d 36 43 40 3f 3d 3c 42 43 3b 41 3f 41 38 42 39 3b 38 32 40 3b 3e 3e 41 3e 3c 3e 3b 41 47 42 43 3e 41 48 37 41 44 43 3f 47 41 47 49 43 46 45 3d 49 49 49 4d 4f 4c 44 49 3d 42 46 44 47 41 44 27 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 1b 42 42 4e 41 4a 48 45 46 45 41 46 4c 45 4c 40 45 4a 40 45 41 3f 41 45 37 44 43 3c 43 3f 3f 41 41 48 43 40 3e 39 3d 38 3e 3e 3e 45 39 3c 44 38 40 47 41 36 45 44 44 3e 42 42 3b 3b 3d 32 28 1f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 1b 22 36 37 3b 38 3b 3e 3b 3b 3c 37 40 3d 35 36 32 39 35 35 31 38 41 40 37 3e 3f 3b 3a 3e 30 3f 43 45 43 40 44 3a 3e 3e 3b 3b 44 41 3b 37 3b 3d 42 42 38 3a 3c 41 41 42 41 3d 3c 3d 45 47 45 48 43 3c 49 38 48 42 45 46 46 46 44 48 43 3c 41 49 3b 40 3e 28 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 19 36 33 4e 49 3e 3c 41 45 48 3c 3a 3b 44 47 44 3f 46 46 47 45 48 3d 3c 3e 3b 3d 35 41 4a 3d 41 40 44 40 41 38 3f 42 44 42 3d 3d 3b 43 3e 3a 3d 40 44 3a 3b 40 46 47 53 43 44 3b 37 32 23 16 0b 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 08 15 24 32 3c 34 34 3e 38 3f 41 38 3e 38 3d 35 40 37 3c 3d 42 39 39 3c 39 3b 3c 46 34 3a 3b 2e 3f 3a 3c 3a 39 3c 3f 3f 44 3c 42 3a 3d 3d 43 3b 40 43 39 3e 46 3a 3f 45 3d 41 3b 3b 41 41 44 41 43 45 46 47 4c 3c 4a 3e 46 4b 41 40 44 46 3e 44 43 49 40 34 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 17 35 49 49 44 3d 39 3d 48 43 42 3c 44 3b 3f 41 3e 41 3f 49 43 4a 46 3f 41 33 3a 3e 46 42 41 46 40 3e 3e 43 4b 46 4a 3b 3b 40 36 39 39 44 37 38 44 3f 40 40 3a 3e 43 3b 40 39 33 2b 1e 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 16 14 26 37 37 36 40 40
 3f 43 3f 3d 39 36 3f 3d 3a 3e 35 3a 38 41 3d 3b 42 3f 3a 3d 44 37 39 3c 39 3b 44 3d 3d 3e 3b 35 3d 3b 3f 42 3c 3f 3c 3a 44 3f 3f 41 37 47 38 40 4a 41 41 4a 4a 43 3f 47 3e 49 42 3f 3e 3f 4b 4a 53 47 4a 42 3f 42 40 41 42 3e 30 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 14 40 4b 4a 47 3d 46 45 48 42 40 42 42 43 42 4a 3e 46 3f 3a 37 3e 40 3c 40 3d 3c 4b 40 41 4c 3d 44 43 3b 46 3d 3e 45 44 3d 43 3d 3e 3a 41 3e 43 45 3a 3c 36 3b 43 40 3b 3a 35 24 1f 0b 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 07 10 15 26 2a 38 3d 43 37 3f 43 3c 41 3e 37 39 3b 39 37 37 34 41 3a 36 3d 3a 3f 3c 34 3b 38 3a 37 40 37 3c 3f 44 3d 3b 38 41 3c 37 3a 39 3f 3e 44 3c 40 3b 3c 45 39 3d 44 41 3e 47 3a 42 4d 3e 44 46 44 45 3c 48 48 46 4b 44 3f 46 41 3f 45 43 40 3e 2a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3b 40 43 4a 48 47 45 42 2d 40 3f 40 46 3f 47 40 3e 47 4b 3f 4f 43 44 3e 3f 48 46 46 45 44 40 38 3e 43 47 47 3c 3b 3b 42 41 3d 3c 41 3b 3f 3f 40 3c 3b 3f 37 37 37 2f 20 25 0f 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 19 21 2b 36 37 3c 44 3d 37 3d 39 39 36 41 34 36 41 3c 3b 37 3a 3f 3a 3f 40 3a 35 3f 3e 3a 30 36 3b 3a 3b 3a 35 3c 37 38 40 39 3a 39 3c 40 39 3c 3f 3f 44 39 41 3b 3a 3d 3c 42 43 42 43 47 3d 45 4a 41 44 49 40 3f 3f 45 44 3f 4a 44 3f 3e 41 2d 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0e 3c 46 4c 45 47 38 3b 39 42 3e 3d 44 42 46 42 3c 47 4b 45 48 44 3b 41 47 3f 40 4b 46 39 41 41 45 3d 41 45 39 43 46 42 3c 3c 3d 40 3f 3e 3d 3a 3b 34 37 35 32 37 2e 25 23 0e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0c 14 1d 27 37
 35 3e 3d 35 37 3b 3c 36 3b 3f 42 44 3a 42 39 35 45 3e 40 40 3b 3f 38 34 41 3e 42 3d 3a 39 3c 44 45 42 46 3c 40 3b 3b 42 38 3a 43 3b 43 3d 38 3f 46 45 47 47 43 41 3b 46 3b 46 49 47 3e 46 47 45 41 42 4c 41 40 41 45 48 43 3b 2f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 09 35 3a 42 4e 43 45 46 4a 4a 43 44 46 49 44 4a 4c 4b 48 49 44 51 48 43 3e 3e 4b 41 44 45 48 44 41 3e 4c 40 45 44 3c 36 3f 43 3c 40 3b 39 42 3a 36 35 31 2d 35 24 17 11 09 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 04 1a 1a 25 2d 33 36 3c 39 41 3f 40 3d 3e 39 41 3c 41 3d 42 36 38 3a 3f 37 36 47 37 41 3b 3b 36 35 40 3d 3e 43 38 37 42 36 3a 3c 3c 3e 39 43 3d 3f 3f 42 47 42 49 47 40 49 47 4a 3f 44 45 43 4b 44 4c 42 42 45 44 45 3e 45 3b 4d 45 3f 35 33 0f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0c 36 3c 43 45 44 4a 4e 46 4d 4e 4a 4c 54 40 4f 54 52 55 4a 56 56 55 56 55 4c 55 4e 4d 4e 4b 4b 48 50 47 38 4c 45 4b 3f 3a 42 45 35 46 38 3d 3e 32 35 2c 2a 1a 17 12 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 07 0e 16 23 2d 32 32 3b 3a 35 33 3f 39 43 3d 3c 3b 3e 46 3d 3b 36 3b 41 42 3f 37 39 35 35 3e 3d 39 3d 3c 3d 3e 3f 3d 39 35 3e 40 3b 3f 42 41 47 3f 3e 3e 47 40 3d 3c 3c 40 44 46 47 40 42 42 42 4a 44 4e 45 40 3e 42 41 39 44 45 3b 41 32 0b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 3b 49 56 50 4c 55 55 4f 5d 5c 62 60 64 62 62 66 63 5f 62 64 6a 6d 6a 5c 65 58 61 5b 54 61 55 59 4b 51 50 4d 4a 4a 4d 4e 48 38 3f 3b 2f 36 2f 2e 26 1a 1b 0f 09 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 12 20 25 2f 2f 3d 38 3f 3a 3c 3d 3f 3b 3c 38 40 3e 3e 3e 3c 3f 41 37 3d 3a 39 3f 3d 38 3e 3c 40 40 3a 41 45 3a 3e 40 39 46 39 45 42 3d 3f 3b 44 4a 45 45 40 40 44 42 48 46 41 46 46 42 51 45 48 3f 3a 46 44 42 46 49 42 49 3e 2a 15 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 48 52 5a 6b 67 65 68 6c 6c 74 6e 6c 74 73 7e 76 79 78 74 7e 79 7a 7b 75 77 76 77 72 74 73 6f 69 64 62 60 5e 56 5f 57 58 51 4b 48 3d 3a 29 20 1f 16 07 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 10 1f 21 25 33 3a 39 38 44 39 3a 3d 36 46 3d 3a 42 37 3b 39 43 40 3b 37 3f 3f 3f 39 3d 3b 3a 43 42 39 43 44 40 40 43 3e 3e 42 37 3f 45 43 42 41 41 47 45 3e 46 3e 42 49 4e 40 42 48 4a 3d 44 47 46 41 3c 42 43 40 45 3d 3b 2d 0d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 14 4f 62 69 7c 73 76 7e 77 7e 71 7b 7a 7e 82 82 83 77 7c 7e 7f 81 7c 84 83 7e 7f 76 7b 78 7e 75 77 75 76 75 71 65 67 60 59 58 47 3f 3b 2f 1d 13 0a 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 06 11 15 22 2b 33 32 3a 35 36 3d 39 44 45 37 3c 39 44 3f 40 3b 30 3c 3e 43 3b 34 3f 3a 3e 3e 3f 3f 3e 3a 43 3f 3a 3f 40 46 42 49 45 3b 41 40 48 41 3e 40 3d 3f 45 42 37 40 46 4a 3e 4a 4d 41 44 45 42 45 3f 43 3d 42 41 38 31 10 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 0b 4f 6e 7e 7e 79 6d 77 7d 7a 7a 79 7d 7a 77 80 7e 81 7e 7d 82 84 7e 81 80 80 7b 84 7f 7e 7e 7b 80 7c 7a 6e 68 68 67 63 5f 56 45 3d 25 1b 16 05 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 02 06 09 16 20 22 28 36 3f 3f 3f 40 43 3e 3e 3b 3e 43 3c 3b 3d 3c 3d 45 3d 3d 3a 33 41 3e 41 45 3d 42 43 44 42 40 4c 3a 3f 43 42 3f 3e 3d 40 47 46 4b 41 47 46 42 49 40 40 49 44 45 4a 47 4a 45 49 45 3d 45 3c 43 44 41 40 37 16 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 56 72 7e 82 7b 78 76 80 77 7b 79 77 7d 7f 80 7c 78 7d 7c 76 81 7f 7d 7b 7f 7a 80 7d 7e 80 74 77 6b 6c 6e 69 65 5f 53 51 38 33 1d 11 06 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0d 0d 19 25 24 31 35 3a 39 3c 3b 3c 36 43 38 3e 3a 3e 40 41 40 3a 43 3c 41 41 41 42 41 3e 46 49 38 45 42 3d 3d 47 48 48 40 4c 3f 46 42 41 4b 47 40 4b 40 45 49 44 47 45 49 42 42 4f 40 4a 49 4a 43 49 4b 43 3a 41 38 1b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 46 6c 71 7e 6f 73 77 71 77 75 7a 7a 7c 7b 7b 78 7d 7c 76 73 74 77 7d 79 76 73 73 76 7f 74 6e 6a 69 6a 64 60 54 47 44 31 24 15 09 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 08 11 1d 2b 26 35 39 3a 44 37 36 3f 3f 44 3f 48 41 3c 49 45 45 3f 40 41 3a 45 40 4b 3f 44 4b 3e 40 45 40 43 48 47 4b 49 48 4a 48 46 49 45 4a 44 48 46 46 43 4e 4c 47 4e 48 49 4b 49 4f 4b 4d 4a 49 4b 47 4f 3f 24 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 45 68 72 72 6f 74 74 70 70 6f 72 71 71 76 71 73 75 71 75 70 72 73 70 72 68 6e 70 67 6f 6a 62 5c 56 55 4d 43 3e 35 24 18 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 01 06 0d 14 24 25 33 3a 3e 3e 44 40 3f 42 49 42 46 3f 44 47 4d 45 42 41 48 44 49 40 42 4a 4f 45 49 4d 49 53 49 4f 4d 48 53 4f 53 57 4d 55 50 4b 50 51 55 51 4b 55 58 5f 54 53 54 52 5a 53 56 52 5c 57 64 5d 53 4a 25 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 3f 5c 6c 75 6d 66 6b 67 6b 69 70 71 76 6d 73 6c 6b 73 71 66 6c 63 6e 66 69 68 63 66 64 5e 5a 53 47 40 3e 2b 1f 1d 0f 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0a 14 1b 25 36 3d 3b 4b 43 45 4a 47 47 4a 4f 4b 55 4f 51 47 4a 50 4a 51 55 57 55 4f 53 56 56 4f 55 53 56 5a 5c 5d 57 57 5f 60 59 5f 67 5d 62 5c 63 61 61 68 69 6f 65 64 68 67 64 66 6a 69 71 6a 68 5f 5e 28 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 38 5a 60 66 65 65 60 71 6b 5e 66 70 67 6b 6e 6a 6f 6f 66 65 68 63 60 64 58 5d 63 51 4d 49 4a 35 36 2b 1f 1a 15 06 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0a 0c 16 21 34 37 40 3c 4a 49 4f 52 4f 55 56 57 5f 51 57 57 53 56 5b 5c 5d 5b 5f 65 64 5e 68 64 5f 5e 6a 65 6c 71 72 6c 69 67 6d 70 78 6e 6d 78 6d 6d 6d 75 76 75 74 71 6d 6c 6e 70 65 72 6e 68 6a 5b 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 32 52 5e 61 5d 5e 61 65 64 5f 5b 62 65 64 65 5a 64 62 60 5a 5b 5b 5b 4e 49 45 4d 43 3f 33 2f 1d 21 0c 02 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 07 12 21 31 3b 42 4b 5b 54 5f 5f 5c 60 68 65 60 5f 5f 69 6f 6c 6b 69 6b 70 76 79 6f 6c 72 71 74 7b 77 76 6c 77 7c 79 7f 84 75 7d 76 78 7c 7b 73 72 75 76 79 79 74 70 6f 79 67 68 75 65 64 5e 55 2e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 2f 56 5e 65 5d 5b 54 5a 54 5e 5f 5d 58 5e 56 4e 52 5b 5b 4d 4a 42 4d 42 39 36 36 2f 26 20 16 14 08 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0c 15 17 24 3c 3f 4a 59 59 63 61 6b 6d 6a 6c 6b 75 76 75 74 72 7b 77 7e 76 80 7c 7a 84 7b 81 7b 79 81 81 7b 81 78 79 7b 78 77 7d 77 76 7a 7d 7e 7a 79 76 6b 73 6c 6e 6c 6c 65 73 73 62 65 5f 2e 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 25 4c 52 5f 5d 4f 5e 54 58 57 52 53 54 50 50 4f 48 45 42 45 41 33 2d 2a 2a 21 1d 17 0c 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0c 0f 22 21 3b 40 4b 51 59 64 62 6d 78 72 77 71 72 74 77 74 79 7b 74 68 7f 76 7d 7b 76 7c 7c 7d 77 7b 74 75 74 75 7b 73 77 77 6a 73 6e 6c 71 71 6f 64 65 6c 69 71 67 6a 5f 6b 69 59 60 5a 2b 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 21 3b 5d 5c 4a 4c 4b 4b 53 55 4c 48 46 43 40 39 3c 3b 2e 29 2b 1d 1d 1c 0c 12 0a 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 0e 20 2a 3b 4e 56 5e 5d 60 66 6e 72 71 74 70 75 71 78 7a 7a 73 6e 70 75 75 7f 72 6b 71 6b 73 70 6d 69 6f 68 6e 6f 6d 64 67 6d 70 74 68 64 68 65 64 65 63 60 5b 62 62 59 5b 50 4b 30 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 0d 3f 45 40 46 3c 3b 41 37 38 40 31 2e 32 29 2b 29 1e 19 0d 11 03 0d 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 07 03 0e 18 2a 2f 42 49 51 5d 62 69 67 62 69 6c 75 71 70 72 72 71 6e 72 6d 71 65 70 6d 69 6d 6d 64 65 62 64 64 64 66 63 57 61 62 6c 68 61 66 5e 61 60 60 5e 5c 60 63 61 54 56 50 52 2f 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 06 30 3b 36 31 31 2f 2c 29 25 1e 24 1c 1b 0a 13 0b 08 09 09 05 0a 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 06 0f 18 1b 2a 28 3b 4e 4f 5a 55 5d 5c 62 66 6c 6d 70 6a 62 69 66 6c 6e 67 62 69 65 5e 60 61 62 63 60 60 60 5f 65 60 5d 5b 64 5f 5a 67 5c 5a 62 58 54 5a 4e 5a 54 59 50 5a 50 2d 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 1b 24 25 17 1a 1e 12 14 0f 0d 06 09 08 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 07 0f 1b 22 20 32 36 3f 4c 54 4b 50 64 5e 60 62 67 63 64 5e 5f 62 60 5a 5c 5e 61 52 58 51 56 54 52 57 5d 5b 59 5c 5a 55 5b 5b 60 57 5f 52 51 54 53 57 53 49 52 47 4b 47 30 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 11 0d 05 0a 0b 06 09 03 00 06 05 03 00 06 06 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 0b 12 15 1c 24 2b 38 47 4a 50 46 4d 50 5b 59 53 52 5c 5f 5a 59 59 53 4a 51 4a 4e 4c 4a 4b 4e 52 56 56 52 5b 4f 5a 57 50 56 52 57 4e 51 4b 4f 51 48 4c 47 44 3f 3e 31 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 02 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 0f 10 12 24 29 26 35 3f 49 40 45 4a 4e 51 4f 49 4b 47 4b 47 44 3c 2d 32 3e 3f 3b 46 46 51 4d 4e 53 54 43 50 49 4c 4e 44 45 43 4a 45 3b 44 35 3b 38 35 37 24 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 05 07 0b 19 10 18 25 31 28 30 39 31 35 38 38 41 3d 3a 38 2b 22 12 1e 1e 23 2f 35 3d 43 47 41 44 39 3f 40 32 3d 3d 3c 37 31 30 33 2c 27 2b 26 24 1c 1d 12 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 04 05 0b 16 15 12 21 1c 2d 26 21 28 2c 29 27 27 16 11 06 11 13 15 19 26 30 29 30 33 29 31 2a 2b 25 27 2b 25 1c 1b 17 14 16 12 10 13 0d 03 07 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 05 00 0c 0e 12 0f 14 11 13 14 12 10 0f 03 06 05 08 02 0b 05 0f 14 19 17 11 10 13 0b 03 0e 06 05 0d 06 06 05 05 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 03 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 04 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 01 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05 03 00 06 05
